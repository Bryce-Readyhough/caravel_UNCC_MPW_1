magic
tech sky130A
timestamp 1608004133
<< metal1 >>
rect 2292 20720 3540 20735
rect 1958 20696 2034 20702
rect 1958 20642 1966 20696
rect 2027 20642 2034 20696
rect 1958 20635 2034 20642
rect 2286 20693 3540 20720
rect 1803 20592 1869 20606
rect 1803 20539 1813 20592
rect 1862 20539 1869 20592
rect 1803 20524 1869 20539
rect 1672 20478 1720 20483
rect 1672 20446 1679 20478
rect 1713 20446 1720 20478
rect 1672 20441 1720 20446
rect 1554 20371 1591 20378
rect 1554 20339 1560 20371
rect 1587 20339 1591 20371
rect 1554 20333 1591 20339
rect 882 20321 938 20332
rect 882 20281 893 20321
rect 927 20281 938 20321
rect 882 20271 938 20281
rect 898 20250 927 20271
rect 894 20145 927 20250
rect 894 20102 923 20145
rect 1566 20143 1588 20333
rect 1555 20125 1597 20143
rect 1686 20136 1705 20441
rect 1823 20138 1840 20524
rect 879 20080 936 20102
rect 1555 20095 1561 20125
rect 1592 20095 1597 20125
rect 1555 20089 1597 20095
rect 1675 20126 1720 20136
rect 1675 20088 1680 20126
rect 1713 20088 1720 20126
rect 1675 20083 1720 20088
rect 1812 20126 1858 20138
rect 1971 20136 1991 20635
rect 879 20045 888 20080
rect 926 20045 936 20080
rect 1812 20081 1816 20126
rect 1854 20081 1858 20126
rect 1812 20077 1858 20081
rect 1953 20123 2011 20136
rect 1953 20071 1957 20123
rect 2006 20071 2011 20123
rect 1953 20066 2011 20071
rect 879 20030 936 20045
rect 2286 10329 2337 20693
rect 4218 20272 4820 20303
rect 2198 10320 2337 10329
rect 2198 10310 2315 10320
rect 4785 10301 4820 20272
rect 4727 10282 4820 10301
rect 4785 10280 4820 10282
<< via1 >>
rect 1966 20642 2027 20696
rect 1813 20539 1862 20592
rect 1679 20446 1713 20478
rect 1560 20339 1587 20371
rect 893 20281 927 20321
rect 1561 20095 1592 20125
rect 1680 20088 1713 20126
rect 888 20045 926 20080
rect 1816 20081 1854 20126
rect 1957 20071 2006 20123
<< metal2 >>
rect 224 20499 260 20836
rect 1243 20821 2039 20825
rect 3664 20821 3694 20824
rect 1243 20796 3694 20821
rect 1243 20793 2039 20796
rect 1246 20508 1283 20793
rect 1960 20697 2037 20705
rect 1960 20642 1965 20697
rect 2030 20642 2037 20697
rect 3664 20691 3694 20796
rect 1960 20636 2037 20642
rect 1801 20596 1871 20604
rect 1801 20533 1807 20596
rect 1863 20533 1871 20596
rect 1801 20527 1871 20533
rect 1245 20499 1283 20508
rect 224 20487 1283 20499
rect 224 20473 1272 20487
rect 224 20052 260 20473
rect 880 20327 937 20345
rect 880 20282 890 20327
rect 929 20282 937 20327
rect 880 20281 893 20282
rect 927 20281 937 20282
rect 880 20272 937 20281
rect 884 20080 940 20085
rect 884 20045 888 20080
rect 926 20045 940 20080
rect 884 20039 940 20045
rect 884 20005 896 20039
rect 928 20005 940 20039
rect 884 19996 940 20005
rect 1245 19948 1272 20473
rect 1674 20485 1723 20491
rect 1674 20444 1677 20485
rect 1719 20444 1723 20485
rect 1674 20439 1723 20444
rect 1547 20404 1605 20417
rect 1547 20368 1555 20404
rect 1594 20368 1605 20404
rect 1547 20358 1560 20368
rect 1552 20339 1560 20358
rect 1587 20358 1605 20368
rect 1587 20339 1598 20358
rect 1552 20332 1598 20339
rect 1554 20127 1599 20134
rect 1554 20093 1560 20127
rect 1591 20125 1599 20127
rect 1592 20095 1599 20125
rect 1591 20093 1599 20095
rect 1554 20087 1599 20093
rect 1676 20126 1719 20132
rect 1676 20088 1680 20126
rect 1713 20088 1719 20126
rect 1676 20083 1719 20088
rect 1811 20126 1861 20135
rect 1811 20081 1816 20126
rect 1854 20081 1861 20126
rect 1811 20077 1861 20081
rect 1953 20123 2011 20128
rect 1953 20071 1957 20123
rect 2006 20071 2011 20123
rect 1953 20066 2011 20071
rect 2163 20025 2786 20056
rect 2169 19950 2219 20025
rect 1483 19948 2227 19950
rect 1243 19920 2227 19948
rect 1243 19919 2106 19920
rect 1243 19912 1516 19919
rect 3773 10237 3829 10240
rect 3689 10230 3829 10237
rect 3668 10196 3829 10230
rect 3668 10194 3801 10196
rect 3668 9949 3716 10194
rect 3306 9948 3716 9949
rect 2918 9946 3716 9948
rect 2852 9936 3716 9946
rect 2852 9891 2862 9936
rect 2909 9916 3716 9936
rect 2909 9914 3714 9916
rect 2909 9913 3326 9914
rect 2909 9891 2926 9913
rect 2852 9877 2926 9891
<< via2 >>
rect 1965 20696 2030 20697
rect 1965 20642 1966 20696
rect 1966 20642 2027 20696
rect 2027 20642 2030 20696
rect 1807 20592 1863 20596
rect 1807 20539 1813 20592
rect 1813 20539 1862 20592
rect 1862 20539 1863 20592
rect 1807 20533 1863 20539
rect 890 20321 929 20327
rect 890 20282 893 20321
rect 893 20282 927 20321
rect 927 20282 929 20321
rect 896 20005 928 20039
rect 1677 20478 1719 20485
rect 1677 20446 1679 20478
rect 1679 20446 1713 20478
rect 1713 20446 1719 20478
rect 1677 20444 1719 20446
rect 1555 20371 1594 20404
rect 1555 20368 1560 20371
rect 1560 20368 1587 20371
rect 1587 20368 1594 20371
rect 1560 20125 1591 20127
rect 1560 20095 1561 20125
rect 1561 20095 1591 20125
rect 1560 20093 1591 20095
rect 1681 20089 1712 20125
rect 1816 20082 1853 20125
rect 1959 20074 2002 20122
rect 2862 9891 2909 9936
<< metal3 >>
rect 1959 20697 2061 20712
rect 1959 20642 1965 20697
rect 2030 20642 2061 20697
rect 1959 20634 2061 20642
rect 1798 20596 1883 20608
rect 1798 20533 1807 20596
rect 1863 20580 1883 20596
rect 1863 20572 2994 20580
rect 1863 20546 3010 20572
rect 1863 20533 1883 20546
rect 1798 20524 1883 20533
rect 1672 20493 1737 20498
rect 1672 20485 2887 20493
rect 1672 20444 1677 20485
rect 1719 20478 2887 20485
rect 1719 20444 2909 20478
rect 1672 20438 1737 20444
rect 1550 20404 1603 20412
rect 1550 20368 1555 20404
rect 1594 20402 1603 20404
rect 1594 20397 2785 20402
rect 1594 20368 2818 20397
rect 875 20327 948 20366
rect 1550 20362 2818 20368
rect 875 20282 890 20327
rect 929 20308 948 20327
rect 929 20294 2730 20308
rect 929 20282 2740 20294
rect 875 20268 2740 20282
rect 875 20266 948 20268
rect 89 20211 2662 20218
rect 89 20187 2664 20211
rect 90 20049 123 20187
rect 1553 20127 1598 20133
rect 1553 20093 1560 20127
rect 1591 20093 1598 20127
rect 1553 20086 1598 20093
rect 1677 20125 1716 20128
rect 1677 20089 1681 20125
rect 1712 20089 1716 20125
rect 1558 19808 1594 20086
rect 1677 19850 1716 20089
rect 1812 20125 1856 20129
rect 1812 20082 1816 20125
rect 1853 20082 1856 20125
rect 1812 19943 1856 20082
rect 1952 20122 2006 20131
rect 1952 20074 1959 20122
rect 2002 20074 2006 20122
rect 1952 20048 2006 20074
rect 1951 20002 2453 20048
rect 2624 20044 2664 20187
rect 2710 20059 2740 20268
rect 2782 20130 2818 20362
rect 2874 20201 2909 20444
rect 2972 20270 3010 20546
rect 4488 20270 4519 20275
rect 2972 20240 4519 20270
rect 2987 20238 4519 20240
rect 2874 20178 4365 20201
rect 2881 20170 4365 20178
rect 2782 20111 4118 20130
rect 2782 20097 4126 20111
rect 2782 20093 2818 20097
rect 2710 20029 3470 20059
rect 2711 20019 3470 20029
rect 4088 20016 4126 20097
rect 1808 19905 2000 19943
rect 1671 19817 1824 19850
rect 1954 19836 1997 19905
rect 1235 10272 1282 10289
rect 2388 10272 2439 20002
rect 4092 19781 4122 20016
rect 4326 19801 4361 20170
rect 4488 19779 4519 20238
rect 1235 10221 2446 10272
rect 1235 10220 1282 10221
rect 1235 10186 1241 10220
rect 1276 10186 1282 10220
rect 1235 10181 1282 10186
rect 2842 9943 2919 9965
rect 2800 9936 2919 9943
rect 2800 9932 2862 9936
rect 2800 9892 2810 9932
rect 2845 9892 2862 9932
rect 2800 9891 2862 9892
rect 2909 9891 2919 9936
rect 2800 9883 2919 9891
<< via3 >>
rect 1241 10186 1276 10220
rect 2810 9892 2845 9932
<< metal4 >>
rect 450 20264 490 20841
rect 1439 20264 3026 20268
rect 450 20259 3026 20264
rect 450 20226 3029 20259
rect 450 20024 490 20226
rect 1439 20224 3029 20226
rect 2991 20174 3029 20224
rect 3797 20174 3835 20322
rect 2991 20133 3868 20174
rect 2991 20038 3029 20133
rect 1233 10225 1288 10228
rect 1223 10220 1289 10225
rect 1223 10186 1241 10220
rect 1276 10209 1289 10220
rect 2271 10209 2317 10214
rect 1276 10186 2317 10209
rect 1223 10167 2317 10186
rect 1289 10154 2317 10167
rect 2271 9923 2317 10154
rect 2802 9932 2852 9953
rect 2802 9923 2810 9932
rect 2271 9892 2810 9923
rect 2845 9892 2852 9932
rect 2271 9883 2852 9892
rect 2271 9880 2317 9883
use 6good  6good_0
timestamp 1608004133
transform 1 0 2 0 1 0
box -3 0 2218 20253
use 6good  6good_1
timestamp 1608004133
transform 1 0 2537 0 1 -28
box -3 0 2218 20253
use Sw-1  Sw-1_0
timestamp 1608004133
transform 1 0 3529 0 1 20226
box -70 45 891 509
<< end >>
