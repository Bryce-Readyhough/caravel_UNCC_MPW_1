* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Include SkyWater sky130 device models
* .include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical__lin.spice"
.include "/foss/pdks/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__cap_var_hvt.model.spice"
* .include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical.spice"
.include "/foss/pdks/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__cap_var_lvt.model.spice"
* .include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"
.include "/foss/pdks/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8__tt.corner.spice"

* DC source for current measure
Vdd vdda1 gnd DC 0.7V
Vgnd vssa1 gnd DC 0.0V
Vth analog_io[10] gnd DC 0.1V
Vk analog_io[9] gnd DC 0.15V
Vw analog_io[11] gnd DC 0.18V
Vr analog_io[8] gnd DC 0.25V
Vau analog_io[12] gnd DC 0.7V
Vad analog_io[7] gnd DC 0.0V

Vdd_aux vdda2 gnd DC 1.8V
Ibias analog_io[6] gnd DC 1n

Vsel analog_io[19] gnd DC 1.8V
Vsyn0 analog_io[13] gnd DC 0.7V
Vsyn1 analog_io[14] gnd DC 0.426V


* Vdd VPWR gnd DC 0.7V
* Vgnd VGND gnd DC 0.0V
* Vth vth gnd DC 0.1V
* Vk vk gnd DC 0.15V
* Vw vw gnd DC 0.01V
* Vr vr gnd DC 0.37V
* Vau vau gnd DC 0.08V
* Vad vad gnd DC 0.25V

Idc vdd analog_io[24] DC 10p

.subckt sky130_fd_pr__nfet_01v8_j74adr VSUBS a_109_249# a_109_337# a_21_289#
X0 a_109_337# a_21_289# a_109_249# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_htftno VSUBS w_n187_n133# a_n184_n57# a_n87_n9# a_n87_n97#
X0 a_n87_n9# a_n184_n57# a_n87_n97# w_n187_n133# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_h5gdbm VSUBS a_n101_295# a_n13_343# a_n13_255#
X0 a_n13_343# a_n101_295# a_n13_255# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_dma3uj VSUBS a_n57_109# a_31_157# a_31_69#
X0 a_31_157# a_n57_109# a_31_69# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_hf7xew VSUBS w_n109_n123# a_n106_n47# a_n9_1# a_n9_n87#
X0 a_n9_1# a_n106_n47# a_n9_n87# w_n109_n123# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_b4l3oq VSUBS a_n11_n3# a_n11_n91# w_n111_n127# a_n108_n51#
X0 a_n11_n3# a_n108_n51# a_n11_n91# w_n111_n127# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_k0ujpa VSUBS a_n151_n105# a_n151_n17# w_n251_n141#
+ a_n248_n65#
X0 a_n151_n17# a_n248_n65# a_n151_n105# w_n251_n141# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lz0viw VSUBS a_n55_313# a_n25_343# a_n25_255#
X0 a_n25_343# a_n55_313# a_n25_255# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt Sw-1 VSUBS li_402_584# w_10_596# w_6_312# li_762_210# w_928_594# w_1442_592#
Xsky130_fd_pr__nfet_01v8_j74adr_0 VSUBS VSUBS li_29_719# li_402_584# sky130_fd_pr__nfet_01v8_j74adr
Xsky130_fd_pr__pfet_01v8_htftno_0 VSUBS w_928_594# li_29_719# w_928_594# w_1442_592#
+ sky130_fd_pr__pfet_01v8_htftno
Xsky130_fd_pr__nfet_01v8_h5gdbm_0 VSUBS li_29_719# w_1442_592# li_762_210# sky130_fd_pr__nfet_01v8_h5gdbm
Xsky130_fd_pr__nfet_01v8_dma3uj_0 VSUBS li_29_719# li_126_470# VSUBS sky130_fd_pr__nfet_01v8_dma3uj
Xsky130_fd_pr__pfet_01v8_hf7xew_0 VSUBS w_10_596# li_29_719# w_10_596# li_126_470#
+ sky130_fd_pr__pfet_01v8_hf7xew
Xsky130_fd_pr__pfet_01v8_b4l3oq_0 VSUBS w_10_596# li_29_719# w_10_596# li_402_584#
+ sky130_fd_pr__pfet_01v8_b4l3oq
Xsky130_fd_pr__pfet_01v8_k0ujpa_0 VSUBS li_762_210# w_1442_592# w_1442_592# li_126_470#
+ sky130_fd_pr__pfet_01v8_k0ujpa
Xsky130_fd_pr__nfet_01v8_lz0viw_0 VSUBS li_126_470# w_928_594# w_1442_592# sky130_fd_pr__nfet_01v8_lz0viw
.ends

* .subckt sky130_fd_pr__res_generic_po_i65fu2 VSUBS a_n33_n244# a_n33_171#
* R0 a_n33_n244# a_n33_171# sky130_fd_pr__res_generic_po w=330000u l=1.71e+06u
* .ends
* 
* .subckt sky130_fd_pr__res_generic_po_kabjgr VSUBS a_n33_n244# a_n33_171#
* R0 a_n33_n244# a_n33_171# sky130_fd_pr__res_generic_po w=330000u l=1.71e+06u
* .ends
* 
* .subckt sky130_fd_pr__res_generic_po_abfehu VSUBS a_n33_n244# a_n33_171#
* R0 a_n33_n244# a_n33_171# sky130_fd_pr__res_generic_po w=330000u l=1.71e+06u
* .ends
* 
* .subckt sky130_fd_pr__res_generic_po_0v6cx5 VSUBS a_n33_n244# a_n33_171#
* R0 a_n33_n244# a_n33_171# sky130_fd_pr__res_generic_po w=330000u l=1.71e+06u
* .ends
* 
* .subckt good VSUBS m3_n30_n637# li_n184_n930# Sw-1_2/w_1442_592# m2_240_n362# li_n184_1324#
* + m4_633_n294# m3_1916_186#
* XSw-1_1 VSUBS m3_n30_n637# m2_240_n362# m4_633_n294# li_n184_n930# li_n184_n588# m1_1880_n536#
* + Sw-1
* XSw-1_0 VSUBS m3_n30_n637# m2_240_n362# m4_633_n294# li_n188_368# li_n188_700# m1_1892_666#
* + Sw-1
* XSw-1_2 VSUBS m3_1916_186# m2_240_n362# m4_633_n294# m1_1880_n536# m1_1892_666# Sw-1_2/w_1442_592#
* + Sw-1
* Xsky130_fd_pr__res_generic_po_i65fu2_0 VSUBS li_n184_n930# li_n184_n588# sky130_fd_pr__res_generic_po_i65fu2
* Xsky130_fd_pr__res_generic_po_kabjgr_0 VSUBS li_n188_368# li_n188_700# sky130_fd_pr__res_generic_po_kabjgr
* Xsky130_fd_pr__res_generic_po_abfehu_0 VSUBS li_n188_700# li_n184_1324# sky130_fd_pr__res_generic_po_abfehu
* Xsky130_fd_pr__res_generic_po_0v6cx5_0 VSUBS li_n184_n588# li_n188_368# sky130_fd_pr__res_generic_po_0v6cx5
* .ends
* 
* .subckt good m4_944_2166# VSUBS m2_426_2318# m3_162_2308# 2good_0/li_n184_n930# m3_1772_2124#
* + m3_2194_2596# Sw-1_0/w_1442_592# 2good_1/li_n184_1324#
* XSw-1_0 VSUBS m3_2194_2596# m2_426_2318# m4_944_2166# m1_3752_2110# m1_3532_3020#
* + Sw-1_0/w_1442_592# Sw-1
* X2good_0 VSUBS m3_162_2308# 2good_0/li_n184_n930# m1_3752_2110# m2_426_2318# 2good_0/li_n184_1324#
* + m4_944_2166# m3_1772_2124# good
* X2good_1 VSUBS m3_162_2308# 2good_0/li_n184_1324# m1_3532_3020# m2_426_2318# 2good_1/li_n184_1324#
* + m4_944_2166# m3_1772_2124# good
* .ends
* 
* .subckt good VSUBS m4_870_4802# Sw-1_0/li_402_584# m3_176_4822# m3_2006_4492# m2_444_4830#
* + m3_1776_4796# 3good_0/2good_0/li_n184_n930# Sw-1_0/w_1442_592# Sw-1_0/w_6_312# Sw-1_0/w_10_596#
* + 3good_1/2good_1/li_n184_1324#
* XSw-1_0 VSUBS Sw-1_0/li_402_584# Sw-1_0/w_10_596# Sw-1_0/w_6_312# m1_3686_4442# m1_3500_5610#
* + Sw-1_0/w_1442_592# Sw-1
* X3good_1 m4_870_4802# VSUBS m2_444_4830# m3_176_4822# 3good_0/2good_1/li_n184_1324#
* + m3_1776_4796# m3_2006_4492# m1_3500_5610# 3good_1/2good_1/li_n184_1324# good
* X3good_0 m4_870_4802# VSUBS m2_444_4830# m3_176_4822# 3good_0/2good_0/li_n184_n930#
* + m3_1776_4796# m3_2006_4492# m1_3686_4442# 3good_0/2good_1/li_n184_1324# good
* .ends
* 
* .subckt good VSUBS Sw-1_0/li_402_584# m3_2200_11718# m3_1870_11066# m3_264_11074#
* + 4good_0/3good_0/2good_0/li_n184_n930# Sw-1_0/w_1442_592# m2_556_6654# 4good_1/3good_1/2good_1/li_n184_1324#
* + m4_958_11006# m3_2296_6328#
* XSw-1_0 VSUBS Sw-1_0/li_402_584# m2_556_6654# m4_958_11006# m1_4054_10970# m1_3814_11892#
* + Sw-1_0/w_1442_592# Sw-1
* X4good_0 VSUBS m4_958_11006# m3_2296_6328# m3_264_11074# m3_2200_11718# m2_556_6654#
* + m3_1870_11066# 4good_0/3good_0/2good_0/li_n184_n930# m1_4054_10970# m4_958_11006#
* + m2_556_6654# 4good_0/3good_1/2good_1/li_n184_1324# good
* X4good_1 VSUBS m4_958_11006# m3_2296_6328# m3_264_11074# m3_2200_11718# m2_556_6654#
* + m3_1870_11066# 4good_0/3good_1/2good_1/li_n184_1324# m1_3814_11892# 4good_1/Sw-1_0/w_6_312#
* + m2_556_6654# 4good_1/3good_1/2good_1/li_n184_1324# good
* .ends
* 
* .subckt good m3_1774_19904# VSUBS m2_458_19930# Sw-1_0/li_402_584# m3_2124_19680#
* + 5good_0/4good_0/3good_0/2good_0/li_n184_n930# m4_850_19908# Sw-1_0/w_1442_592# m3_188_19952#
* + 5good_1/4good_1/3good_1/2good_1/li_n184_1324# m3_2310_19816# m3_1968_19534#
* XSw-1_0 VSUBS Sw-1_0/li_402_584# m2_458_19930# m4_850_19908# m1_4002_19952# m1_3768_20868#
* + Sw-1_0/w_1442_592# Sw-1
* X5good_0 VSUBS m3_2310_19816# m3_1968_19534# m3_1774_19904# m3_188_19952# 5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + m1_4002_19952# m2_458_19930# m1_14_20144# m4_850_19908# m3_2124_19680# good
* X5good_1 VSUBS m3_2310_19816# m3_1968_19534# m3_1774_19904# m3_188_19952# m1_14_20144#
* + m1_3768_20868# m2_458_19930# 5good_1/4good_1/3good_1/2good_1/li_n184_1324# m4_850_19908#
* + m3_2124_19680# good
* .ends
* 
* .subckt good VSUBS Sw-1_0/li_402_584# 6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + 6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930# m1_3606_41048# 6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + m4_900_40048# m1_3108_40666# Sw-1_0/w_1442_592# m1_3906_40132# m1_3344_40882# m3_178_40374#
* + m1_1758_40060# m2_448_40104# 6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* X6good_0 m1_1758_40060# VSUBS m2_448_40104# m1_3906_40132# m1_3344_40882# 6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + m4_900_40048# m1_4396_20620# m3_178_40374# 6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + m1_3606_41048# m1_3108_40666# good
* XSw-1_0 VSUBS Sw-1_0/li_402_584# m2_448_40104# m4_900_40048# m1_8436_40544# m1_4396_20620#
* + Sw-1_0/w_1442_592# Sw-1
* X6good_1 m1_1758_40060# VSUBS m2_448_40104# m1_3906_40132# m1_3344_40882# 6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + m4_900_40048# m1_8436_40544# m3_178_40374# 6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + m1_3606_41048# m1_3108_40666# good
* .ends
* 
* .subckt good VSUBS Sw-1_0/li_402_584# m4_7606_40582# m1_14280_42472# 7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + 7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324# m3_3892_42710# 7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + m1_13190_42260# m2_7304_41624# Sw-1_0/w_1442_592# m1_13882_42250# 7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + m1_12816_42246# 7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930# 7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930# 7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + m1_13522_42238# m1_12404_42242#
* X7good_0 VSUBS m1_14280_42472# 7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + 7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930# m1_13882_42250# 7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + m4_7606_40582# m1_13190_42260# m1_8774_43264# m3_3892_42710# m1_13522_42238# m1_12404_42242#
* + m1_12816_42246# m2_7304_41624# 7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + good
* X7good_1 VSUBS m1_14280_42472# 7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + 7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930# m1_13882_42250# 7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + m4_7606_40582# m1_13190_42260# m1_18694_42308# m3_3892_42710# m1_13522_42238# m1_12404_42242#
* + m1_12816_42246# m2_7304_41624# 7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + good
* XSw-1_0 VSUBS Sw-1_0/li_402_584# m2_7304_41624# m4_7606_40582# m1_18694_42308# m1_8774_43264#
* + Sw-1_0/w_1442_592# Sw-1
* .ends
* 
* .subckt good 8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + VSUBS m1_34870_45168# Sw-1_0/li_402_584# m1_33182_44672# 8good_0/m4_7606_40582#
* + 8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324# m3_15256_44922#
* + m2_36872_44966# 8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324# 8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930# 8good_0/m2_7304_41624#
* + 8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324# m2_32394_46370#
* + 8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930# 8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + m2_32742_46204# m4_37832_42440# Sw-1_0/w_1442_592# 8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + m1_33960_44694# m1_33592_44702# 8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324# 8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324# 8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + m1_34434_44684# 8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* X8good_0 VSUBS m3_15256_44922# 8good_0/m4_7606_40582# m1_34870_45168# 8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + 8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324# m1_34434_44684#
* + 8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324# m1_33182_44672#
* + 8good_0/m2_7304_41624# m1_19068_42976# m1_33960_44694# 8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + m2_32742_46204# 8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930# 8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930# m1_33592_44702#
* + m2_32394_46370# good
* X8good_1 VSUBS m3_15256_44922# m4_37832_42440# m1_34870_45168# 8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + 8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_1324# m1_34434_44684#
* + 8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324# m1_33182_44672#
* + m2_36872_44966# m1_38716_44140# m1_33960_44694# 8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_1324#
* + m1_32720_44664# 8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930# 8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n930#
* + 8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n930# m1_33592_44702#
* + m1_32342_44672# good
* XSw-1_0 VSUBS Sw-1_0/li_402_584# m2_36872_44966# m4_37832_42440# m1_38716_44140# m1_19068_42976#
* + Sw-1_0/w_1442_592# Sw-1
* .ends
* 
* .subckt good VSUBS GND VDD D0 D1 D2 D3 D4 D5 D6 D7 D8 D9
* X9good_0 m1_31884_48# VSUBS D6 D8 D2 GND m1_11882_62# D7 VDD m1_6754_8# m1_16966_2#
* + m1_1684_72# m1_16966_2# VDD m1_26760_28# D0 m1_11882_62# m1_21660_68# D1 GND m1_39076_44800#
* + m1_31884_48# D4 D3 m1_26760_28# VDD m1_21660_68# m1_6754_8# m1_36912_2# D5 m1_1684_72#
* + good
* X9good_1 m1_71736_52# VSUBS D6 D8 D2 GND m1_51780_62# D7 VDD m1_46616_8# m1_56844_12#
* + m1_41532_78# m1_56844_12# VDD m1_66618_22# D0 m1_51780_62# m1_61528_92# D1 GND m1_78452_45530#
* + m1_71736_52# D4 D3 m1_66618_22# m1_36912_2# m1_61528_92# m1_46616_8# m1_76798_18#
* + D5 m1_41532_78# good
* XSw-1_0 VSUBS D9 VDD GND m1_78452_45530# m1_39076_44800# Sw-1_0/w_1442_592# Sw-1
* .ends

.subckt sky130_fd_pr__pfet_01v8_owy61o VSUBS a_n73_n61# w_n109_n123# a_15_n61# a_n33_54#
X0 a_15_n61# a_n33_54# a_n73_n61# w_n109_n123# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_63vi9a VSUBS a_15_n11# a_n33_n99# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt one-way VSUBS li_12_16# w_n37_405# li_100_394#
Xsky130_fd_pr__pfet_01v8_owy61o_0 VSUBS li_12_16# w_n37_405# li_100_394# li_100_394#
+ sky130_fd_pr__pfet_01v8_owy61o
Xsky130_fd_pr__nfet_01v8_63vi9a_0 VSUBS li_100_394# li_12_16# li_12_16# sky130_fd_pr__nfet_01v8_63vi9a
.ends

.subckt sky130_fd_pr__nfet_01v8_8mr83b VSUBS a_n73_n42# a_n15_n68# a_15_n42#
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_ykwexw VSUBS a_n73_n42# w_n109_n104# a_n15_n68# a_15_n42#
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt inverter in out vdd vss
Xsky130_fd_pr__nfet_01v8_8mr83b_0 vss vss in out sky130_fd_pr__nfet_01v8_8mr83b
Xsky130_fd_pr__pfet_01v8_ykwexw_0 vss vdd vdd in out sky130_fd_pr__pfet_01v8_ykwexw
.ends

* .subckt sky130_fd_bs_flash__special_sonosfet_star_ocehe0 VSUBS a_15_n11# a_n33_n99#
* + dw_n429_n439# a_n73_n11#
* X0 a_15_n11# a_n33_n99# a_n73_n11# VSUBS sky130_fd_bs_flash__special_sonosfet_star w=420000u l=150000u
* .ends
* 
* .subckt T-cell gate drain source body sky130_fd_bs_flash__special_sonosfet_star_ocehe0_0/dw_n429_n439#
* Xsky130_fd_bs_flash__special_sonosfet_star_ocehe0_0 body source gate sky130_fd_bs_flash__special_sonosfet_star_ocehe0_0/dw_n429_n439#
* + drain sky130_fd_bs_flash__special_sonosfet_star_ocehe0
* .ends
* 
* .subckt x2-array WL0 WL1 BL0 SL0 BL1 SL1 body nwell body SL1 BL1 BL0 SL0 SL1 body
* + BL1 SL0 body BL0
* X1T-cell_0[0|0] WL1 BL0 SL0 body nwell T-cell
* X1T-cell_0[1|0] WL0 BL0 SL0 body nwell T-cell
* X1T-cell_0[0|1] WL1 BL1 SL1 body nwell T-cell
* X1T-cell_0[1|1] WL0 BL1 SL1 body nwell T-cell
* .ends

.subckt sky130_fd_pr__nfet_01v8_r0atdz VSUBS a_n40_n107# a_n98_n81# a_40_n81#
X0 a_40_n81# a_n40_n107# a_n98_n81# VSUBS sky130_fd_pr__nfet_01v8 w=500000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4pknhj VSUBS a_n98_n86# w_n134_n148# a_40_n86# a_n40_n112#
X0 a_40_n86# a_n40_n112# a_n98_n86# w_n134_n148# sky130_fd_pr__pfet_01v8 w=500000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4ujh9u VSUBS w_n144_n198# a_n50_n162# a_n108_n136#
+ a_50_n136#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_01v8 w=1e+06u l=500000u
.ends

.subckt pmos-diff-amp in_1 in_2 out i_bias vdd vss
Xsky130_fd_pr__nfet_01v8_r0atdz_0 vss m1_91_n137# m1_91_n137# vss sky130_fd_pr__nfet_01v8_r0atdz
Xsky130_fd_pr__nfet_01v8_r0atdz_1 vss m1_91_n137# vss out sky130_fd_pr__nfet_01v8_r0atdz
Xsky130_fd_pr__pfet_01v8_4pknhj_0 vss m1_91_n137# vdd li_184_186# in_1 sky130_fd_pr__pfet_01v8_4pknhj
Xsky130_fd_pr__pfet_01v8_4ujh9u_0 vss vdd i_bias li_184_186# vdd sky130_fd_pr__pfet_01v8_4ujh9u
Xsky130_fd_pr__pfet_01v8_4pknhj_1 vss li_184_186# vdd out in_2 sky130_fd_pr__pfet_01v8_4pknhj
Xsky130_fd_pr__pfet_01v8_4ujh9u_1 vss vdd i_bias vdd i_bias sky130_fd_pr__pfet_01v8_4ujh9u
.ends

.subckt sky130_fd_pr__nfet_01v8_dlksd1 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_s3efqo VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lca7f7 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_u061qr VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_h2n75u VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_zt2j7p VSUBS a_n98_n120# a_n40_n146# a_40_n120# w_n134_n182#
X0 a_40_n120# a_n40_n146# a_n98_n120# w_n134_n182# sky130_fd_pr__pfet_01v8 w=1.2e+06u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ckptud VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_2vaynq VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_wpylm8 VSUBS a_n388_n400# a_n330_n426# a_330_n400#
X0 a_330_n400# a_n330_n426# a_n388_n400# VSUBS sky130_fd_pr__nfet_01v8 w=4e+06u l=3.3e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_9i6r5e VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_9hqhhq VSUBS a_n498_n500# a_n440_n526# a_440_n500#
X0 a_440_n500# a_n440_n526# a_n498_n500# VSUBS sky130_fd_pr__nfet_01v8 w=5e+06u l=4.4e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_h43ndc VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_6z4qh8 VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_tb02ql VSUBS a_n618_n800# a_n560_n826# a_560_n800#
X0 a_560_n800# a_n560_n826# a_n618_n800# VSUBS sky130_fd_pr__nfet_01v8 w=8e+06u l=5.6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_zgaw3c VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt neuron-labeled VPWR VGND vth vk vw vr vau vad v u# a# axon
XM10 VGND VGND vad a# sky130_fd_pr__nfet_01v8_dlksd1
XM11 VGND v a# VGND sky130_fd_pr__nfet_01v8_s3efqo
XM1 VGND a_35_1497# v vth sky130_fd_pr__nfet_01v8_lca7f7
XM2 VGND a_35_1497# VPWR VPWR a_35_1497# sky130_fd_pr__pfet_01v8_u061qr
XM3 VGND a_35_1497# VPWR VPWR v sky130_fd_pr__pfet_01v8_h2n75u
XM4 VGND VPWR a_35_1497# axon VPWR sky130_fd_pr__pfet_01v8_zt2j7p
XM5 VGND VGND a_35_1497# axon sky130_fd_pr__nfet_01v8_ckptud
XM6 VGND vw axon VPWR u# sky130_fd_pr__pfet_01v8_2vaynq
XCu VGND VGND u# VGND sky130_fd_pr__nfet_01v8_wpylm8
XM7 VGND VGND vr u# sky130_fd_pr__nfet_01v8_9i6r5e
XCv VGND VGND v VGND sky130_fd_pr__nfet_01v8_9hqhhq
XM8 VGND v u# VGND sky130_fd_pr__nfet_01v8_h43ndc
XM9 VGND vau axon VPWR a# sky130_fd_pr__pfet_01v8_6z4qh8
XCa VGND VGND a# VGND sky130_fd_pr__nfet_01v8_tb02ql
XMk VGND v vk VGND sky130_fd_pr__nfet_01v8_zgaw3c
.ends

.subckt neuron-labeled-extended-opamp v u a vau vw vth vk vr vad vdd vss axon i_bias
+ v_buff u_buff a_buff axon_buff vdd_aux vss vdd v vss
Xpmos-diff-amp_0 v v_buff v_buff i_bias vdd_aux vss pmos-diff-amp
Xpmos-diff-amp_1 u u_buff u_buff i_bias vdd_aux vss pmos-diff-amp
Xpmos-diff-amp_2 a a_buff a_buff i_bias vdd_aux vss pmos-diff-amp
Xpmos-diff-amp_3 axon axon_buff axon_buff i_bias vdd_aux vss pmos-diff-amp
Xneuron-labeled_0 vdd vss vth vk vw vr vau vad v u a axon neuron-labeled
.ends

.subckt sky130_fd_pr__nfet_01v8_5mkfxl VSUBS a_n73_n42# a_15_n42# a_n33_n130#
X0 a_15_n42# a_n33_n130# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_pa2hmj VSUBS a_n33_n177# a_15_n80# w_n109_n180# a_n73_n80#
X0 a_15_n80# a_n33_n177# a_n73_n80# w_n109_n180# sky130_fd_pr__pfet_01v8 w=800000u l=150000u
.ends

.subckt pass-gate clk clk_bar v_in v_out v_newll v_sub v_out
Xsky130_fd_pr__nfet_01v8_5mkfxl_0 v_sub v_out v_in clk sky130_fd_pr__nfet_01v8_5mkfxl
Xsky130_fd_pr__pfet_01v8_pa2hmj_0 v_sub clk_bar v_out v_newll v_in sky130_fd_pr__pfet_01v8_pa2hmj
.ends

.subckt pass-gate-inv-2 in_1 in_2 clk clk_bar out vdd vss vss vdd clk out in_1 clk
+ vss vss
Xinverter_0 clk clk_bar vdd vss inverter
Xpass-gate_0 clk clk_bar in_1 out vdd vss out pass-gate
Xpass-gate_1 clk_bar clk in_2 out vdd vss out pass-gate
.ends

.subckt chip-w-opamp i_bias vad vr vk vth vw vau vsyn0 vsyn1 vdd vss vdd_aux sel v_syn
+ u_syn a_syn axon_syn v_buff u_buff a_buff axon_buff WL0 WL1 BL0 SL0 BL1 SL1 i_in
+ nwell vdd_aux vss BL0 BL1 SL0 vdd_aux BL0 vdd_aux BL1 WL0 BL0 SL1 SL0 BL1 SL1
Xone-way_0 vss inverter_0/out vdd neuron-labeled-extended-opamp_0/v one-way
Xone-way_1 vss inverter_1/out vdd neuron-labeled-extended-opamp_1/v one-way
Xinverter_0 vsyn0 inverter_0/out vdd vss inverter
Xinverter_1 vsyn1 inverter_1/out vdd vss inverter
* X2x2-array_0 WL0 WL1 BL0 SL0 BL1 SL1 vss nwell vss SL1 BL1 BL0 SL0 SL1 vss BL1 SL0
* + vss BL0 x2-array
Xneuron-labeled-extended-opamp_0 neuron-labeled-extended-opamp_0/v neuron-labeled-extended-opamp_0/u
+ neuron-labeled-extended-opamp_0/a vau vw vth vk vr vad vdd vss neuron-labeled-extended-opamp_0/axon
+ i_bias pass-gate-inv-2_0/in_2 pass-gate-inv-2_1/in_2 pass-gate-inv-2_2/in_2 pass-gate-inv-2_3/in_2
+ vdd_aux vss vdd neuron-labeled-extended-opamp_0/v vss neuron-labeled-extended-opamp
Xneuron-labeled-extended-opamp_1 neuron-labeled-extended-opamp_1/v neuron-labeled-extended-opamp_1/u
+ neuron-labeled-extended-opamp_1/a vau vw vth vk vr vad vdd vss neuron-labeled-extended-opamp_1/axon
+ i_bias pass-gate-inv-2_0/in_1 pass-gate-inv-2_1/in_1 pass-gate-inv-2_2/in_1 pass-gate-inv-2_3/in_1
+ vdd_aux vss vdd neuron-labeled-extended-opamp_1/v vss neuron-labeled-extended-opamp
Xneuron-labeled-extended-opamp_2 i_in neuron-labeled-extended-opamp_2/u neuron-labeled-extended-opamp_2/a
+ vau vw vth vk vr vad vdd vss neuron-labeled-extended-opamp_2/axon i_bias v_buff
+ u_buff a_buff axon_buff vdd_aux vss vdd i_in vss neuron-labeled-extended-opamp
Xpass-gate-inv-2_0 pass-gate-inv-2_0/in_1 pass-gate-inv-2_0/in_2 sel pass-gate-inv-2_0/clk_bar
+ v_syn vdd_aux vss vss vdd_aux sel v_syn pass-gate-inv-2_0/in_1 sel vss vss pass-gate-inv-2
Xpass-gate-inv-2_1 pass-gate-inv-2_1/in_1 pass-gate-inv-2_1/in_2 sel pass-gate-inv-2_1/clk_bar
+ u_syn vdd_aux vss vss vdd_aux sel u_syn pass-gate-inv-2_1/in_1 sel vss vss pass-gate-inv-2
Xpass-gate-inv-2_2 pass-gate-inv-2_2/in_1 pass-gate-inv-2_2/in_2 sel pass-gate-inv-2_2/clk_bar
+ a_syn vdd_aux vss vss vdd_aux sel a_syn pass-gate-inv-2_2/in_1 sel vss vss pass-gate-inv-2
Xpass-gate-inv-2_3 pass-gate-inv-2_3/in_1 pass-gate-inv-2_3/in_2 sel pass-gate-inv-2_3/clk_bar
+ axon_syn vdd_aux vss vss vdd_aux sel axon_syn pass-gate-inv-2_3/in_1 sel vss vss
+ pass-gate-inv-2
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[29]
+ analog_io[2] analog_io[30] analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7]
+ analog_io[8] analog_io[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] user_clock2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2
* X10good_0 vssa1 vssa1 vdda1 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
* + io_in[6] io_in[7] io_in[8] io_in[9] good
Xchip-w-opamp_0 analog_io[6] analog_io[7] analog_io[8] analog_io[9] analog_io[10]
+ analog_io[11] analog_io[12] analog_io[13] analog_io[14] vdda1 vssa1 vdda2 analog_io[19]
+ analog_io[20] analog_io[21] analog_io[22] analog_io[23] analog_io[15] analog_io[16]
+ analog_io[17] analog_io[18] analog_io[1] analog_io[0] analog_io[2] analog_io[3]
+ analog_io[4] analog_io[5] analog_io[24] analog_io[26] vdda2 vssa1 analog_io[2] analog_io[4]
+ analog_io[3] vdda2 analog_io[2] vdda2 analog_io[4] analog_io[1] analog_io[2] analog_io[5]
+ analog_io[3] analog_io[4] analog_io[5] chip-w-opamp
.ends


Xckt analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[29]
+ analog_io[2] analog_io[30] analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7]
+ analog_io[8] analog_io[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] user_clock2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2 user_project_wrapper

.control
* Sweep tran
tran 1u 20m uic
plot v("analog_io[24]") v("analog_io[15]")
.endc
.end
