**.subckt restest
XR1 __UNCONNECTED_PIN__ __UNCONNECTED_PIN__ __UNCONNECTED_PIN__ sky130_fd_pr__res_generic_po W=1 L=1
+ mult=1 m=1
**.ends
.end
