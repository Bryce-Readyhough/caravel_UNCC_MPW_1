magic
tech sky130A
magscale 1 2
timestamp 1606706450
<< error_s >>
rect 430 374 442 380
rect 392 368 448 374
rect 386 362 454 368
rect 386 356 404 362
rect 398 330 404 356
rect 436 356 454 362
rect 436 330 448 356
rect 398 324 448 330
rect 430 318 448 324
rect 430 312 442 318
rect 2404 -116 2416 -110
rect 2366 -122 2422 -116
rect 2360 -128 2428 -122
rect 2360 -134 2378 -128
rect 2372 -160 2378 -134
rect 2410 -134 2428 -128
rect 2410 -160 2422 -134
rect 2372 -166 2422 -160
rect 2404 -172 2422 -166
rect 2404 -178 2416 -172
rect 424 -974 436 -968
rect 386 -980 442 -974
rect 380 -986 448 -980
rect 380 -992 398 -986
rect 392 -1018 398 -992
rect 430 -992 448 -986
rect 430 -1018 442 -992
rect 392 -1024 442 -1018
rect 424 -1030 442 -1024
rect 424 -1036 436 -1030
<< locali >>
rect -66 -12 0 28
rect -70 -54 -60 -12
rect -4 -54 6 -12
rect -66 -70 0 -54
rect -66 -352 2 -346
rect -72 -392 -62 -352
rect -2 -392 8 -352
rect -66 -414 2 -392
<< viali >>
rect -60 -54 -4 -12
rect -62 -392 -2 -352
<< metal1 >>
rect 1894 686 2124 730
rect 2068 448 2124 686
rect -78 -8 14 0
rect 72 -8 118 56
rect -78 -12 118 -8
rect -78 -54 -60 -12
rect -4 -48 118 -12
rect -4 -54 88 -48
rect -78 -58 88 -54
rect -78 -68 14 -58
rect -78 -328 14 -324
rect -78 -334 76 -328
rect -78 -352 112 -334
rect -78 -392 -62 -352
rect -2 -370 112 -352
rect -2 -392 14 -370
rect -78 -408 14 -392
rect 68 -432 112 -370
rect 2072 -618 2114 -428
rect 1878 -662 2114 -618
<< metal2 >>
rect 372 458 442 912
rect 372 390 2424 458
rect 372 388 2022 390
rect 372 -466 442 388
<< metal4 >>
rect 650 -320 728 170
rect 650 -390 2711 -320
rect 650 -1224 728 -390
use sky130_fd_pr__res_generic_po_9ekftz  sky130_fd_pr__res_generic_po_9ekftz_0
timestamp 1606706199
transform 1 0 -33 0 1 -200
box -33 -244 33 244
use Sw-1  Sw-1_0
timestamp 1606706242
transform 1 0 118 0 1 -66
box -140 90 1782 1018
use Sw-1  Sw-1_1
timestamp 1606706242
transform 1 0 112 0 1 -1414
box -140 90 1782 1018
use Sw-1  Sw-1_2
timestamp 1606706242
transform 1 0 2092 0 1 -556
box -140 90 1782 1018
<< end >>
