magic
tech sky130A
timestamp 1607535698
<< metal1 >>
rect 36077 24683 36179 24689
rect 36077 24624 36087 24683
rect 36169 24624 36179 24683
rect 36077 24615 36179 24624
rect 36088 23541 36144 24615
rect 36247 24550 36349 24557
rect 36247 24491 36256 24550
rect 36338 24491 36349 24550
rect 36247 24483 36349 24491
rect 36069 23527 36190 23541
rect 36268 23538 36326 24483
rect 36492 24423 36594 24432
rect 36492 24364 36501 24423
rect 36583 24364 36594 24423
rect 36492 24358 36594 24364
rect 36069 23462 36077 23527
rect 36180 23462 36190 23527
rect 36069 23456 36190 23462
rect 36267 23526 36388 23538
rect 36503 23531 36556 24358
rect 36703 24294 36805 24301
rect 36703 24235 36712 24294
rect 36794 24235 36805 24294
rect 36703 24227 36805 24235
rect 36712 23536 36778 24227
rect 36884 24160 36986 24167
rect 36884 24101 36894 24160
rect 36976 24101 36986 24160
rect 36884 24093 36986 24101
rect 36267 23461 36276 23526
rect 36379 23461 36388 23526
rect 36267 23453 36388 23461
rect 36482 23518 36603 23531
rect 36482 23453 36491 23518
rect 36594 23453 36603 23518
rect 36482 23446 36603 23453
rect 36687 23522 36808 23536
rect 36902 23533 36960 24093
rect 37125 24039 37227 24048
rect 37125 23980 37134 24039
rect 37216 23980 37227 24039
rect 37125 23974 37227 23980
rect 37146 23536 37202 23974
rect 37321 23926 37423 23931
rect 37321 23867 37330 23926
rect 37412 23867 37423 23926
rect 37321 23857 37423 23867
rect 36687 23457 36696 23522
rect 36799 23457 36808 23522
rect 36687 23451 36808 23457
rect 36888 23520 37009 23533
rect 36888 23455 36897 23520
rect 37000 23455 37009 23520
rect 36888 23448 37009 23455
rect 37107 23522 37228 23536
rect 37339 23534 37392 23857
rect 37894 23808 37996 23813
rect 37894 23749 37904 23808
rect 37986 23749 37996 23808
rect 37894 23739 37996 23749
rect 37922 23542 37973 23739
rect 37107 23457 37117 23522
rect 37220 23457 37228 23522
rect 37107 23451 37228 23457
rect 37313 23525 37434 23534
rect 37313 23460 37323 23525
rect 37426 23460 37434 23525
rect 37313 23449 37434 23460
rect 37890 23532 38011 23542
rect 37890 23467 37899 23532
rect 38002 23467 38011 23532
rect 37890 23457 38011 23467
rect 38116 23240 38623 23252
rect 38080 23218 38623 23240
rect 19538 22400 19845 22437
rect 19811 22238 19844 22400
rect 25000 22238 35867 22247
rect 19811 22223 35867 22238
rect 38080 22223 38134 23218
rect 39226 22765 39506 22811
rect 39466 22399 39506 22765
rect 19811 22211 38134 22223
rect 19811 22202 30678 22211
rect 19811 22199 19844 22202
rect 35540 22171 38134 22211
rect 35540 22165 38116 22171
rect 10 20301 67 21446
rect 10 20277 340 20301
rect 2552 20277 2809 20284
rect 19 20269 340 20277
rect 310 20116 340 20269
rect 2402 20274 2809 20277
rect 2402 20252 2822 20274
rect 576 20116 681 20162
rect 310 20082 681 20116
rect 310 20079 587 20082
rect 310 20077 340 20079
rect 2406 73 2424 20252
rect 2552 20247 2822 20252
rect 2787 20100 2822 20247
rect 2785 20065 2822 20100
rect 2798 20058 3093 20065
rect 3182 20058 3236 20337
rect 5131 20309 5187 20497
rect 5001 20298 5187 20309
rect 5001 20263 5226 20298
rect 7528 20265 7688 20284
rect 8269 20281 8343 20396
rect 9994 20304 10041 20400
rect 9953 20301 10041 20304
rect 9953 20288 10059 20301
rect 7828 20265 8343 20281
rect 5001 20261 5187 20263
rect 5001 20251 5161 20261
rect 4999 20229 5161 20251
rect 7528 20236 8343 20265
rect 7521 20232 8343 20236
rect 2798 20030 3607 20058
rect 2798 20029 2812 20030
rect 3083 20028 3607 20030
rect 842 36 2443 73
rect 4999 61 5017 20229
rect 7521 20204 7688 20232
rect 7828 20230 8343 20232
rect 8269 20223 8343 20230
rect 9945 20273 10059 20288
rect 9945 20264 10035 20273
rect 7521 69 7539 20204
rect 9945 128 9963 20264
rect 12534 20262 12807 20269
rect 2406 35 2424 36
rect 3377 12 5017 61
rect 5941 31 7539 69
rect 3377 4 5009 12
rect 7521 -3 7539 31
rect 9923 49 9963 128
rect 12450 20239 12807 20262
rect 12450 20219 12565 20239
rect 12450 66 12468 20219
rect 12774 20068 12806 20239
rect 13208 20069 13265 20371
rect 15096 20292 15161 20415
rect 19866 20403 19915 20411
rect 19866 20371 19875 20403
rect 19906 20386 19915 20403
rect 19948 20386 19986 20393
rect 19906 20377 19986 20386
rect 19906 20372 19973 20377
rect 19906 20371 19915 20372
rect 19866 20364 19915 20371
rect 19953 20302 19973 20372
rect 29887 20303 30013 20308
rect 15024 20271 15175 20292
rect 13039 20068 13265 20069
rect 12774 20048 13265 20068
rect 15023 20263 15175 20271
rect 17642 20265 17895 20269
rect 19948 20266 20339 20302
rect 24988 20285 25114 20295
rect 29887 20289 30269 20303
rect 15023 20249 15139 20263
rect 17584 20258 17895 20265
rect 12774 20041 13261 20048
rect 12774 20039 13062 20041
rect 12774 20034 12806 20039
rect 9923 24 9958 49
rect 10830 34 12482 66
rect 15023 46 15041 20249
rect 17584 20240 17898 20258
rect 17582 20235 17898 20240
rect 17582 20222 17699 20235
rect 17582 56 17600 20222
rect 17867 20061 17898 20235
rect 20304 20099 20338 20266
rect 22390 20264 22516 20267
rect 22390 20262 22731 20264
rect 22390 20232 22758 20262
rect 24988 20256 25435 20285
rect 29887 20282 30275 20289
rect 29880 20270 30275 20282
rect 27517 20258 27643 20270
rect 24988 20236 25114 20256
rect 22390 20208 22516 20232
rect 20304 20068 20575 20099
rect 20320 20067 20575 20068
rect 17863 20031 17899 20061
rect 17863 20021 18232 20031
rect 17866 20001 18232 20021
rect 19866 10259 19912 10266
rect 19866 10225 19872 10259
rect 19904 10225 19912 10259
rect 19866 10220 19912 10225
rect 19875 10219 19908 10220
rect 19893 56 19908 10219
rect 22391 59 22408 20208
rect 22715 20076 22758 20232
rect 22715 20045 23476 20076
rect 24993 71 25010 20236
rect 25395 20098 25431 20256
rect 27517 20224 27983 20258
rect 27517 20211 27643 20224
rect 25395 20064 25786 20098
rect 25395 20062 25431 20064
rect 8483 1 9963 24
rect 12450 12 12468 34
rect 13380 32 15041 46
rect 13380 14 15032 32
rect 15942 24 17600 56
rect 19864 35 19908 56
rect 20766 39 22408 59
rect 19864 29 19906 35
rect 17582 1 17600 24
rect 18456 1 19906 29
rect 22391 26 22408 39
rect 24945 27 25010 71
rect 27520 54 27537 20211
rect 27930 20068 27983 20224
rect 29880 20249 30013 20270
rect 27930 20037 28675 20068
rect 27930 20031 27983 20037
rect 29880 93 29897 20249
rect 30216 20126 30275 20270
rect 32391 20284 32517 20303
rect 34963 20297 35089 20303
rect 32391 20267 32865 20284
rect 32389 20262 32865 20267
rect 32389 20244 32866 20262
rect 34963 20260 35460 20297
rect 37503 20260 37629 20278
rect 34963 20244 35089 20260
rect 30216 20080 30640 20126
rect 30243 20078 30640 20080
rect 25890 31 27542 54
rect 29872 44 29897 93
rect 32389 74 32406 20244
rect 32468 20236 32866 20244
rect 32811 20092 32866 20236
rect 32811 20055 33787 20092
rect 32823 20053 33787 20055
rect 34971 116 34988 20244
rect 35403 20102 35454 20260
rect 37503 20222 37934 20260
rect 37503 20219 37629 20222
rect 35403 20064 35777 20102
rect 30764 46 32406 74
rect 23308 4 25010 27
rect 27520 1 27537 31
rect 29872 29 29890 44
rect 32389 29 32406 46
rect 34891 84 34988 116
rect 34891 36 34983 84
rect 37503 51 37520 20219
rect 37906 20096 37933 20222
rect 37906 20064 38785 20096
rect 37906 20059 37933 20064
rect 28422 6 29902 29
rect 33309 16 34983 36
rect 35868 26 37520 51
rect 39939 39 39969 24870
rect 37503 21 37520 26
rect 33309 11 34921 16
rect 38399 9 39997 39
rect 9923 -4 9958 1
rect 19864 -11 19906 1
<< via1 >>
rect 36087 24624 36169 24683
rect 36256 24491 36338 24550
rect 36501 24364 36583 24423
rect 36077 23462 36180 23527
rect 36712 24235 36794 24294
rect 36894 24101 36976 24160
rect 36276 23461 36379 23526
rect 36491 23453 36594 23518
rect 37134 23980 37216 24039
rect 37330 23867 37412 23926
rect 36696 23457 36799 23522
rect 36897 23455 37000 23520
rect 37904 23749 37986 23808
rect 37117 23457 37220 23522
rect 37323 23460 37426 23525
rect 37899 23467 38002 23532
rect 19875 20371 19906 20403
rect 19872 10225 19904 10259
<< metal2 >>
rect 36077 24683 36178 24690
rect 36077 24624 36087 24683
rect 36169 24624 36178 24683
rect 36077 24622 36088 24624
rect 36166 24622 36178 24624
rect 36077 24615 36178 24622
rect 36249 24550 36350 24558
rect 36249 24491 36256 24550
rect 36338 24491 36350 24550
rect 36249 24483 36350 24491
rect 36491 24424 36592 24432
rect 36491 24366 36500 24424
rect 36578 24423 36592 24424
rect 36491 24364 36501 24366
rect 36583 24364 36592 24423
rect 36491 24357 36592 24364
rect 36701 24294 36802 24301
rect 36701 24235 36712 24294
rect 36794 24235 36802 24294
rect 36701 24226 36802 24235
rect 36883 24162 36984 24168
rect 36883 24160 36896 24162
rect 36974 24160 36984 24162
rect 36883 24101 36894 24160
rect 36976 24101 36984 24160
rect 36883 24093 36984 24101
rect 37123 24040 37224 24049
rect 37123 24039 37135 24040
rect 37213 24039 37224 24040
rect 37123 23980 37134 24039
rect 37216 23980 37224 24039
rect 37123 23974 37224 23980
rect 37322 23926 37423 23935
rect 37322 23868 37329 23926
rect 37322 23867 37330 23868
rect 37412 23867 37423 23926
rect 37322 23860 37423 23867
rect 37895 23808 37996 23814
rect 37895 23749 37904 23808
rect 37986 23749 37996 23808
rect 37895 23739 37996 23749
rect 36069 23527 36191 23537
rect 36069 23462 36077 23527
rect 36180 23462 36191 23527
rect 36069 23455 36191 23462
rect 36266 23526 36388 23537
rect 36266 23461 36276 23526
rect 36379 23461 36388 23526
rect 36266 23455 36388 23461
rect 36478 23518 36600 23528
rect 36478 23515 36491 23518
rect 36478 23453 36488 23515
rect 36594 23453 36600 23518
rect 36478 23446 36600 23453
rect 36686 23522 36808 23531
rect 36686 23457 36696 23522
rect 36799 23457 36808 23522
rect 36686 23449 36808 23457
rect 36886 23520 37008 23529
rect 36886 23455 36897 23520
rect 37000 23455 37008 23520
rect 36886 23447 37008 23455
rect 37106 23522 37228 23533
rect 37890 23532 38012 23540
rect 37106 23521 37117 23522
rect 37106 23459 37116 23521
rect 37106 23457 37117 23459
rect 37220 23457 37228 23522
rect 37106 23451 37228 23457
rect 37312 23525 37434 23531
rect 37312 23518 37323 23525
rect 37312 23456 37322 23518
rect 37426 23460 37434 23525
rect 37424 23456 37434 23460
rect 37890 23465 37899 23532
rect 38002 23467 38012 23532
rect 38001 23465 38012 23467
rect 37890 23458 38012 23465
rect 37312 23449 37434 23456
rect 38362 23301 38701 23313
rect 38362 23274 38709 23301
rect 38363 22418 38403 23274
rect 38664 23192 38709 23274
rect -369 20778 258 20863
rect 8763 20821 10246 20854
rect 18754 20819 20188 20860
rect 28696 20812 30174 20873
rect 19869 20403 19913 20413
rect 19869 20371 19875 20403
rect 19906 20371 19913 20403
rect 19869 20365 19913 20371
rect 19879 10266 19898 20365
rect 19868 10259 19914 10266
rect 19868 10225 19872 10259
rect 19904 10225 19914 10259
rect 19868 10217 19914 10225
<< via2 >>
rect 36088 24624 36166 24680
rect 36088 24622 36166 24624
rect 36257 24491 36335 24549
rect 36500 24423 36578 24424
rect 36500 24366 36501 24423
rect 36501 24366 36578 24423
rect 36713 24236 36791 24294
rect 36896 24160 36974 24162
rect 36896 24104 36974 24160
rect 37135 24039 37213 24040
rect 37135 23982 37213 24039
rect 37329 23868 37330 23926
rect 37330 23868 37407 23926
rect 37905 23749 37983 23807
rect 36078 23465 36180 23527
rect 36277 23461 36379 23523
rect 36488 23453 36491 23515
rect 36491 23453 36590 23515
rect 36697 23459 36799 23521
rect 36897 23456 36999 23518
rect 37116 23459 37117 23521
rect 37117 23459 37218 23521
rect 37322 23460 37323 23518
rect 37323 23460 37424 23518
rect 37322 23456 37424 23460
rect 37899 23467 38001 23527
rect 37899 23465 38001 23467
<< metal3 >>
rect 16185 24680 36178 24687
rect 16185 24622 36088 24680
rect 36166 24622 36178 24680
rect 16185 24615 36178 24622
rect 16197 24475 16275 24615
rect 16354 24549 36347 24556
rect 16354 24491 36257 24549
rect 36335 24491 36347 24549
rect 16354 24484 36347 24491
rect 16188 24457 16275 24475
rect 16188 23184 16272 24457
rect 16372 24393 16461 24484
rect 16366 24384 16461 24393
rect 16597 24424 36590 24432
rect 16366 23102 16450 24384
rect 16597 24366 36500 24424
rect 36578 24366 36590 24424
rect 16597 24360 36590 24366
rect 16606 24270 16695 24360
rect 16809 24294 36802 24301
rect 16610 23000 16694 24270
rect 16809 24244 36713 24294
rect 16799 24236 36713 24244
rect 36791 24236 36802 24294
rect 16799 24229 36802 24236
rect 16799 24160 16893 24229
rect 16990 24162 36983 24170
rect 16803 22890 16887 24160
rect 16990 24135 36896 24162
rect 16988 24104 36896 24135
rect 36974 24104 36983 24162
rect 16988 24098 36983 24104
rect 16988 24082 17082 24098
rect 16987 24051 17082 24082
rect 16987 22791 17071 24051
rect 17227 24040 37220 24048
rect 17227 23982 37135 24040
rect 37213 23982 37220 24040
rect 17227 23976 37220 23982
rect 17227 22691 17311 23976
rect 17424 23926 37417 23933
rect 17424 23868 37329 23926
rect 37407 23868 37417 23926
rect 17424 23861 37417 23868
rect 17433 22582 17517 23861
rect 17998 23807 37991 23814
rect 17998 23764 37905 23807
rect 17995 23749 37905 23764
rect 37983 23749 37991 23807
rect 17995 23742 37991 23749
rect 17995 22466 18079 23742
rect 18294 23682 38207 23686
rect 18294 23670 38263 23682
rect 18180 23599 38263 23670
rect 18180 22382 18260 23599
rect 36066 23527 36193 23539
rect 36066 23465 36078 23527
rect 36180 23465 36193 23527
rect 36066 23451 36193 23465
rect 36263 23523 36390 23539
rect 36263 23461 36277 23523
rect 36379 23461 36390 23523
rect 36263 23451 36390 23461
rect 36477 23515 36604 23532
rect 36477 23453 36488 23515
rect 36590 23453 36604 23515
rect 36116 23205 36171 23451
rect 36308 23122 36358 23451
rect 36477 23444 36604 23453
rect 36685 23521 36812 23537
rect 36685 23459 36697 23521
rect 36799 23459 36812 23521
rect 36685 23449 36812 23459
rect 36884 23518 37011 23530
rect 36884 23456 36897 23518
rect 36999 23456 37011 23518
rect 36540 23023 36601 23444
rect 36741 22911 36802 23449
rect 36884 23442 37011 23456
rect 37104 23521 37231 23534
rect 37104 23459 37116 23521
rect 37218 23459 37231 23521
rect 37104 23446 37231 23459
rect 37312 23518 37439 23534
rect 37312 23456 37322 23518
rect 37424 23456 37439 23518
rect 37312 23446 37439 23456
rect 37886 23527 38013 23540
rect 37886 23465 37899 23527
rect 38001 23465 38013 23527
rect 37886 23452 38013 23465
rect 36916 22810 36988 23442
rect 37150 22702 37215 23446
rect 37355 22594 37433 23446
rect 37922 22468 38002 23452
rect 38188 22393 38263 23599
rect 38430 23023 38495 23635
rect 18180 22322 18618 22382
rect 38188 22333 38551 22393
rect 18180 22319 18260 22322
<< metal4 >>
rect 38809 22844 38877 22859
rect 38809 22775 38912 22844
rect 38854 22090 38912 22775
rect -355 21041 499 21110
rect 449 20823 499 21041
rect 8923 20137 9004 20218
rect 8923 20087 10466 20137
rect 18759 20110 20417 20186
rect 28739 20130 30397 20206
rect 8944 20078 10466 20087
use 9good  9good_1
timestamp 1607535698
transform 1 0 19934 0 1 3
box -3 -1 19911 23259
use 9good  9good_0
timestamp 1607535698
transform 1 0 2 0 1 1
box -3 -1 19911 23259
use Sw-1  Sw-1_0
timestamp 1607535698
transform 1 0 38534 0 1 22730
box -70 45 891 509
<< labels >>
rlabel metal4 -339 21054 -292 21094 1 GND
rlabel metal2 -349 20793 -302 20833 1 VDD
rlabel metal1 22 21391 53 21431 1 VREF
rlabel metal3 36018 24628 36049 24668 1 D0
rlabel metal3 36201 24502 36232 24542 1 D1
rlabel metal3 36429 24379 36460 24419 1 D2
rlabel metal3 36648 24238 36679 24278 1 D3
rlabel metal3 36842 24111 36873 24151 1 D4
rlabel metal3 37059 23993 37090 24033 1 D5
rlabel metal3 37254 23880 37285 23920 1 D6
rlabel metal3 37446 23756 37477 23796 1 D7
rlabel metal3 37591 23618 37622 23658 1 D8
rlabel metal3 38444 23562 38475 23602 1 D9
<< end >>
