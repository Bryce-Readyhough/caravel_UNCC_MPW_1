.include "/shared/PDK-ROOT-11242020/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"
.model sky130_fd_pr__res_generic_po1 R ( TC1=0 TC2=0 Rsh = 48.2 NARROW=0.0 TNOM=27 )

valpha  VREF Gnd 3.3
vbeta  VDD Gnd 3.3
vzero D0 Gnd pulse(0 1.8 0.1m 60p 60p 0.1m 0.2m)
vone  D1 Gnd pulse(0 1.8 0.2m 60p 60p 0.2m 0.4m)
vtwo  D2 Gnd pulse(0 1.8 0.4m 60p 60p 0.4m 0.8m)
vthree D3 Gnd pulse(0 1.8 0.8m 60p 60p 0.8m 1.6m)
vfour D4 Gnd pulse (0 1.8 1.6m 60p 60p 1.6m 3.2m)
vfive D5 Gnd pulse (0 1.8 3.2m 60p 60p 3.2m 6.4m)
vsix D6 Gnd pulse (0 1.8 6.4m 60p 60p 6.4m 12.8m)
vseven D7 Gnd pulse (0 1.8 12.8m 60p 60p 12.8m 25.6m)
veight D8 Gnd pulse (0 1.8 25.6m 60p 60p 25.6m 51.2m)
vnine D9 Gnd pulse (0 1.8 51.2m 60p 60p 51.2m 102.4m)
.tran 0.01m 102.4m
.control
run

plot V(Y) V(D0)

.endc
.end




* SPICE3 file created from 10good.ext - technology: sky130A

.option scale=5000u

X0 9good_0/8good_0/7good_0/Sw-1_0/li_29_719# D6 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1 9good_0/8good_0/7good_0/m1_4396_20620# 9good_0/8good_0/7good_0/Sw-1_0/li_29_719# 9good_0/8good_0/m1_8774_43264# 9good_0/8good_0/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X2 9good_0/8good_0/m1_8774_43264# 9good_0/8good_0/7good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3 9good_0/8good_0/7good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4 VDD 9good_0/8good_0/7good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5 VDD D6 9good_0/8good_0/7good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6 9good_0/8good_0/m1_8774_43264# 9good_0/8good_0/7good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/m1_8436_40544# 9good_0/8good_0/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X7 9good_0/8good_0/7good_0/m1_4396_20620# 9good_0/8good_0/7good_0/Sw-1_0/li_126_470# 9good_0/8good_0/m1_8774_43264# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X9 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/m1_4396_20620# 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X10 9good_0/8good_0/7good_0/m1_4396_20620# 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X11 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X12 VDD 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X13 VDD D5 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X14 9good_0/8good_0/7good_0/m1_4396_20620# 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 9good_0/8good_0/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X15 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/m1_4396_20620# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X16 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X17 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X18 9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X19 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X20 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X21 VDD D4 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X22 9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 9good_0/8good_0/7good_0/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X23 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X24 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X25 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X26 9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X27 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X28 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X29 VDD D3 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X30 9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X31 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X32 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X33 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X34 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X35 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X36 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X37 VDD D2 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X38 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X39 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X40 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X41 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X42 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X43 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X44 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X45 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X46 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X47 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X48 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X49 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X50 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_1684_72# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X51 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X52 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X53 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X54 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_1684_72# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X55 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X56 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X57 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X58 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X59 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X60 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X61 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X62 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X63 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R0 m1_1684_72# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R2 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R3 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X64 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X65 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X66 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X67 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X68 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X69 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X70 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X71 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X72 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X73 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X74 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X75 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X76 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X77 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X78 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X79 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X80 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X81 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X82 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X83 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X84 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X85 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X86 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X87 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R4 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R5 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R6 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R7 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X88 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X89 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X90 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X91 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X92 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X93 VDD D2 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X94 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X95 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X96 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X97 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X98 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X99 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X100 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X101 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X102 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X103 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X104 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X105 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X106 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X107 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X108 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X109 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X110 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X111 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X112 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X113 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X114 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X115 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X116 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X117 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X118 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X119 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R8 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R9 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R10 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R11 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X120 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X121 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X122 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X123 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X124 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X125 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X126 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X127 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X128 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X129 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X130 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X131 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X132 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X133 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X134 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X135 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X136 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X137 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X138 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X139 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X140 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X141 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X142 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X143 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R12 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R13 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R14 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R15 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X144 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X145 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X146 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X147 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X148 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X149 VDD D3 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X150 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X151 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X152 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X153 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X154 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X155 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X156 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X157 VDD D2 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X158 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X159 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X160 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X161 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X162 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X163 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X164 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X165 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X166 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X167 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X168 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X169 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X170 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X171 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X172 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X173 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X174 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X175 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X176 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X177 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X178 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X179 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X180 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X181 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X182 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X183 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R16 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R17 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R18 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R19 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X184 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X185 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X186 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X187 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X188 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X189 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X190 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X191 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X192 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X193 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X194 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X195 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X196 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X197 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X198 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X199 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X200 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X201 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X202 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X203 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X204 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X205 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X206 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X207 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R20 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R21 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R22 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R23 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X208 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X209 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X210 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X211 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X212 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X213 VDD D2 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X214 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X215 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X216 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X217 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X218 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X219 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X220 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X221 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X222 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X223 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X224 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X225 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X226 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X227 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X228 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X229 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X230 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X231 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X232 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X233 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X234 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X235 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X236 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X237 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X238 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X239 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R24 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R25 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R26 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R27 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X240 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X241 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X242 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X243 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X244 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X245 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X246 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X247 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X248 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X249 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X250 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X251 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X252 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X253 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X254 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X255 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X256 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X257 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X258 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X259 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X260 VDD 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X261 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X262 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X263 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R28 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R29 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R30 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R31 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X264 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X265 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X266 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X267 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X268 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X269 VDD D4 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X270 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X271 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X272 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X273 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X274 9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X275 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X276 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X277 VDD D3 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X278 9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X279 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X280 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X281 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X282 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X283 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X284 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X285 VDD D2 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X286 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X287 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X288 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X289 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X290 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X291 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X292 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X293 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X294 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X295 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X296 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X297 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X298 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X299 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X300 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X301 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X302 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/m1_14_20144# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X303 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X304 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X305 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X306 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X307 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X308 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X309 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X310 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X311 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R32 9good_0/8good_0/7good_0/6good_0/m1_14_20144# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R33 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R34 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R35 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X312 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X313 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X314 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X315 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X316 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X317 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X318 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X319 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X320 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X321 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X322 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X323 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X324 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X325 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X326 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X327 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X328 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X329 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X330 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X331 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X332 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X333 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X334 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X335 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R36 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R37 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R38 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R39 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X336 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X337 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X338 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X339 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X340 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X341 VDD D2 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X342 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X343 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X344 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X345 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X346 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X347 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X348 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X349 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X350 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X351 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X352 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X353 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X354 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X355 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X356 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X357 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X358 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X359 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X360 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X361 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X362 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X363 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X364 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X365 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X366 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X367 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R40 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R41 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R42 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R43 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X368 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X369 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X370 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X371 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X372 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X373 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X374 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X375 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X376 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X377 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X378 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X379 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X380 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X381 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X382 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X383 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X384 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X385 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X386 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X387 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X388 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X389 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X390 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X391 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R44 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R45 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R46 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R47 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X392 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X393 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X394 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X395 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X396 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X397 VDD D3 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X398 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X399 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X400 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X401 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X402 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X403 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X404 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X405 VDD D2 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X406 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X407 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X408 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X409 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X410 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X411 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X412 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X413 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X414 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X415 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X416 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X417 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X418 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X419 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X420 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X421 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X422 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X423 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X424 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X425 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X426 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X427 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X428 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X429 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X430 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X431 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R48 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R49 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R50 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R51 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X432 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X433 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X434 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X435 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X436 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X437 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X438 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X439 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X440 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X441 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X442 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X443 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X444 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X445 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X446 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X447 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X448 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X449 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X450 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X451 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X452 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X453 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X454 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X455 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R52 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R53 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R54 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R55 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X456 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X457 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X458 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X459 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X460 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X461 VDD D2 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X462 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X463 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X464 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X465 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X466 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X467 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X468 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X469 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X470 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X471 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X472 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X473 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X474 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X475 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X476 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X477 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X478 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X479 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X480 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X481 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X482 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X483 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X484 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X485 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X486 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X487 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R56 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R57 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R58 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R59 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X488 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X489 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X490 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X491 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X492 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X493 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X494 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X495 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X496 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X497 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X498 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X499 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X500 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X501 VDD D0 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X502 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X503 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X504 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X505 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X506 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X507 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X508 VDD 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X509 VDD D1 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X510 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X511 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R60 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R61 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R62 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# VREF sky130_fd_pr__res_generic_po1 w=66 l=342
R63 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X512 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X513 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/m1_8436_40544# 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X514 9good_0/8good_0/7good_0/m1_8436_40544# 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X515 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X516 VDD 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X517 VDD D5 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X518 9good_0/8good_0/7good_0/m1_8436_40544# 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 9good_0/8good_0/7good_0/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X519 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X520 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X521 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X522 9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X523 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X524 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X525 VDD D4 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X526 9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 9good_0/8good_0/7good_0/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X527 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X528 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X529 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X530 9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X531 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X532 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X533 VDD D3 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X534 9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X535 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X536 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X537 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X538 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X539 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X540 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X541 VDD D2 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X542 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X543 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X544 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X545 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X546 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X547 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X548 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X549 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X550 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X551 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X552 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X553 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X554 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_6754_8# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X555 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X556 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X557 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X558 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_6754_8# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X559 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X560 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X561 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X562 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X563 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X564 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X565 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X566 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X567 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R64 m1_6754_8# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R65 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R66 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R67 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X568 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X569 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X570 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X571 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X572 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X573 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X574 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X575 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X576 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X577 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X578 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X579 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X580 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X581 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X582 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X583 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X584 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X585 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X586 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X587 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X588 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X589 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X590 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X591 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R68 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R69 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R70 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R71 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X592 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X593 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X594 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X595 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X596 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X597 VDD D2 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X598 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X599 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X600 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X601 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X602 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X603 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X604 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X605 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X606 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X607 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X608 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X609 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X610 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X611 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X612 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X613 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X614 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X615 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X616 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X617 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X618 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X619 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X620 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X621 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X622 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X623 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R72 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R73 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R74 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R75 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X624 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X625 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X626 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X627 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X628 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X629 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X630 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X631 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X632 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X633 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X634 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X635 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X636 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X637 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X638 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X639 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X640 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X641 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X642 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X643 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X644 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X645 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X646 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X647 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R76 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R77 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R78 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R79 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X648 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X649 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X650 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X651 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X652 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X653 VDD D3 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X654 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X655 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X656 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X657 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X658 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X659 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X660 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X661 VDD D2 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X662 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X663 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X664 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X665 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X666 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X667 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X668 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X669 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X670 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X671 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X672 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X673 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X674 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X675 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X676 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X677 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X678 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X679 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X680 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X681 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X682 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X683 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X684 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X685 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X686 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X687 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R80 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R81 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R82 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R83 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X688 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X689 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X690 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X691 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X692 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X693 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X694 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X695 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X696 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X697 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X698 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X699 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X700 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X701 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X702 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X703 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X704 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X705 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X706 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X707 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X708 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X709 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X710 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X711 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R84 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R85 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R86 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R87 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X712 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X713 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X714 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X715 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X716 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X717 VDD D2 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X718 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X719 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X720 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X721 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X722 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X723 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X724 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X725 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X726 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X727 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X728 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X729 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X730 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X731 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X732 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X733 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X734 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X735 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X736 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X737 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X738 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X739 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X740 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X741 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X742 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X743 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R88 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R89 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R90 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R91 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X744 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X745 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X746 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X747 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X748 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X749 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X750 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X751 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X752 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X753 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X754 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X755 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X756 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X757 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X758 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X759 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X760 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X761 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X762 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X763 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X764 VDD 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X765 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X766 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X767 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R92 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R93 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R94 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R95 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X768 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X769 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X770 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X771 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X772 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X773 VDD D4 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X774 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X775 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X776 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X777 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X778 9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X779 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X780 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X781 VDD D3 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X782 9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X783 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X784 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X785 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X786 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X787 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X788 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X789 VDD D2 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X790 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X791 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X792 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X793 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X794 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X795 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X796 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X797 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X798 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X799 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X800 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X801 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X802 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X803 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X804 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X805 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X806 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/m1_14_20144# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X807 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X808 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X809 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X810 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X811 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X812 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X813 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X814 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X815 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R96 9good_0/8good_0/7good_0/6good_1/m1_14_20144# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R97 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R98 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R99 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X816 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X817 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X818 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X819 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X820 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X821 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X822 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X823 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X824 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X825 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X826 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X827 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X828 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X829 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X830 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X831 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X832 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X833 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X834 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X835 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X836 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X837 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X838 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X839 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R100 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R101 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R102 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R103 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X840 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X841 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X842 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X843 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X844 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X845 VDD D2 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X846 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X847 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X848 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X849 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X850 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X851 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X852 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X853 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X854 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X855 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X856 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X857 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X858 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X859 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X860 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X861 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X862 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X863 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X864 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X865 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X866 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X867 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X868 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X869 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X870 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X871 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R104 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R105 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R106 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R107 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X872 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X873 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X874 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X875 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X876 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X877 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X878 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X879 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X880 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X881 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X882 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X883 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X884 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X885 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X886 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X887 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X888 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X889 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X890 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X891 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X892 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X893 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X894 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X895 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R108 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R109 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R110 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R111 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X896 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X897 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X898 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X899 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X900 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X901 VDD D3 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X902 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X903 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X904 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X905 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X906 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X907 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X908 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X909 VDD D2 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X910 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X911 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X912 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X913 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X914 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X915 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X916 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X917 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X918 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X919 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X920 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X921 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X922 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X923 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X924 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X925 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X926 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X927 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X928 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X929 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X930 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X931 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X932 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X933 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X934 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X935 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R112 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R113 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R114 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R115 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X936 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X937 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X938 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X939 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X940 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X941 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X942 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X943 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X944 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X945 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X946 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X947 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X948 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X949 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X950 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X951 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X952 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X953 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X954 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X955 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X956 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X957 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X958 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X959 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R116 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R117 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R118 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R119 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X960 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X961 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X962 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X963 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X964 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X965 VDD D2 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X966 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X967 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X968 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X969 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X970 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X971 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X972 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X973 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X974 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X975 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X976 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X977 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X978 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X979 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X980 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X981 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X982 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X983 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X984 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X985 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X986 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X987 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X988 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X989 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X990 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X991 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R120 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R121 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R122 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R123 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X992 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X993 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X994 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X995 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X996 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X997 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X998 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X999 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1000 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1001 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1002 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1003 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1004 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1005 VDD D0 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1006 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1007 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1008 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1009 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1010 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1011 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1012 VDD 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1013 VDD D1 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1014 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1015 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R124 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R125 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R126 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_1684_72# sky130_fd_pr__res_generic_po1 w=66 l=342
R127 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1016 9good_0/8good_0/Sw-1_0/li_29_719# D7 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1017 9good_0/8good_0/m1_8774_43264# 9good_0/8good_0/Sw-1_0/li_29_719# 9good_0/m1_19068_42976# 9good_0/8good_0/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X1018 9good_0/m1_19068_42976# 9good_0/8good_0/Sw-1_0/li_29_719# 9good_0/8good_0/m1_18694_42308# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1019 9good_0/8good_0/Sw-1_0/li_126_470# 9good_0/8good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1020 VDD 9good_0/8good_0/Sw-1_0/li_29_719# 9good_0/8good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1021 VDD D7 9good_0/8good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1022 9good_0/m1_19068_42976# 9good_0/8good_0/Sw-1_0/li_126_470# 9good_0/8good_0/m1_18694_42308# 9good_0/m1_19068_42976# sky130_fd_pr__pfet_01v8 w=84 l=30
X1023 9good_0/8good_0/m1_8774_43264# 9good_0/8good_0/Sw-1_0/li_126_470# 9good_0/m1_19068_42976# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1024 9good_0/8good_0/7good_1/Sw-1_0/li_29_719# D6 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1025 9good_0/8good_0/7good_1/m1_4396_20620# 9good_0/8good_0/7good_1/Sw-1_0/li_29_719# 9good_0/8good_0/m1_18694_42308# 9good_0/8good_0/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X1026 9good_0/8good_0/m1_18694_42308# 9good_0/8good_0/7good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1027 9good_0/8good_0/7good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1028 VDD 9good_0/8good_0/7good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1029 VDD D6 9good_0/8good_0/7good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1030 9good_0/8good_0/m1_18694_42308# 9good_0/8good_0/7good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/m1_8436_40544# 9good_0/8good_0/m1_18694_42308# sky130_fd_pr__pfet_01v8 w=84 l=30
X1031 9good_0/8good_0/7good_1/m1_4396_20620# 9good_0/8good_0/7good_1/Sw-1_0/li_126_470# 9good_0/8good_0/m1_18694_42308# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1032 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1033 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/m1_4396_20620# 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X1034 9good_0/8good_0/7good_1/m1_4396_20620# 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1035 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1036 VDD 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1037 VDD D5 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1038 9good_0/8good_0/7good_1/m1_4396_20620# 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 9good_0/8good_0/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X1039 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/m1_4396_20620# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1040 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1041 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1042 9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1043 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1044 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1045 VDD D4 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1046 9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X1047 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1048 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1049 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1050 9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1051 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1052 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1053 VDD D3 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1054 9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X1055 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1056 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1057 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1058 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1059 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1060 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1061 VDD D2 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1062 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1063 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1064 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1065 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1066 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1067 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1068 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1069 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1070 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1071 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1072 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1073 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1074 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_11882_62# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1075 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1076 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1077 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1078 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_11882_62# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1079 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1080 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1081 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1082 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1083 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1084 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1085 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1086 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1087 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R128 m1_11882_62# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R129 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R130 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R131 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1088 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1089 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1090 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1091 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1092 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1093 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1094 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1095 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1096 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1097 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1098 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1099 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1100 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1101 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1102 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1103 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1104 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1105 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1106 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1107 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1108 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1109 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1110 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1111 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R132 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R133 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R134 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R135 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1112 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1113 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1114 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1115 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1116 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1117 VDD D2 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1118 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1119 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1120 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1121 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1122 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1123 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1124 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1125 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1126 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1127 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1128 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1129 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1130 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1131 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1132 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1133 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1134 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1135 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1136 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1137 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1138 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1139 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1140 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1141 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1142 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1143 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R136 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R137 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R138 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R139 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1144 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1145 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1146 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1147 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1148 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1149 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1150 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1151 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1152 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1153 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1154 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1155 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1156 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1157 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1158 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1159 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1160 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1161 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1162 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1163 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1164 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1165 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1166 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1167 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R140 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R141 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R142 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R143 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1168 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1169 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1170 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1171 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1172 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1173 VDD D3 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1174 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1175 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1176 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1177 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1178 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1179 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1180 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1181 VDD D2 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1182 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1183 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1184 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1185 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1186 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1187 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1188 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1189 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1190 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1191 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1192 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1193 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1194 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1195 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1196 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1197 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1198 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1199 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1200 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1201 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1202 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1203 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1204 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1205 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1206 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1207 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R144 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R145 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R146 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R147 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1208 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1209 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1210 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1211 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1212 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1213 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1214 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1215 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1216 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1217 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1218 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1219 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1220 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1221 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1222 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1223 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1224 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1225 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1226 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1227 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1228 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1229 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1230 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1231 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R148 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R149 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R150 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R151 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1232 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1233 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1234 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1235 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1236 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1237 VDD D2 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1238 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1239 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1240 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1241 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1242 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1243 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1244 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1245 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1246 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1247 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1248 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1249 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1250 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1251 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1252 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1253 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1254 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1255 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1256 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1257 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1258 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1259 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1260 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1261 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1262 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1263 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R152 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R153 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R154 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R155 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1264 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1265 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1266 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1267 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1268 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1269 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1270 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1271 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1272 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1273 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1274 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1275 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1276 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1277 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1278 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1279 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1280 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1281 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1282 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1283 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1284 VDD 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1285 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1286 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1287 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R156 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R157 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R158 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R159 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1288 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1289 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1290 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1291 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1292 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1293 VDD D4 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1294 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X1295 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1296 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1297 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1298 9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1299 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1300 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1301 VDD D3 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1302 9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X1303 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1304 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1305 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1306 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1307 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1308 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1309 VDD D2 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1310 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1311 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1312 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1313 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1314 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1315 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1316 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1317 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1318 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1319 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1320 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1321 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1322 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1323 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1324 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1325 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1326 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/m1_14_20144# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1327 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1328 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1329 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1330 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1331 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1332 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1333 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1334 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1335 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R160 9good_0/8good_0/7good_1/6good_0/m1_14_20144# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R161 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R162 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R163 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1336 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1337 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1338 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1339 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1340 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1341 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1342 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1343 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1344 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1345 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1346 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1347 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1348 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1349 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1350 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1351 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1352 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1353 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1354 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1355 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1356 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1357 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1358 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1359 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R164 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R165 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R166 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R167 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1360 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1361 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1362 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1363 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1364 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1365 VDD D2 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1366 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1367 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1368 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1369 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1370 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1371 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1372 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1373 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1374 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1375 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1376 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1377 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1378 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1379 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1380 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1381 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1382 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1383 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1384 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1385 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1386 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1387 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1388 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1389 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1390 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1391 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R168 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R169 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R170 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R171 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1392 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1393 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1394 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1395 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1396 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1397 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1398 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1399 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1400 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1401 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1402 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1403 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1404 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1405 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1406 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1407 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1408 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1409 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1410 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1411 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1412 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1413 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1414 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1415 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R172 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R173 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R174 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R175 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1416 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1417 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1418 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1419 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1420 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1421 VDD D3 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1422 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1423 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1424 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1425 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1426 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1427 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1428 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1429 VDD D2 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1430 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1431 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1432 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1433 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1434 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1435 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1436 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1437 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1438 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1439 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1440 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1441 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1442 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1443 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1444 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1445 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1446 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1447 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1448 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1449 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1450 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1451 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1452 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1453 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1454 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1455 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R176 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R177 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R178 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R179 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1456 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1457 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1458 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1459 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1460 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1461 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1462 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1463 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1464 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1465 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1466 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1467 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1468 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1469 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1470 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1471 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1472 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1473 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1474 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1475 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1476 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1477 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1478 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1479 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R180 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R181 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R182 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R183 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1480 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1481 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1482 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1483 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1484 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1485 VDD D2 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1486 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1487 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1488 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1489 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1490 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1491 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1492 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1493 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1494 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1495 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1496 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1497 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1498 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1499 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1500 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1501 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1502 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1503 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1504 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1505 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1506 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1507 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1508 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1509 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1510 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1511 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R184 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R185 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R186 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R187 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1512 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1513 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1514 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1515 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1516 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1517 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1518 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1519 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1520 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1521 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1522 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1523 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1524 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1525 VDD D0 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1526 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1527 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1528 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1529 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1530 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1531 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1532 VDD 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1533 VDD D1 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1534 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1535 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R188 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R189 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R190 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_6754_8# sky130_fd_pr__res_generic_po1 w=66 l=342
R191 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1536 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1537 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/m1_8436_40544# 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X1538 9good_0/8good_0/7good_1/m1_8436_40544# 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1539 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1540 VDD 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1541 VDD D5 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1542 9good_0/8good_0/7good_1/m1_8436_40544# 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 9good_0/8good_0/7good_1/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X1543 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1544 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1545 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1546 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1547 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1548 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1549 VDD D4 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1550 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X1551 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1552 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1553 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1554 9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1555 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1556 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1557 VDD D3 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1558 9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X1559 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1560 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1561 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1562 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1563 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1564 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1565 VDD D2 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1566 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1567 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1568 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1569 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1570 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1571 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1572 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1573 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1574 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1575 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1576 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1577 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1578 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_16966_2# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1579 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1580 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1581 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1582 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_16966_2# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1583 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1584 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1585 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1586 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1587 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1588 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1589 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1590 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1591 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R192 m1_16966_2# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R193 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R194 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R195 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1592 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1593 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1594 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1595 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1596 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1597 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1598 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1599 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1600 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1601 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1602 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1603 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1604 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1605 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1606 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1607 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1608 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1609 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1610 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1611 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1612 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1613 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1614 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1615 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R196 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R197 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R198 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R199 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1616 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1617 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1618 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1619 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1620 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1621 VDD D2 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1622 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1623 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1624 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1625 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1626 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1627 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1628 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1629 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1630 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1631 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1632 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1633 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1634 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1635 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1636 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1637 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1638 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1639 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1640 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1641 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1642 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1643 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1644 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1645 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1646 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1647 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R200 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R201 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R202 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R203 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1648 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1649 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1650 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1651 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1652 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1653 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1654 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1655 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1656 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1657 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1658 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1659 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1660 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1661 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1662 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1663 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1664 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1665 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1666 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1667 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1668 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1669 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1670 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1671 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R204 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R205 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R206 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R207 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1672 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1673 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1674 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1675 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1676 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1677 VDD D3 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1678 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1679 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1680 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1681 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1682 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1683 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1684 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1685 VDD D2 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1686 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1687 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1688 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1689 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1690 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1691 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1692 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1693 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1694 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1695 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1696 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1697 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1698 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1699 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1700 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1701 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1702 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1703 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1704 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1705 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1706 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1707 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1708 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1709 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1710 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1711 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R208 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R209 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R210 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R211 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1712 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1713 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1714 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1715 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1716 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1717 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1718 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1719 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1720 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1721 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1722 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1723 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1724 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1725 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1726 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1727 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1728 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1729 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1730 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1731 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1732 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1733 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1734 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1735 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R212 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R213 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R214 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R215 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1736 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1737 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1738 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1739 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1740 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1741 VDD D2 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1742 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1743 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1744 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1745 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1746 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1747 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1748 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1749 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1750 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1751 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1752 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1753 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1754 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1755 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1756 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1757 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1758 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1759 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1760 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1761 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1762 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1763 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1764 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1765 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1766 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1767 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R216 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R217 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R218 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R219 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1768 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1769 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1770 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1771 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1772 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1773 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1774 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1775 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1776 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1777 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1778 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1779 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1780 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1781 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1782 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1783 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1784 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1785 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1786 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1787 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1788 VDD 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1789 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1790 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1791 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R220 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R221 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R222 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R223 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1792 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1793 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1794 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1795 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1796 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1797 VDD D4 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1798 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X1799 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1800 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1801 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1802 9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1803 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1804 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1805 VDD D3 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1806 9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X1807 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1808 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1809 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1810 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1811 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1812 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1813 VDD D2 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1814 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1815 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1816 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1817 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1818 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1819 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1820 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1821 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1822 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1823 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1824 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1825 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1826 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1827 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1828 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1829 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1830 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/m1_14_20144# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1831 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1832 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1833 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1834 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1835 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1836 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1837 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1838 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1839 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R224 9good_0/8good_0/7good_1/6good_1/m1_14_20144# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R225 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R226 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R227 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1840 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1841 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1842 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1843 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1844 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1845 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1846 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1847 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1848 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1849 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1850 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1851 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1852 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1853 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1854 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1855 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1856 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1857 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1858 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1859 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1860 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1861 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1862 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1863 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R228 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R229 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R230 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R231 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1864 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1865 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1866 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1867 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1868 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1869 VDD D2 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1870 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1871 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1872 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1873 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1874 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1875 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1876 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1877 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1878 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1879 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1880 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1881 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1882 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1883 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1884 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1885 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1886 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1887 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1888 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1889 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1890 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1891 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1892 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1893 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1894 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1895 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R232 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R233 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R234 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R235 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1896 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1897 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1898 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1899 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1900 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1901 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1902 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1903 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1904 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1905 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1906 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1907 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1908 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1909 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1910 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1911 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1912 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1913 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1914 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1915 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1916 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1917 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1918 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1919 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R236 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R237 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R238 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R239 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1920 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1921 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1922 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1923 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1924 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1925 VDD D3 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1926 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1927 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1928 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1929 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1930 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1931 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1932 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1933 VDD D2 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1934 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1935 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1936 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1937 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1938 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1939 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1940 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1941 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1942 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1943 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1944 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1945 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1946 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1947 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1948 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1949 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1950 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1951 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1952 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1953 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1954 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1955 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1956 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1957 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1958 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1959 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R240 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R241 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R242 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R243 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1960 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1961 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1962 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1963 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1964 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1965 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1966 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1967 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1968 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1969 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1970 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1971 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1972 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1973 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1974 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1975 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1976 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1977 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1978 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1979 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1980 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1981 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1982 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1983 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R244 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R245 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R246 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R247 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X1984 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1985 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1986 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1987 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1988 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1989 VDD D2 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1990 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1991 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1992 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1993 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1994 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1995 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X1996 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1997 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X1998 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1999 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2000 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2001 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2002 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2003 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2004 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2005 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2006 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2007 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2008 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2009 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2010 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2011 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2012 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2013 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2014 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2015 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R248 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R249 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R250 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R251 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2016 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2017 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2018 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2019 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2020 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2021 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2022 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2023 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2024 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2025 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2026 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2027 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2028 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2029 VDD D0 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2030 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2031 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2032 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2033 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2034 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2035 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2036 VDD 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2037 VDD D1 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2038 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2039 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R252 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R253 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R254 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_11882_62# sky130_fd_pr__res_generic_po1 w=66 l=342
R255 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2040 9good_0/8good_1/7good_0/Sw-1_0/li_29_719# D6 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2041 9good_0/8good_1/7good_0/m1_4396_20620# 9good_0/8good_1/7good_0/Sw-1_0/li_29_719# 9good_0/8good_1/m1_8774_43264# 9good_0/8good_1/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X2042 9good_0/8good_1/m1_8774_43264# 9good_0/8good_1/7good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2043 9good_0/8good_1/7good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2044 VDD 9good_0/8good_1/7good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2045 VDD D6 9good_0/8good_1/7good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2046 9good_0/8good_1/m1_8774_43264# 9good_0/8good_1/7good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/m1_8436_40544# 9good_0/8good_1/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X2047 9good_0/8good_1/7good_0/m1_4396_20620# 9good_0/8good_1/7good_0/Sw-1_0/li_126_470# 9good_0/8good_1/m1_8774_43264# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2048 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2049 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/m1_4396_20620# 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2050 9good_0/8good_1/7good_0/m1_4396_20620# 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2051 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2052 VDD 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2053 VDD D5 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2054 9good_0/8good_1/7good_0/m1_4396_20620# 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 9good_0/8good_1/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X2055 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/m1_4396_20620# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2056 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2057 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2058 9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2059 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2060 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2061 VDD D4 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2062 9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X2063 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2064 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2065 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2066 9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2067 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2068 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2069 VDD D3 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2070 9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X2071 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2072 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2073 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2074 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2075 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2076 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2077 VDD D2 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2078 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2079 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2080 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2081 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2082 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2083 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2084 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2085 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2086 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2087 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2088 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2089 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2090 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_21660_68# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2091 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2092 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2093 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2094 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_21660_68# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2095 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2096 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2097 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2098 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2099 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2100 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2101 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2102 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2103 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R256 m1_21660_68# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R257 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R258 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R259 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2104 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2105 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2106 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2107 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2108 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2109 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2110 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2111 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2112 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2113 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2114 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2115 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2116 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2117 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2118 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2119 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2120 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2121 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2122 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2123 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2124 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2125 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2126 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2127 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R260 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R261 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R262 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R263 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2128 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2129 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2130 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2131 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2132 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2133 VDD D2 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2134 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2135 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2136 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2137 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2138 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2139 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2140 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2141 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2142 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2143 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2144 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2145 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2146 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2147 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2148 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2149 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2150 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2151 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2152 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2153 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2154 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2155 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2156 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2157 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2158 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2159 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R264 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R265 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R266 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R267 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2160 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2161 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2162 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2163 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2164 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2165 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2166 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2167 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2168 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2169 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2170 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2171 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2172 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2173 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2174 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2175 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2176 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2177 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2178 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2179 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2180 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2181 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2182 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2183 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R268 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R269 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R270 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R271 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2184 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2185 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2186 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2187 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2188 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2189 VDD D3 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2190 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2191 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2192 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2193 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2194 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2195 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2196 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2197 VDD D2 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2198 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2199 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2200 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2201 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2202 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2203 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2204 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2205 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2206 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2207 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2208 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2209 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2210 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2211 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2212 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2213 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2214 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2215 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2216 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2217 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2218 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2219 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2220 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2221 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2222 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2223 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R272 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R273 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R274 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R275 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2224 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2225 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2226 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2227 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2228 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2229 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2230 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2231 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2232 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2233 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2234 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2235 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2236 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2237 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2238 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2239 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2240 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2241 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2242 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2243 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2244 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2245 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2246 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2247 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R276 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R277 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R278 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R279 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2248 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2249 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2250 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2251 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2252 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2253 VDD D2 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2254 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2255 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2256 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2257 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2258 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2259 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2260 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2261 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2262 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2263 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2264 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2265 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2266 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2267 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2268 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2269 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2270 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2271 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2272 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2273 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2274 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2275 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2276 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2277 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2278 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2279 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R280 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R281 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R282 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R283 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2280 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2281 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2282 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2283 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2284 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2285 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2286 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2287 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2288 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2289 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2290 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2291 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2292 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2293 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2294 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2295 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2296 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2297 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2298 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2299 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2300 VDD 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2301 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2302 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2303 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R284 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R285 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R286 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R287 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2304 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2305 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2306 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2307 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2308 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2309 VDD D4 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2310 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2311 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2312 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2313 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2314 9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2315 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2316 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2317 VDD D3 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2318 9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X2319 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2320 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2321 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2322 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2323 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2324 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2325 VDD D2 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2326 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2327 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2328 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2329 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2330 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2331 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2332 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2333 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2334 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2335 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2336 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2337 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2338 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2339 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2340 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2341 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2342 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/m1_14_20144# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2343 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2344 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2345 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2346 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2347 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2348 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2349 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2350 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2351 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R288 9good_0/8good_1/7good_0/6good_0/m1_14_20144# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R289 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R290 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R291 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2352 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2353 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2354 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2355 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2356 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2357 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2358 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2359 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2360 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2361 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2362 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2363 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2364 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2365 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2366 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2367 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2368 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2369 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2370 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2371 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2372 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2373 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2374 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2375 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R292 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R293 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R294 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R295 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2376 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2377 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2378 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2379 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2380 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2381 VDD D2 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2382 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2383 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2384 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2385 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2386 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2387 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2388 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2389 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2390 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2391 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2392 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2393 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2394 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2395 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2396 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2397 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2398 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2399 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2400 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2401 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2402 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2403 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2404 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2405 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2406 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2407 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R296 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R297 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R298 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R299 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2408 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2409 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2410 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2411 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2412 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2413 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2414 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2415 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2416 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2417 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2418 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2419 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2420 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2421 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2422 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2423 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2424 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2425 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2426 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2427 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2428 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2429 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2430 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2431 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R300 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R301 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R302 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R303 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2432 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2433 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2434 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2435 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2436 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2437 VDD D3 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2438 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2439 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2440 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2441 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2442 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2443 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2444 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2445 VDD D2 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2446 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2447 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2448 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2449 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2450 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2451 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2452 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2453 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2454 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2455 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2456 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2457 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2458 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2459 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2460 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2461 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2462 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2463 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2464 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2465 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2466 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2467 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2468 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2469 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2470 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2471 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R304 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R305 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R306 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R307 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2472 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2473 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2474 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2475 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2476 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2477 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2478 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2479 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2480 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2481 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2482 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2483 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2484 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2485 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2486 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2487 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2488 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2489 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2490 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2491 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2492 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2493 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2494 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2495 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R308 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R309 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R310 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R311 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2496 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2497 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2498 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2499 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2500 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2501 VDD D2 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2502 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2503 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2504 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2505 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2506 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2507 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2508 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2509 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2510 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2511 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2512 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2513 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2514 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2515 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2516 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2517 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2518 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2519 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2520 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2521 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2522 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2523 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2524 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2525 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2526 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2527 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R312 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R313 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R314 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R315 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2528 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2529 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2530 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2531 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2532 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2533 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2534 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2535 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2536 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2537 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2538 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2539 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2540 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2541 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2542 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2543 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2544 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2545 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2546 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2547 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2548 VDD 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2549 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2550 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2551 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R316 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R317 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R318 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_16966_2# sky130_fd_pr__res_generic_po1 w=66 l=342
R319 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2552 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2553 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/m1_8436_40544# 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2554 9good_0/8good_1/7good_0/m1_8436_40544# 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2555 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2556 VDD 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2557 VDD D5 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2558 9good_0/8good_1/7good_0/m1_8436_40544# 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 9good_0/8good_1/7good_0/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X2559 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2560 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2561 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2562 9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2563 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2564 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2565 VDD D4 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2566 9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X2567 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2568 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2569 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2570 9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2571 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2572 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2573 VDD D3 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2574 9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X2575 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2576 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2577 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2578 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2579 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2580 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2581 VDD D2 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2582 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2583 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2584 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2585 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2586 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2587 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2588 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2589 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2590 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2591 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2592 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2593 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2594 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_26760_28# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2595 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2596 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2597 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2598 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_26760_28# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2599 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2600 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2601 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2602 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2603 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2604 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2605 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2606 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2607 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R320 m1_26760_28# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R321 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R322 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R323 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2608 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2609 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2610 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2611 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2612 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2613 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2614 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2615 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2616 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2617 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2618 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2619 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2620 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2621 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2622 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2623 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2624 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2625 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2626 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2627 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2628 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2629 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2630 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2631 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R324 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R325 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R326 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R327 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2632 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2633 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2634 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2635 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2636 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2637 VDD D2 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2638 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2639 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2640 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2641 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2642 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2643 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2644 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2645 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2646 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2647 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2648 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2649 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2650 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2651 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2652 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2653 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2654 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2655 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2656 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2657 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2658 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2659 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2660 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2661 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2662 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2663 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R328 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R329 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R330 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R331 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2664 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2665 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2666 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2667 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2668 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2669 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2670 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2671 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2672 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2673 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2674 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2675 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2676 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2677 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2678 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2679 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2680 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2681 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2682 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2683 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2684 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2685 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2686 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2687 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R332 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R333 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R334 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R335 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2688 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2689 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2690 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2691 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2692 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2693 VDD D3 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2694 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2695 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2696 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2697 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2698 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2699 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2700 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2701 VDD D2 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2702 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2703 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2704 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2705 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2706 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2707 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2708 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2709 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2710 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2711 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2712 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2713 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2714 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2715 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2716 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2717 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2718 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2719 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2720 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2721 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2722 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2723 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2724 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2725 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2726 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2727 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R336 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R337 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R338 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R339 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2728 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2729 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2730 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2731 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2732 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2733 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2734 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2735 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2736 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2737 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2738 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2739 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2740 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2741 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2742 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2743 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2744 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2745 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2746 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2747 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2748 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2749 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2750 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2751 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R340 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R341 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R342 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R343 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2752 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2753 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2754 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2755 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2756 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2757 VDD D2 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2758 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2759 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2760 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2761 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2762 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2763 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2764 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2765 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2766 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2767 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2768 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2769 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2770 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2771 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2772 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2773 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2774 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2775 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2776 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2777 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2778 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2779 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2780 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2781 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2782 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2783 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R344 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R345 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R346 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R347 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2784 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2785 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2786 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2787 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2788 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2789 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2790 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2791 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2792 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2793 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2794 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2795 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2796 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2797 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2798 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2799 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2800 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2801 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2802 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2803 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2804 VDD 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2805 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2806 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2807 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R348 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R349 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R350 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R351 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2808 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2809 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2810 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2811 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2812 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2813 VDD D4 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2814 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2815 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2816 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2817 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2818 9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2819 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2820 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2821 VDD D3 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2822 9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X2823 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2824 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2825 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2826 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2827 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2828 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2829 VDD D2 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2830 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2831 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2832 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2833 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2834 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2835 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2836 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2837 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2838 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2839 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2840 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2841 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2842 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2843 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2844 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2845 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2846 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/m1_14_20144# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2847 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2848 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2849 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2850 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2851 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2852 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2853 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2854 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2855 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R352 9good_0/8good_1/7good_0/6good_1/m1_14_20144# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R353 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R354 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R355 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2856 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2857 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2858 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2859 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2860 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2861 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2862 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2863 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2864 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2865 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2866 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2867 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2868 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2869 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2870 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2871 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2872 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2873 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2874 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2875 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2876 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2877 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2878 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2879 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R356 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R357 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R358 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R359 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2880 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2881 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2882 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2883 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2884 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2885 VDD D2 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2886 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2887 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2888 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2889 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2890 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2891 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2892 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2893 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2894 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2895 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2896 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2897 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2898 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2899 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2900 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2901 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2902 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2903 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2904 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2905 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2906 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2907 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2908 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2909 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2910 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2911 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R360 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R361 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R362 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R363 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2912 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2913 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2914 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2915 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2916 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2917 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2918 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2919 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2920 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2921 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2922 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2923 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2924 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2925 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2926 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2927 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2928 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2929 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2930 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2931 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2932 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2933 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2934 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2935 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R364 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R365 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R366 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R367 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2936 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2937 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2938 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2939 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2940 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2941 VDD D3 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2942 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2943 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2944 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2945 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2946 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2947 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2948 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2949 VDD D2 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2950 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2951 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2952 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2953 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2954 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2955 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2956 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2957 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2958 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2959 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2960 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2961 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2962 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2963 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2964 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2965 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2966 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2967 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2968 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2969 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2970 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2971 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2972 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2973 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2974 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2975 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R368 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R369 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R370 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R371 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X2976 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2977 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2978 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2979 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2980 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2981 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2982 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2983 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2984 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2985 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2986 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2987 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2988 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2989 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2990 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2991 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2992 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2993 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2994 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2995 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X2996 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2997 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X2998 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2999 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R372 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R373 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R374 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R375 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3000 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3001 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3002 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3003 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3004 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3005 VDD D2 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3006 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3007 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3008 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3009 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3010 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3011 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3012 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3013 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3014 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3015 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3016 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3017 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3018 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3019 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3020 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3021 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3022 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3023 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3024 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3025 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3026 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3027 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3028 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3029 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3030 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3031 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R376 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R377 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R378 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R379 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3032 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3033 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3034 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3035 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3036 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3037 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3038 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3039 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3040 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3041 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3042 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3043 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3044 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3045 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3046 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3047 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3048 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3049 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3050 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3051 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3052 VDD 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3053 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3054 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3055 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R380 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R381 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R382 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_21660_68# sky130_fd_pr__res_generic_po1 w=66 l=342
R383 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3056 9good_0/8good_1/Sw-1_0/li_29_719# D7 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3057 9good_0/8good_1/m1_8774_43264# 9good_0/8good_1/Sw-1_0/li_29_719# 9good_0/m1_38716_44140# 9good_0/8good_1/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X3058 9good_0/m1_38716_44140# 9good_0/8good_1/Sw-1_0/li_29_719# 9good_0/8good_1/m1_18694_42308# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3059 9good_0/8good_1/Sw-1_0/li_126_470# 9good_0/8good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3060 VDD 9good_0/8good_1/Sw-1_0/li_29_719# 9good_0/8good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3061 VDD D7 9good_0/8good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3062 9good_0/m1_38716_44140# 9good_0/8good_1/Sw-1_0/li_126_470# 9good_0/8good_1/m1_18694_42308# 9good_0/m1_38716_44140# sky130_fd_pr__pfet_01v8 w=84 l=30
X3063 9good_0/8good_1/m1_8774_43264# 9good_0/8good_1/Sw-1_0/li_126_470# 9good_0/m1_38716_44140# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3064 9good_0/8good_1/7good_1/Sw-1_0/li_29_719# D6 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3065 9good_0/8good_1/7good_1/m1_4396_20620# 9good_0/8good_1/7good_1/Sw-1_0/li_29_719# 9good_0/8good_1/m1_18694_42308# 9good_0/8good_1/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X3066 9good_0/8good_1/m1_18694_42308# 9good_0/8good_1/7good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3067 9good_0/8good_1/7good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3068 VDD 9good_0/8good_1/7good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3069 VDD D6 9good_0/8good_1/7good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3070 9good_0/8good_1/m1_18694_42308# 9good_0/8good_1/7good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/m1_8436_40544# 9good_0/8good_1/m1_18694_42308# sky130_fd_pr__pfet_01v8 w=84 l=30
X3071 9good_0/8good_1/7good_1/m1_4396_20620# 9good_0/8good_1/7good_1/Sw-1_0/li_126_470# 9good_0/8good_1/m1_18694_42308# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3072 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3073 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/m1_4396_20620# 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X3074 9good_0/8good_1/7good_1/m1_4396_20620# 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3075 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3076 VDD 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3077 VDD D5 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3078 9good_0/8good_1/7good_1/m1_4396_20620# 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 9good_0/8good_1/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X3079 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/m1_4396_20620# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3080 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3081 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3082 9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3083 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3084 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3085 VDD D4 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3086 9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 9good_0/8good_1/7good_1/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X3087 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3088 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3089 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3090 9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3091 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3092 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3093 VDD D3 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3094 9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X3095 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3096 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3097 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3098 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3099 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3100 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3101 VDD D2 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3102 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3103 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3104 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3105 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3106 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3107 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3108 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3109 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3110 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3111 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3112 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3113 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3114 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_31884_48# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3115 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3116 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3117 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3118 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_31884_48# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3119 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3120 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3121 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3122 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3123 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3124 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3125 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3126 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3127 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R384 m1_31884_48# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R385 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R386 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R387 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3128 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3129 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3130 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3131 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3132 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3133 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3134 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3135 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3136 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3137 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3138 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3139 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3140 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3141 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3142 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3143 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3144 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3145 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3146 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3147 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3148 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3149 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3150 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3151 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R388 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R389 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R390 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R391 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3152 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3153 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3154 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3155 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3156 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3157 VDD D2 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3158 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3159 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3160 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3161 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3162 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3163 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3164 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3165 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3166 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3167 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3168 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3169 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3170 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3171 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3172 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3173 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3174 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3175 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3176 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3177 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3178 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3179 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3180 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3181 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3182 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3183 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R392 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R393 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R394 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R395 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3184 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3185 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3186 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3187 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3188 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3189 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3190 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3191 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3192 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3193 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3194 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3195 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3196 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3197 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3198 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3199 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3200 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3201 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3202 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3203 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3204 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3205 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3206 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3207 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R396 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R397 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R398 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R399 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3208 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3209 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3210 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3211 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3212 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3213 VDD D3 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3214 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3215 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3216 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3217 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3218 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3219 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3220 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3221 VDD D2 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3222 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3223 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3224 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3225 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3226 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3227 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3228 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3229 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3230 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3231 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3232 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3233 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3234 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3235 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3236 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3237 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3238 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3239 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3240 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3241 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3242 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3243 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3244 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3245 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3246 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3247 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R400 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R401 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R402 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R403 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3248 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3249 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3250 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3251 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3252 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3253 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3254 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3255 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3256 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3257 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3258 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3259 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3260 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3261 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3262 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3263 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3264 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3265 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3266 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3267 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3268 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3269 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3270 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3271 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R404 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R405 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R406 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R407 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3272 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3273 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3274 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3275 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3276 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3277 VDD D2 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3278 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3279 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3280 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3281 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3282 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3283 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3284 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3285 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3286 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3287 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3288 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3289 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3290 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3291 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3292 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3293 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3294 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3295 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3296 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3297 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3298 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3299 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3300 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3301 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3302 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3303 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R408 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R409 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R410 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R411 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3304 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3305 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3306 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3307 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3308 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3309 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3310 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3311 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3312 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3313 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3314 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3315 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3316 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3317 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3318 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3319 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3320 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3321 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3322 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3323 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3324 VDD 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3325 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3326 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3327 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R412 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R413 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R414 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R415 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3328 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3329 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3330 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3331 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3332 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3333 VDD D4 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3334 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X3335 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3336 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3337 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3338 9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3339 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3340 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3341 VDD D3 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3342 9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X3343 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3344 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3345 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3346 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3347 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3348 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3349 VDD D2 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3350 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3351 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3352 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3353 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3354 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3355 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3356 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3357 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3358 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3359 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3360 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3361 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3362 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3363 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3364 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3365 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3366 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/m1_14_20144# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3367 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3368 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3369 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3370 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3371 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3372 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3373 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3374 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3375 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R416 9good_0/8good_1/7good_1/6good_0/m1_14_20144# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R417 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R418 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R419 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3376 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3377 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3378 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3379 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3380 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3381 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3382 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3383 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3384 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3385 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3386 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3387 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3388 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3389 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3390 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3391 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3392 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3393 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3394 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3395 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3396 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3397 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3398 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3399 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R420 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R421 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R422 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R423 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3400 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3401 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3402 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3403 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3404 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3405 VDD D2 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3406 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3407 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3408 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3409 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3410 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3411 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3412 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3413 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3414 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3415 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3416 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3417 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3418 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3419 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3420 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3421 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3422 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3423 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3424 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3425 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3426 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3427 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3428 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3429 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3430 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3431 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R424 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R425 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R426 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R427 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3432 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3433 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3434 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3435 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3436 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3437 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3438 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3439 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3440 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3441 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3442 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3443 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3444 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3445 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3446 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3447 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3448 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3449 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3450 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3451 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3452 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3453 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3454 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3455 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R428 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R429 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R430 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R431 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3456 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3457 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3458 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3459 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3460 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3461 VDD D3 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3462 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3463 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3464 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3465 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3466 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3467 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3468 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3469 VDD D2 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3470 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3471 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3472 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3473 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3474 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3475 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3476 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3477 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3478 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3479 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3480 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3481 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3482 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3483 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3484 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3485 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3486 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3487 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3488 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3489 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3490 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3491 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3492 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3493 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3494 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3495 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R432 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R433 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R434 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R435 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3496 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3497 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3498 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3499 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3500 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3501 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3502 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3503 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3504 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3505 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3506 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3507 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3508 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3509 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3510 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3511 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3512 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3513 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3514 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3515 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3516 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3517 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3518 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3519 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R436 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R437 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R438 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R439 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3520 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3521 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3522 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3523 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3524 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3525 VDD D2 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3526 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3527 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3528 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3529 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3530 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3531 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3532 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3533 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3534 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3535 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3536 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3537 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3538 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3539 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3540 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3541 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3542 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3543 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3544 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3545 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3546 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3547 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3548 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3549 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3550 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3551 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R440 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R441 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R442 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R443 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3552 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3553 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3554 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3555 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3556 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3557 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3558 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3559 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3560 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3561 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3562 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3563 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3564 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3565 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3566 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3567 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3568 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3569 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3570 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3571 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3572 VDD 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3573 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3574 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3575 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R444 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R445 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R446 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_26760_28# sky130_fd_pr__res_generic_po1 w=66 l=342
R447 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3576 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3577 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/m1_8436_40544# 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X3578 9good_0/8good_1/7good_1/m1_8436_40544# 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3579 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3580 VDD 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3581 VDD D5 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3582 9good_0/8good_1/7good_1/m1_8436_40544# 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 9good_0/8good_1/7good_1/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X3583 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3584 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3585 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3586 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3587 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3588 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3589 VDD D4 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3590 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X3591 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3592 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3593 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3594 9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3595 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3596 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3597 VDD D3 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3598 9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X3599 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3600 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3601 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3602 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3603 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3604 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3605 VDD D2 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3606 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3607 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3608 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3609 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3610 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3611 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3612 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3613 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3614 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3615 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3616 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3617 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3618 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_36912_2# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3619 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3620 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3621 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3622 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_36912_2# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3623 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3624 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3625 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3626 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3627 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3628 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3629 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3630 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3631 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R448 m1_36912_2# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R449 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R450 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R451 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3632 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3633 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3634 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3635 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3636 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3637 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3638 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3639 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3640 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3641 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3642 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3643 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3644 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3645 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3646 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3647 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3648 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3649 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3650 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3651 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3652 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3653 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3654 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3655 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R452 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R453 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R454 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R455 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3656 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3657 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3658 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3659 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3660 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3661 VDD D2 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3662 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3663 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3664 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3665 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3666 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3667 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3668 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3669 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3670 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3671 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3672 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3673 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3674 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3675 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3676 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3677 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3678 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3679 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3680 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3681 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3682 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3683 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3684 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3685 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3686 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3687 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R456 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R457 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R458 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R459 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3688 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3689 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3690 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3691 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3692 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3693 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3694 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3695 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3696 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3697 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3698 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3699 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3700 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3701 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3702 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3703 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3704 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3705 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3706 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3707 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3708 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3709 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3710 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3711 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R460 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R461 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R462 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R463 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3712 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3713 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3714 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3715 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3716 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3717 VDD D3 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3718 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3719 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3720 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3721 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3722 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3723 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3724 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3725 VDD D2 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3726 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3727 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3728 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3729 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3730 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3731 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3732 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3733 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3734 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3735 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3736 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3737 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3738 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3739 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3740 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3741 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3742 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3743 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3744 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3745 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3746 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3747 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3748 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3749 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3750 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3751 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R464 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R465 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R466 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R467 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3752 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3753 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3754 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3755 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3756 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3757 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3758 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3759 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3760 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3761 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3762 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3763 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3764 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3765 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3766 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3767 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3768 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3769 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3770 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3771 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3772 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3773 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3774 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3775 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R468 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R469 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R470 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R471 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3776 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3777 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3778 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3779 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3780 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3781 VDD D2 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3782 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3783 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3784 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3785 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3786 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3787 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3788 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3789 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3790 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3791 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3792 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3793 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3794 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3795 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3796 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3797 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3798 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3799 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3800 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3801 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3802 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3803 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3804 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3805 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3806 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3807 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R472 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R473 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R474 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R475 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3808 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3809 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3810 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3811 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3812 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3813 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3814 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3815 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3816 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3817 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3818 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3819 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3820 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3821 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3822 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3823 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3824 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3825 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3826 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3827 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3828 VDD 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3829 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3830 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3831 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R476 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R477 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R478 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R479 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3832 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3833 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3834 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3835 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3836 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3837 VDD D4 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3838 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X3839 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3840 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3841 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3842 9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3843 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3844 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3845 VDD D3 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3846 9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X3847 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3848 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3849 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3850 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3851 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3852 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3853 VDD D2 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3854 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3855 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3856 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3857 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3858 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3859 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3860 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3861 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3862 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3863 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3864 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3865 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3866 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3867 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3868 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3869 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3870 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/m1_14_20144# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3871 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3872 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3873 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3874 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3875 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3876 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3877 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3878 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3879 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R480 9good_0/8good_1/7good_1/6good_1/m1_14_20144# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R481 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R482 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R483 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3880 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3881 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3882 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3883 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3884 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3885 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3886 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3887 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3888 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3889 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3890 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3891 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3892 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3893 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3894 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3895 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3896 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3897 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3898 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3899 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3900 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3901 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3902 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3903 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R484 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R485 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R486 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R487 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3904 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3905 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3906 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3907 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3908 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3909 VDD D2 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3910 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3911 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3912 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3913 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3914 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3915 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3916 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3917 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3918 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3919 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3920 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3921 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3922 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3923 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3924 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3925 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3926 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3927 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3928 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3929 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3930 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3931 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3932 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3933 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3934 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3935 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R488 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R489 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R490 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R491 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3936 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3937 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3938 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3939 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3940 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3941 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3942 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3943 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3944 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3945 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3946 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3947 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3948 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3949 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3950 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3951 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3952 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3953 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3954 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3955 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3956 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3957 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3958 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3959 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R492 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R493 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R494 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R495 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X3960 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3961 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3962 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3963 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3964 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3965 VDD D3 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3966 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3967 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3968 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3969 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3970 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3971 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3972 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3973 VDD D2 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3974 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3975 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3976 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3977 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3978 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3979 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3980 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3981 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3982 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3983 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3984 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3985 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3986 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3987 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3988 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3989 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3990 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3991 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3992 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3993 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3994 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3995 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X3996 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3997 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X3998 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3999 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R496 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R497 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R498 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R499 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4000 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4001 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4002 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4003 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4004 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4005 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4006 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4007 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4008 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4009 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4010 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4011 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4012 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4013 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4014 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4015 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4016 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4017 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4018 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4019 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4020 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4021 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4022 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4023 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R500 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R501 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R502 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R503 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4024 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4025 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4026 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4027 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4028 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4029 VDD D2 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4030 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4031 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4032 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4033 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4034 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4035 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4036 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4037 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4038 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4039 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4040 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4041 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4042 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4043 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4044 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4045 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4046 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4047 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4048 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4049 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4050 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4051 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4052 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4053 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4054 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4055 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R504 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R505 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R506 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R507 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4056 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4057 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4058 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4059 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4060 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4061 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4062 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4063 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4064 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4065 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4066 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4067 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4068 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4069 VDD 9good_0/m1_32342_44672# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4070 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4071 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4072 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4073 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4074 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4075 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4076 VDD 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4077 VDD 9good_0/m1_32720_44664# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4078 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4079 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R508 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R509 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R510 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_31884_48# sky130_fd_pr__res_generic_po1 w=66 l=342
R511 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4080 9good_0/Sw-1_0/li_29_719# D8 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4081 9good_0/m1_19068_42976# 9good_0/Sw-1_0/li_29_719# m1_39076_44800# 9good_0/m1_19068_42976# sky130_fd_pr__pfet_01v8 w=84 l=30
X4082 m1_39076_44800# 9good_0/Sw-1_0/li_29_719# 9good_0/m1_38716_44140# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4083 9good_0/Sw-1_0/li_126_470# 9good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4084 VDD 9good_0/Sw-1_0/li_29_719# 9good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4085 VDD D8 9good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4086 m1_39076_44800# 9good_0/Sw-1_0/li_126_470# 9good_0/m1_38716_44140# m1_39076_44800# sky130_fd_pr__pfet_01v8 w=84 l=30
X4087 9good_0/m1_19068_42976# 9good_0/Sw-1_0/li_126_470# m1_39076_44800# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4088 9good_1/8good_0/7good_0/Sw-1_0/li_29_719# D6 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4089 9good_1/8good_0/7good_0/m1_4396_20620# 9good_1/8good_0/7good_0/Sw-1_0/li_29_719# 9good_1/8good_0/m1_8774_43264# 9good_1/8good_0/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X4090 9good_1/8good_0/m1_8774_43264# 9good_1/8good_0/7good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4091 9good_1/8good_0/7good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4092 VDD 9good_1/8good_0/7good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4093 VDD D6 9good_1/8good_0/7good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4094 9good_1/8good_0/m1_8774_43264# 9good_1/8good_0/7good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/m1_8436_40544# 9good_1/8good_0/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X4095 9good_1/8good_0/7good_0/m1_4396_20620# 9good_1/8good_0/7good_0/Sw-1_0/li_126_470# 9good_1/8good_0/m1_8774_43264# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4096 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4097 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/m1_4396_20620# 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X4098 9good_1/8good_0/7good_0/m1_4396_20620# 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4099 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4100 VDD 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4101 VDD D5 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4102 9good_1/8good_0/7good_0/m1_4396_20620# 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 9good_1/8good_0/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X4103 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/m1_4396_20620# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4104 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4105 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4106 9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4107 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4108 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4109 VDD D4 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4110 9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 9good_1/8good_0/7good_0/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X4111 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4112 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4113 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4114 9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4115 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4116 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4117 VDD D3 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4118 9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X4119 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4120 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4121 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4122 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4123 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4124 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4125 VDD D2 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4126 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4127 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4128 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4129 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4130 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4131 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4132 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4133 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4134 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4135 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4136 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4137 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4138 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_41532_78# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4139 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4140 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4141 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4142 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_41532_78# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4143 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4144 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4145 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4146 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4147 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4148 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4149 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4150 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4151 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R512 m1_41532_78# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R513 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R514 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R515 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4152 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4153 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4154 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4155 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4156 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4157 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4158 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4159 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4160 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4161 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4162 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4163 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4164 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4165 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4166 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4167 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4168 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4169 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4170 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4171 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4172 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4173 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4174 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4175 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R516 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R517 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R518 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R519 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4176 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4177 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4178 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4179 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4180 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4181 VDD D2 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4182 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4183 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4184 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4185 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4186 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4187 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4188 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4189 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4190 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4191 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4192 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4193 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4194 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4195 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4196 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4197 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4198 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4199 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4200 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4201 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4202 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4203 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4204 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4205 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4206 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4207 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R520 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R521 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R522 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R523 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4208 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4209 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4210 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4211 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4212 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4213 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4214 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4215 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4216 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4217 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4218 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4219 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4220 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4221 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4222 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4223 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4224 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4225 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4226 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4227 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4228 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4229 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4230 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4231 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R524 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R525 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R526 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R527 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4232 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4233 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4234 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4235 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4236 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4237 VDD D3 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4238 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4239 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4240 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4241 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4242 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4243 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4244 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4245 VDD D2 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4246 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4247 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4248 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4249 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4250 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4251 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4252 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4253 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4254 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4255 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4256 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4257 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4258 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4259 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4260 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4261 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4262 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4263 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4264 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4265 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4266 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4267 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4268 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4269 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4270 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4271 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R528 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R529 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R530 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R531 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4272 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4273 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4274 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4275 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4276 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4277 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4278 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4279 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4280 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4281 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4282 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4283 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4284 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4285 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4286 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4287 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4288 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4289 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4290 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4291 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4292 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4293 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4294 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4295 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R532 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R533 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R534 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R535 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4296 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4297 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4298 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4299 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4300 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4301 VDD D2 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4302 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4303 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4304 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4305 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4306 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4307 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4308 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4309 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4310 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4311 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4312 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4313 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4314 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4315 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4316 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4317 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4318 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4319 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4320 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4321 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4322 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4323 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4324 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4325 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4326 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4327 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R536 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R537 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R538 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R539 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4328 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4329 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4330 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4331 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4332 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4333 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4334 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4335 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4336 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4337 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4338 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4339 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4340 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4341 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4342 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4343 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4344 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4345 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4346 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4347 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4348 VDD 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4349 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4350 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4351 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R540 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R541 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R542 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R543 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4352 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4353 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4354 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4355 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4356 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4357 VDD D4 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4358 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X4359 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4360 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4361 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4362 9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4363 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4364 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4365 VDD D3 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4366 9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X4367 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4368 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4369 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4370 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4371 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4372 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4373 VDD D2 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4374 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4375 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4376 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4377 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4378 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4379 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4380 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4381 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4382 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4383 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4384 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4385 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4386 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4387 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4388 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4389 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4390 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/m1_14_20144# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4391 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4392 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4393 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4394 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4395 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4396 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4397 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4398 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4399 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R544 9good_1/8good_0/7good_0/6good_0/m1_14_20144# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R545 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R546 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R547 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4400 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4401 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4402 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4403 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4404 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4405 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4406 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4407 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4408 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4409 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4410 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4411 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4412 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4413 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4414 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4415 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4416 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4417 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4418 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4419 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4420 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4421 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4422 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4423 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R548 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R549 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R550 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R551 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4424 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4425 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4426 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4427 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4428 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4429 VDD D2 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4430 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4431 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4432 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4433 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4434 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4435 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4436 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4437 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4438 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4439 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4440 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4441 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4442 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4443 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4444 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4445 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4446 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4447 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4448 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4449 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4450 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4451 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4452 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4453 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4454 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4455 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R552 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R553 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R554 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R555 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4456 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4457 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4458 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4459 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4460 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4461 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4462 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4463 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4464 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4465 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4466 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4467 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4468 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4469 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4470 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4471 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4472 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4473 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4474 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4475 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4476 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4477 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4478 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4479 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R556 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R557 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R558 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R559 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4480 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4481 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4482 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4483 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4484 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4485 VDD D3 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4486 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4487 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4488 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4489 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4490 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4491 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4492 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4493 VDD D2 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4494 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4495 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4496 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4497 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4498 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4499 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4500 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4501 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4502 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4503 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4504 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4505 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4506 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4507 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4508 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4509 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4510 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4511 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4512 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4513 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4514 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4515 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4516 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4517 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4518 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4519 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R560 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R561 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R562 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R563 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4520 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4521 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4522 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4523 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4524 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4525 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4526 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4527 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4528 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4529 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4530 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4531 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4532 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4533 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4534 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4535 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4536 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4537 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4538 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4539 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4540 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4541 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4542 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4543 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R564 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R565 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R566 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R567 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4544 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4545 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4546 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4547 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4548 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4549 VDD D2 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4550 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4551 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4552 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4553 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4554 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4555 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4556 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4557 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4558 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4559 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4560 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4561 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4562 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4563 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4564 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4565 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4566 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4567 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4568 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4569 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4570 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4571 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4572 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4573 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4574 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4575 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R568 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R569 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R570 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R571 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4576 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4577 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4578 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4579 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4580 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4581 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4582 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4583 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4584 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4585 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4586 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4587 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4588 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4589 VDD D0 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4590 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4591 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4592 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4593 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4594 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4595 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4596 VDD 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4597 VDD D1 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4598 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4599 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R572 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R573 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R574 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_36912_2# sky130_fd_pr__res_generic_po1 w=66 l=342
R575 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4600 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4601 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/m1_8436_40544# 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X4602 9good_1/8good_0/7good_0/m1_8436_40544# 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4603 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4604 VDD 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4605 VDD D5 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4606 9good_1/8good_0/7good_0/m1_8436_40544# 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 9good_1/8good_0/7good_0/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X4607 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4608 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4609 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4610 9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4611 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4612 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4613 VDD D4 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4614 9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X4615 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4616 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4617 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4618 9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4619 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4620 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4621 VDD D3 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4622 9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X4623 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4624 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4625 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4626 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4627 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4628 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4629 VDD D2 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4630 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4631 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4632 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4633 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4634 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4635 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4636 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4637 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4638 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4639 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4640 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4641 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4642 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_46616_8# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4643 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4644 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4645 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4646 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_46616_8# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4647 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4648 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4649 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4650 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4651 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4652 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4653 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4654 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4655 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R576 m1_46616_8# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R577 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R578 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R579 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4656 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4657 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4658 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4659 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4660 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4661 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4662 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4663 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4664 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4665 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4666 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4667 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4668 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4669 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4670 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4671 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4672 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4673 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4674 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4675 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4676 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4677 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4678 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4679 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R580 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R581 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R582 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R583 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4680 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4681 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4682 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4683 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4684 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4685 VDD D2 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4686 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4687 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4688 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4689 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4690 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4691 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4692 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4693 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4694 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4695 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4696 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4697 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4698 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4699 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4700 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4701 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4702 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4703 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4704 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4705 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4706 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4707 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4708 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4709 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4710 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4711 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R584 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R585 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R586 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R587 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4712 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4713 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4714 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4715 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4716 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4717 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4718 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4719 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4720 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4721 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4722 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4723 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4724 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4725 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4726 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4727 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4728 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4729 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4730 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4731 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4732 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4733 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4734 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4735 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R588 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R589 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R590 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R591 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4736 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4737 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4738 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4739 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4740 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4741 VDD D3 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4742 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4743 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4744 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4745 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4746 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4747 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4748 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4749 VDD D2 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4750 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4751 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4752 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4753 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4754 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4755 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4756 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4757 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4758 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4759 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4760 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4761 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4762 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4763 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4764 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4765 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4766 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4767 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4768 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4769 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4770 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4771 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4772 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4773 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4774 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4775 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R592 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R593 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R594 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R595 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4776 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4777 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4778 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4779 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4780 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4781 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4782 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4783 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4784 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4785 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4786 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4787 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4788 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4789 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4790 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4791 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4792 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4793 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4794 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4795 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4796 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4797 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4798 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4799 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R596 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R597 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R598 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R599 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4800 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4801 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4802 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4803 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4804 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4805 VDD D2 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4806 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4807 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4808 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4809 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4810 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4811 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4812 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4813 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4814 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4815 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4816 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4817 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4818 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4819 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4820 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4821 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4822 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4823 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4824 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4825 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4826 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4827 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4828 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4829 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4830 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4831 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R600 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R601 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R602 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R603 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4832 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4833 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4834 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4835 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4836 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4837 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4838 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4839 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4840 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4841 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4842 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4843 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4844 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4845 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4846 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4847 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4848 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4849 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4850 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4851 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4852 VDD 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4853 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4854 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4855 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R604 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R605 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R606 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R607 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4856 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4857 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4858 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4859 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4860 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4861 VDD D4 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4862 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X4863 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4864 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4865 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4866 9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4867 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4868 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4869 VDD D3 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4870 9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X4871 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4872 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4873 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4874 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4875 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4876 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4877 VDD D2 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4878 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4879 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4880 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4881 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4882 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4883 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4884 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4885 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4886 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4887 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4888 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4889 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4890 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4891 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4892 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4893 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4894 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/m1_14_20144# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4895 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4896 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4897 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4898 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4899 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4900 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4901 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4902 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4903 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R608 9good_1/8good_0/7good_0/6good_1/m1_14_20144# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R609 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R610 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R611 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4904 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4905 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4906 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4907 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4908 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4909 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4910 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4911 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4912 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4913 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4914 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4915 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4916 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4917 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4918 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4919 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4920 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4921 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4922 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4923 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4924 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4925 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4926 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4927 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R612 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R613 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R614 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R615 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4928 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4929 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4930 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4931 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4932 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4933 VDD D2 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4934 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4935 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4936 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4937 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4938 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4939 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4940 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4941 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4942 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4943 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4944 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4945 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4946 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4947 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4948 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4949 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4950 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4951 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4952 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4953 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4954 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4955 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4956 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4957 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4958 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4959 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R616 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R617 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R618 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R619 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4960 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4961 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4962 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4963 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4964 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4965 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4966 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4967 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4968 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4969 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4970 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4971 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4972 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4973 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4974 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4975 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4976 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4977 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4978 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4979 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4980 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4981 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4982 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4983 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R620 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R621 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R622 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R623 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X4984 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4985 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4986 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4987 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4988 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4989 VDD D3 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4990 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4991 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4992 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4993 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4994 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4995 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X4996 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4997 VDD D2 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X4998 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4999 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5000 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5001 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5002 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5003 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5004 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5005 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5006 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5007 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5008 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5009 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5010 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5011 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5012 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5013 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5014 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5015 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5016 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5017 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5018 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5019 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5020 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5021 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5022 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5023 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R624 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R625 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R626 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R627 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5024 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5025 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5026 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5027 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5028 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5029 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5030 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5031 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5032 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5033 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5034 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5035 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5036 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5037 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5038 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5039 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5040 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5041 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5042 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5043 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5044 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5045 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5046 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5047 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R628 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R629 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R630 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R631 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5048 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5049 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5050 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5051 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5052 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5053 VDD D2 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5054 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5055 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5056 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5057 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5058 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5059 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5060 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5061 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5062 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5063 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5064 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5065 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5066 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5067 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5068 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5069 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5070 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5071 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5072 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5073 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5074 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5075 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5076 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5077 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5078 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5079 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R632 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R633 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R634 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R635 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5080 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5081 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5082 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5083 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5084 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5085 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5086 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5087 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5088 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5089 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5090 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5091 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5092 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5093 VDD D0 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5094 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5095 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5096 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5097 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5098 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5099 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5100 VDD 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5101 VDD D1 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5102 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5103 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R636 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R637 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R638 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_41532_78# sky130_fd_pr__res_generic_po1 w=66 l=342
R639 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5104 9good_1/8good_0/Sw-1_0/li_29_719# D7 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5105 9good_1/8good_0/m1_8774_43264# 9good_1/8good_0/Sw-1_0/li_29_719# 9good_1/m1_19068_42976# 9good_1/8good_0/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X5106 9good_1/m1_19068_42976# 9good_1/8good_0/Sw-1_0/li_29_719# 9good_1/8good_0/m1_18694_42308# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5107 9good_1/8good_0/Sw-1_0/li_126_470# 9good_1/8good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5108 VDD 9good_1/8good_0/Sw-1_0/li_29_719# 9good_1/8good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5109 VDD D7 9good_1/8good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5110 9good_1/m1_19068_42976# 9good_1/8good_0/Sw-1_0/li_126_470# 9good_1/8good_0/m1_18694_42308# 9good_1/m1_19068_42976# sky130_fd_pr__pfet_01v8 w=84 l=30
X5111 9good_1/8good_0/m1_8774_43264# 9good_1/8good_0/Sw-1_0/li_126_470# 9good_1/m1_19068_42976# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5112 9good_1/8good_0/7good_1/Sw-1_0/li_29_719# D6 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5113 9good_1/8good_0/7good_1/m1_4396_20620# 9good_1/8good_0/7good_1/Sw-1_0/li_29_719# 9good_1/8good_0/m1_18694_42308# 9good_1/8good_0/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X5114 9good_1/8good_0/m1_18694_42308# 9good_1/8good_0/7good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5115 9good_1/8good_0/7good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5116 VDD 9good_1/8good_0/7good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5117 VDD D6 9good_1/8good_0/7good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5118 9good_1/8good_0/m1_18694_42308# 9good_1/8good_0/7good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/m1_8436_40544# 9good_1/8good_0/m1_18694_42308# sky130_fd_pr__pfet_01v8 w=84 l=30
X5119 9good_1/8good_0/7good_1/m1_4396_20620# 9good_1/8good_0/7good_1/Sw-1_0/li_126_470# 9good_1/8good_0/m1_18694_42308# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5120 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5121 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/m1_4396_20620# 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X5122 9good_1/8good_0/7good_1/m1_4396_20620# 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5123 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5124 VDD 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5125 VDD D5 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5126 9good_1/8good_0/7good_1/m1_4396_20620# 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 9good_1/8good_0/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X5127 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/m1_4396_20620# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5128 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5129 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5130 9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5131 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5132 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5133 VDD D4 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5134 9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 9good_1/8good_0/7good_1/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X5135 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5136 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5137 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5138 9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5139 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5140 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5141 VDD D3 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5142 9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X5143 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5144 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5145 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5146 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5147 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5148 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5149 VDD D2 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5150 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5151 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5152 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5153 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5154 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5155 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5156 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5157 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5158 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5159 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5160 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5161 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5162 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_51780_62# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5163 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5164 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5165 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5166 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_51780_62# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5167 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5168 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5169 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5170 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5171 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5172 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5173 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5174 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5175 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R640 m1_51780_62# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R641 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R642 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R643 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5176 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5177 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5178 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5179 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5180 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5181 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5182 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5183 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5184 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5185 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5186 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5187 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5188 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5189 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5190 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5191 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5192 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5193 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5194 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5195 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5196 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5197 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5198 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5199 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R644 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R645 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R646 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R647 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5200 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5201 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5202 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5203 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5204 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5205 VDD D2 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5206 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5207 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5208 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5209 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5210 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5211 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5212 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5213 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5214 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5215 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5216 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5217 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5218 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5219 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5220 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5221 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5222 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5223 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5224 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5225 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5226 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5227 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5228 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5229 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5230 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5231 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R648 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R649 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R650 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R651 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5232 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5233 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5234 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5235 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5236 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5237 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5238 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5239 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5240 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5241 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5242 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5243 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5244 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5245 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5246 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5247 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5248 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5249 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5250 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5251 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5252 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5253 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5254 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5255 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R652 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R653 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R654 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R655 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5256 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5257 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5258 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5259 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5260 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5261 VDD D3 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5262 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5263 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5264 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5265 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5266 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5267 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5268 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5269 VDD D2 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5270 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5271 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5272 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5273 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5274 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5275 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5276 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5277 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5278 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5279 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5280 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5281 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5282 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5283 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5284 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5285 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5286 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5287 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5288 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5289 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5290 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5291 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5292 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5293 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5294 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5295 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R656 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R657 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R658 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R659 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5296 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5297 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5298 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5299 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5300 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5301 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5302 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5303 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5304 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5305 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5306 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5307 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5308 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5309 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5310 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5311 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5312 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5313 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5314 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5315 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5316 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5317 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5318 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5319 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R660 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R661 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R662 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R663 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5320 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5321 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5322 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5323 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5324 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5325 VDD D2 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5326 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5327 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5328 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5329 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5330 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5331 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5332 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5333 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5334 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5335 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5336 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5337 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5338 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5339 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5340 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5341 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5342 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5343 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5344 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5345 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5346 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5347 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5348 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5349 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5350 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5351 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R664 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R665 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R666 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R667 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5352 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5353 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5354 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5355 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5356 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5357 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5358 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5359 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5360 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5361 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5362 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5363 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5364 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5365 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5366 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5367 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5368 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5369 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5370 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5371 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5372 VDD 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5373 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5374 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5375 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R668 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R669 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R670 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R671 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5376 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5377 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5378 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5379 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5380 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5381 VDD D4 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5382 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X5383 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5384 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5385 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5386 9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5387 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5388 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5389 VDD D3 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5390 9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X5391 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5392 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5393 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5394 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5395 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5396 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5397 VDD D2 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5398 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5399 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5400 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5401 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5402 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5403 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5404 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5405 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5406 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5407 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5408 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5409 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5410 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5411 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5412 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5413 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5414 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/m1_14_20144# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5415 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5416 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5417 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5418 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5419 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5420 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5421 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5422 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5423 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R672 9good_1/8good_0/7good_1/6good_0/m1_14_20144# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R673 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R674 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R675 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5424 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5425 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5426 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5427 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5428 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5429 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5430 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5431 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5432 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5433 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5434 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5435 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5436 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5437 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5438 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5439 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5440 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5441 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5442 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5443 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5444 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5445 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5446 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5447 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R676 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R677 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R678 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R679 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5448 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5449 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5450 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5451 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5452 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5453 VDD D2 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5454 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5455 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5456 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5457 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5458 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5459 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5460 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5461 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5462 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5463 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5464 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5465 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5466 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5467 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5468 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5469 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5470 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5471 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5472 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5473 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5474 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5475 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5476 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5477 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5478 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5479 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R680 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R681 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R682 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R683 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5480 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5481 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5482 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5483 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5484 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5485 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5486 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5487 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5488 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5489 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5490 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5491 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5492 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5493 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5494 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5495 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5496 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5497 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5498 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5499 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5500 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5501 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5502 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5503 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R684 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R685 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R686 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R687 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5504 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5505 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5506 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5507 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5508 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5509 VDD D3 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5510 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5511 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5512 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5513 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5514 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5515 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5516 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5517 VDD D2 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5518 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5519 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5520 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5521 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5522 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5523 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5524 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5525 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5526 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5527 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5528 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5529 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5530 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5531 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5532 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5533 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5534 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5535 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5536 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5537 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5538 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5539 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5540 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5541 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5542 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5543 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R688 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R689 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R690 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R691 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5544 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5545 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5546 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5547 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5548 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5549 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5550 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5551 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5552 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5553 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5554 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5555 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5556 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5557 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5558 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5559 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5560 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5561 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5562 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5563 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5564 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5565 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5566 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5567 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R692 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R693 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R694 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R695 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5568 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5569 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5570 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5571 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5572 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5573 VDD D2 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5574 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5575 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5576 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5577 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5578 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5579 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5580 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5581 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5582 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5583 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5584 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5585 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5586 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5587 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5588 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5589 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5590 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5591 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5592 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5593 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5594 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5595 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5596 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5597 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5598 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5599 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R696 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R697 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R698 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R699 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5600 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5601 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5602 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5603 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5604 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5605 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5606 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5607 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5608 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5609 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5610 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5611 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5612 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5613 VDD D0 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5614 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5615 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5616 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5617 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5618 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5619 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5620 VDD 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5621 VDD D1 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5622 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5623 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R700 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R701 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R702 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_46616_8# sky130_fd_pr__res_generic_po1 w=66 l=342
R703 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5624 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5625 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/m1_8436_40544# 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X5626 9good_1/8good_0/7good_1/m1_8436_40544# 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5627 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5628 VDD 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5629 VDD D5 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5630 9good_1/8good_0/7good_1/m1_8436_40544# 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 9good_1/8good_0/7good_1/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X5631 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5632 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5633 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5634 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5635 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5636 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5637 VDD D4 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5638 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X5639 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5640 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5641 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5642 9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5643 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5644 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5645 VDD D3 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5646 9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X5647 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5648 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5649 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5650 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5651 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5652 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5653 VDD D2 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5654 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5655 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5656 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5657 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5658 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5659 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5660 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5661 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5662 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5663 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5664 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5665 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5666 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_56844_12# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5667 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5668 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5669 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5670 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_56844_12# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5671 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5672 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5673 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5674 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5675 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5676 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5677 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5678 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5679 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R704 m1_56844_12# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R705 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R706 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R707 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5680 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5681 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5682 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5683 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5684 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5685 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5686 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5687 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5688 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5689 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5690 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5691 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5692 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5693 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5694 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5695 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5696 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5697 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5698 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5699 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5700 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5701 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5702 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5703 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R708 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R709 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R710 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R711 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5704 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5705 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5706 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5707 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5708 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5709 VDD D2 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5710 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5711 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5712 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5713 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5714 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5715 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5716 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5717 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5718 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5719 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5720 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5721 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5722 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5723 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5724 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5725 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5726 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5727 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5728 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5729 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5730 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5731 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5732 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5733 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5734 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5735 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R712 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R713 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R714 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R715 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5736 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5737 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5738 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5739 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5740 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5741 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5742 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5743 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5744 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5745 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5746 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5747 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5748 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5749 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5750 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5751 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5752 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5753 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5754 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5755 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5756 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5757 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5758 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5759 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R716 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R717 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R718 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R719 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5760 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5761 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5762 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5763 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5764 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5765 VDD D3 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5766 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5767 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5768 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5769 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5770 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5771 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5772 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5773 VDD D2 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5774 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5775 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5776 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5777 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5778 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5779 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5780 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5781 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5782 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5783 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5784 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5785 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5786 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5787 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5788 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5789 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5790 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5791 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5792 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5793 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5794 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5795 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5796 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5797 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5798 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5799 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R720 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R721 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R722 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R723 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5800 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5801 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5802 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5803 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5804 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5805 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5806 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5807 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5808 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5809 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5810 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5811 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5812 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5813 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5814 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5815 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5816 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5817 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5818 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5819 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5820 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5821 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5822 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5823 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R724 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R725 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R726 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R727 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5824 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5825 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5826 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5827 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5828 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5829 VDD D2 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5830 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5831 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5832 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5833 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5834 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5835 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5836 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5837 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5838 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5839 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5840 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5841 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5842 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5843 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5844 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5845 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5846 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5847 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5848 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5849 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5850 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5851 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5852 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5853 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5854 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5855 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R728 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R729 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R730 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R731 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5856 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5857 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5858 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5859 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5860 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5861 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5862 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5863 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5864 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5865 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5866 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5867 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5868 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5869 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5870 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5871 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5872 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5873 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5874 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5875 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5876 VDD 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5877 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5878 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5879 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R732 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R733 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R734 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R735 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5880 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5881 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5882 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5883 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5884 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5885 VDD D4 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5886 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X5887 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5888 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5889 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5890 9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5891 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5892 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5893 VDD D3 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5894 9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X5895 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5896 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5897 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5898 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5899 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5900 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5901 VDD D2 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5902 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5903 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5904 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5905 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5906 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5907 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5908 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5909 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5910 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5911 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5912 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5913 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5914 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5915 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5916 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5917 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5918 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/m1_14_20144# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5919 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5920 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5921 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5922 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5923 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5924 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5925 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5926 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5927 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R736 9good_1/8good_0/7good_1/6good_1/m1_14_20144# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R737 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R738 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R739 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5928 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5929 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5930 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5931 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5932 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5933 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5934 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5935 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5936 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5937 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5938 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5939 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5940 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5941 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5942 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5943 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5944 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5945 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5946 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5947 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5948 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5949 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5950 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5951 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R740 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R741 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R742 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R743 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5952 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5953 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5954 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5955 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5956 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5957 VDD D2 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5958 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5959 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5960 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5961 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5962 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5963 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5964 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5965 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5966 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5967 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5968 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5969 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5970 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5971 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5972 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5973 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5974 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5975 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5976 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5977 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5978 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5979 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5980 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5981 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5982 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5983 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R744 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R745 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R746 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R747 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X5984 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5985 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5986 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5987 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5988 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5989 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5990 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5991 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5992 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5993 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5994 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5995 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X5996 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5997 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X5998 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5999 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6000 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6001 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6002 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6003 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6004 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6005 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6006 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6007 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R748 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R749 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R750 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R751 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6008 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6009 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6010 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6011 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6012 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6013 VDD D3 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6014 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6015 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6016 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6017 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6018 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6019 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6020 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6021 VDD D2 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6022 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6023 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6024 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6025 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6026 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6027 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6028 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6029 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6030 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6031 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6032 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6033 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6034 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6035 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6036 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6037 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6038 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6039 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6040 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6041 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6042 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6043 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6044 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6045 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6046 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6047 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R752 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R753 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R754 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R755 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6048 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6049 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6050 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6051 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6052 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6053 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6054 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6055 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6056 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6057 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6058 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6059 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6060 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6061 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6062 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6063 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6064 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6065 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6066 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6067 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6068 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6069 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6070 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6071 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R756 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R757 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R758 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R759 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6072 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6073 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6074 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6075 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6076 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6077 VDD D2 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6078 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6079 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6080 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6081 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6082 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6083 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6084 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6085 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6086 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6087 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6088 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6089 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6090 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6091 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6092 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6093 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6094 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6095 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6096 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6097 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6098 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6099 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6100 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6101 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6102 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6103 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R760 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R761 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R762 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R763 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6104 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6105 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6106 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6107 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6108 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6109 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6110 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6111 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6112 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# D0 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6113 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6114 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6115 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6116 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6117 VDD D0 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6118 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6119 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6120 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# D1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6121 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6122 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6123 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6124 VDD 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6125 VDD D1 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6126 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6127 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R764 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R765 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R766 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_51780_62# sky130_fd_pr__res_generic_po1 w=66 l=342
R767 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6128 9good_1/8good_1/7good_0/Sw-1_0/li_29_719# D6 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6129 9good_1/8good_1/7good_0/m1_4396_20620# 9good_1/8good_1/7good_0/Sw-1_0/li_29_719# 9good_1/8good_1/m1_8774_43264# 9good_1/8good_1/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X6130 9good_1/8good_1/m1_8774_43264# 9good_1/8good_1/7good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6131 9good_1/8good_1/7good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6132 VDD 9good_1/8good_1/7good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6133 VDD D6 9good_1/8good_1/7good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6134 9good_1/8good_1/m1_8774_43264# 9good_1/8good_1/7good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/m1_8436_40544# 9good_1/8good_1/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X6135 9good_1/8good_1/7good_0/m1_4396_20620# 9good_1/8good_1/7good_0/Sw-1_0/li_126_470# 9good_1/8good_1/m1_8774_43264# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6136 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6137 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/m1_4396_20620# 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X6138 9good_1/8good_1/7good_0/m1_4396_20620# 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6139 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6140 VDD 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6141 VDD D5 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6142 9good_1/8good_1/7good_0/m1_4396_20620# 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 9good_1/8good_1/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X6143 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/m1_4396_20620# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6144 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6145 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6146 9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6147 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6148 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6149 VDD D4 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6150 9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 9good_1/8good_1/7good_0/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X6151 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6152 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6153 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6154 9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6155 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6156 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6157 VDD D3 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6158 9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X6159 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6160 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6161 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6162 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6163 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6164 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6165 VDD D2 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6166 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6167 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6168 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6169 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6170 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6171 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6172 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6173 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6174 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6175 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6176 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6177 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6178 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_61528_92# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6179 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6180 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6181 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6182 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_61528_92# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6183 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6184 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6185 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6186 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6187 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6188 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6189 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6190 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6191 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R768 m1_61528_92# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R769 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R770 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R771 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6192 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6193 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6194 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6195 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6196 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6197 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6198 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6199 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6200 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6201 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6202 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6203 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6204 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6205 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6206 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6207 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6208 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6209 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6210 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6211 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6212 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6213 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6214 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6215 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R772 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R773 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R774 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R775 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6216 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6217 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6218 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6219 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6220 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6221 VDD D2 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6222 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6223 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6224 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6225 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6226 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6227 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6228 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6229 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6230 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6231 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6232 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6233 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6234 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6235 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6236 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6237 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6238 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6239 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6240 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6241 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6242 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6243 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6244 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6245 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6246 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6247 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R776 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R777 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R778 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R779 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6248 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6249 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6250 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6251 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6252 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6253 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6254 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6255 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6256 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6257 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6258 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6259 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6260 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6261 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6262 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6263 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6264 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6265 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6266 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6267 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6268 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6269 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6270 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6271 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R780 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R781 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R782 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R783 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6272 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6273 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6274 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6275 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6276 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6277 VDD D3 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6278 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6279 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6280 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6281 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6282 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6283 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6284 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6285 VDD D2 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6286 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6287 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6288 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6289 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6290 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6291 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6292 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6293 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6294 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6295 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6296 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6297 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6298 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6299 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6300 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6301 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6302 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6303 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6304 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6305 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6306 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6307 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6308 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6309 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6310 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6311 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R784 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R785 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R786 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R787 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6312 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6313 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6314 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6315 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6316 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6317 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6318 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6319 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6320 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6321 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6322 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6323 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6324 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6325 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6326 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6327 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6328 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6329 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6330 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6331 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6332 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6333 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6334 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6335 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R788 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R789 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R790 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R791 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6336 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6337 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6338 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6339 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6340 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6341 VDD D2 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6342 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6343 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6344 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6345 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6346 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6347 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6348 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6349 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6350 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6351 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6352 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6353 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6354 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6355 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6356 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6357 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6358 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6359 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6360 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6361 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6362 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6363 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6364 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6365 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6366 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6367 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R792 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R793 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R794 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R795 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6368 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6369 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6370 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6371 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6372 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6373 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6374 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6375 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6376 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6377 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6378 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6379 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6380 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6381 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6382 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6383 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6384 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6385 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6386 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6387 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6388 VDD 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6389 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6390 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6391 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R796 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R797 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R798 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R799 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6392 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6393 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6394 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6395 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6396 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6397 VDD D4 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6398 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X6399 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6400 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6401 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6402 9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6403 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6404 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6405 VDD D3 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6406 9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X6407 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6408 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6409 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6410 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6411 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6412 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6413 VDD D2 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6414 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6415 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6416 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6417 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6418 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6419 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6420 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6421 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6422 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6423 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6424 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6425 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6426 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6427 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6428 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6429 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6430 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/m1_14_20144# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6431 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6432 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6433 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6434 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6435 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6436 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6437 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6438 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6439 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R800 9good_1/8good_1/7good_0/6good_0/m1_14_20144# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R801 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R802 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R803 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6440 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6441 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6442 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6443 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6444 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6445 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6446 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6447 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6448 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6449 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6450 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6451 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6452 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6453 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6454 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6455 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6456 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6457 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6458 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6459 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6460 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6461 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6462 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6463 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R804 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R805 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R806 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R807 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6464 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6465 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6466 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6467 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6468 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6469 VDD D2 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6470 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6471 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6472 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6473 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6474 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6475 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6476 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6477 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6478 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6479 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6480 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6481 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6482 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6483 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6484 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6485 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6486 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6487 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6488 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6489 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6490 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6491 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6492 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6493 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6494 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6495 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R808 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R809 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R810 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R811 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6496 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6497 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6498 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6499 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6500 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6501 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6502 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6503 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6504 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6505 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6506 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6507 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6508 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6509 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6510 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6511 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6512 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6513 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6514 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6515 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6516 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6517 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6518 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6519 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R812 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R813 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R814 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R815 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6520 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6521 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6522 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6523 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6524 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6525 VDD D3 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6526 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6527 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6528 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6529 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6530 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6531 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6532 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6533 VDD D2 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6534 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6535 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6536 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6537 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6538 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6539 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6540 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6541 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6542 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6543 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6544 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6545 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6546 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6547 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6548 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6549 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6550 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6551 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6552 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6553 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6554 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6555 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6556 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6557 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6558 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6559 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R816 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R817 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R818 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R819 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6560 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6561 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6562 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6563 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6564 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6565 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6566 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6567 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6568 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6569 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6570 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6571 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6572 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6573 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6574 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6575 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6576 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6577 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6578 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6579 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6580 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6581 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6582 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6583 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R820 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R821 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R822 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R823 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6584 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6585 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6586 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6587 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6588 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6589 VDD D2 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6590 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6591 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6592 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6593 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6594 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6595 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6596 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6597 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6598 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6599 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6600 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6601 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6602 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6603 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6604 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6605 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6606 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6607 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6608 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6609 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6610 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6611 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6612 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6613 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6614 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6615 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R824 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R825 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R826 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R827 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6616 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6617 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6618 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6619 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6620 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6621 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6622 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6623 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6624 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6625 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6626 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6627 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6628 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6629 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6630 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6631 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6632 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6633 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6634 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6635 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6636 VDD 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6637 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6638 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6639 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R828 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R829 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R830 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_56844_12# sky130_fd_pr__res_generic_po1 w=66 l=342
R831 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6640 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6641 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/m1_8436_40544# 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X6642 9good_1/8good_1/7good_0/m1_8436_40544# 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6643 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6644 VDD 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6645 VDD D5 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6646 9good_1/8good_1/7good_0/m1_8436_40544# 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 9good_1/8good_1/7good_0/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X6647 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6648 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6649 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6650 9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6651 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6652 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6653 VDD D4 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6654 9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 9good_1/8good_1/7good_0/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X6655 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6656 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6657 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6658 9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6659 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6660 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6661 VDD D3 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6662 9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X6663 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6664 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6665 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6666 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6667 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6668 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6669 VDD D2 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6670 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6671 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6672 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6673 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6674 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6675 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6676 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6677 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6678 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6679 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6680 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6681 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6682 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_66618_22# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6683 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6684 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6685 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6686 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_66618_22# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6687 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6688 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6689 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6690 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6691 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6692 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6693 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6694 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6695 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R832 m1_66618_22# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R833 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R834 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R835 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6696 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6697 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6698 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6699 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6700 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6701 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6702 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6703 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6704 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6705 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6706 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6707 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6708 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6709 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6710 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6711 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6712 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6713 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6714 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6715 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6716 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6717 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6718 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6719 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R836 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R837 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R838 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R839 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6720 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6721 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6722 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6723 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6724 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6725 VDD D2 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6726 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6727 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6728 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6729 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6730 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6731 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6732 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6733 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6734 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6735 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6736 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6737 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6738 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6739 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6740 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6741 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6742 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6743 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6744 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6745 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6746 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6747 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6748 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6749 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6750 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6751 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R840 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R841 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R842 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R843 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6752 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6753 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6754 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6755 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6756 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6757 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6758 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6759 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6760 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6761 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6762 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6763 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6764 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6765 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6766 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6767 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6768 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6769 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6770 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6771 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6772 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6773 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6774 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6775 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R844 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R845 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R846 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R847 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6776 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6777 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6778 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6779 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6780 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6781 VDD D3 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6782 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6783 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6784 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6785 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6786 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6787 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6788 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6789 VDD D2 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6790 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6791 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6792 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6793 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6794 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6795 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6796 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6797 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6798 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6799 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6800 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6801 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6802 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6803 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6804 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6805 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6806 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6807 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6808 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6809 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6810 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6811 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6812 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6813 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6814 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6815 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R848 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R849 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R850 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R851 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6816 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6817 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6818 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6819 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6820 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6821 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6822 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6823 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6824 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6825 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6826 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6827 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6828 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6829 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6830 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6831 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6832 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6833 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6834 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6835 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6836 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6837 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6838 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6839 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R852 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R853 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R854 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R855 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6840 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6841 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6842 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6843 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6844 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6845 VDD D2 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6846 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6847 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6848 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6849 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6850 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6851 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6852 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6853 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6854 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6855 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6856 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6857 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6858 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6859 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6860 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6861 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6862 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6863 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6864 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6865 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6866 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6867 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6868 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6869 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6870 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6871 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R856 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R857 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R858 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R859 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6872 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6873 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6874 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6875 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6876 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6877 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6878 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6879 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6880 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6881 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6882 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6883 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6884 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6885 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6886 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6887 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6888 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6889 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6890 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6891 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6892 VDD 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6893 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6894 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6895 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R860 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R861 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R862 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R863 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6896 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6897 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6898 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6899 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6900 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6901 VDD D4 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6902 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X6903 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6904 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6905 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6906 9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6907 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6908 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6909 VDD D3 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6910 9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X6911 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6912 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6913 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6914 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6915 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6916 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6917 VDD D2 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6918 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6919 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6920 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6921 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6922 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6923 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6924 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6925 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6926 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6927 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6928 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6929 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6930 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6931 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6932 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6933 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6934 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/m1_14_20144# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6935 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6936 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6937 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6938 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6939 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6940 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6941 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6942 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6943 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R864 9good_1/8good_1/7good_0/6good_1/m1_14_20144# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R865 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R866 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R867 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6944 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6945 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6946 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6947 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6948 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6949 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6950 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6951 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6952 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6953 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6954 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6955 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6956 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6957 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6958 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6959 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6960 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6961 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6962 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6963 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6964 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6965 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6966 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6967 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R868 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R869 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R870 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R871 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X6968 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6969 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6970 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6971 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6972 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6973 VDD D2 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6974 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6975 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6976 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6977 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6978 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6979 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6980 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6981 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6982 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6983 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6984 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6985 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6986 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6987 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6988 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6989 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6990 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6991 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6992 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6993 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6994 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6995 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X6996 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6997 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X6998 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6999 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R872 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R873 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R874 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R875 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7000 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7001 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7002 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7003 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7004 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7005 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7006 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7007 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7008 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7009 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7010 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7011 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7012 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7013 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7014 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7015 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7016 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7017 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7018 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7019 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7020 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7021 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7022 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7023 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R876 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R877 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R878 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R879 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7024 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7025 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7026 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7027 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7028 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7029 VDD D3 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7030 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7031 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7032 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7033 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7034 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7035 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7036 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7037 VDD D2 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7038 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7039 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7040 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7041 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7042 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7043 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7044 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7045 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7046 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7047 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7048 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7049 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7050 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7051 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7052 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7053 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7054 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7055 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7056 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7057 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7058 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7059 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7060 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7061 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7062 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7063 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R880 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R881 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R882 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R883 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7064 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7065 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7066 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7067 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7068 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7069 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7070 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7071 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7072 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7073 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7074 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7075 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7076 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7077 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7078 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7079 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7080 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7081 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7082 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7083 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7084 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7085 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7086 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7087 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R884 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R885 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R886 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R887 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7088 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7089 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7090 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7091 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7092 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7093 VDD D2 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7094 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7095 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7096 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7097 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7098 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7099 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7100 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7101 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7102 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7103 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7104 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7105 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7106 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7107 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7108 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7109 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7110 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7111 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7112 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7113 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7114 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7115 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7116 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7117 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7118 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7119 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R888 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R889 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R890 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R891 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7120 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7121 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7122 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7123 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7124 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7125 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7126 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7127 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7128 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7129 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7130 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7131 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7132 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7133 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7134 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7135 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7136 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7137 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7138 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7139 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7140 VDD 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7141 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7142 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7143 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R892 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R893 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R894 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_61528_92# sky130_fd_pr__res_generic_po1 w=66 l=342
R895 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7144 9good_1/8good_1/Sw-1_0/li_29_719# D7 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7145 9good_1/8good_1/m1_8774_43264# 9good_1/8good_1/Sw-1_0/li_29_719# 9good_1/m1_38716_44140# 9good_1/8good_1/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X7146 9good_1/m1_38716_44140# 9good_1/8good_1/Sw-1_0/li_29_719# 9good_1/8good_1/m1_18694_42308# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7147 9good_1/8good_1/Sw-1_0/li_126_470# 9good_1/8good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7148 VDD 9good_1/8good_1/Sw-1_0/li_29_719# 9good_1/8good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7149 VDD D7 9good_1/8good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7150 9good_1/m1_38716_44140# 9good_1/8good_1/Sw-1_0/li_126_470# 9good_1/8good_1/m1_18694_42308# 9good_1/m1_38716_44140# sky130_fd_pr__pfet_01v8 w=84 l=30
X7151 9good_1/8good_1/m1_8774_43264# 9good_1/8good_1/Sw-1_0/li_126_470# 9good_1/m1_38716_44140# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7152 9good_1/8good_1/7good_1/Sw-1_0/li_29_719# D6 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7153 9good_1/8good_1/7good_1/m1_4396_20620# 9good_1/8good_1/7good_1/Sw-1_0/li_29_719# 9good_1/8good_1/m1_18694_42308# 9good_1/8good_1/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X7154 9good_1/8good_1/m1_18694_42308# 9good_1/8good_1/7good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7155 9good_1/8good_1/7good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7156 VDD 9good_1/8good_1/7good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7157 VDD D6 9good_1/8good_1/7good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7158 9good_1/8good_1/m1_18694_42308# 9good_1/8good_1/7good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/m1_8436_40544# 9good_1/8good_1/m1_18694_42308# sky130_fd_pr__pfet_01v8 w=84 l=30
X7159 9good_1/8good_1/7good_1/m1_4396_20620# 9good_1/8good_1/7good_1/Sw-1_0/li_126_470# 9good_1/8good_1/m1_18694_42308# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7160 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7161 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/m1_4396_20620# 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X7162 9good_1/8good_1/7good_1/m1_4396_20620# 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7163 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7164 VDD 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7165 VDD D5 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7166 9good_1/8good_1/7good_1/m1_4396_20620# 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 9good_1/8good_1/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X7167 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/m1_4396_20620# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7168 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7169 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7170 9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7171 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7172 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7173 VDD D4 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7174 9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 9good_1/8good_1/7good_1/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X7175 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7176 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7177 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7178 9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7179 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7180 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7181 VDD D3 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7182 9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X7183 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7184 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7185 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7186 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7187 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7188 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7189 VDD D2 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7190 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7191 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7192 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7193 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7194 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7195 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7196 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7197 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7198 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7199 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7200 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7201 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7202 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_71736_52# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7203 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7204 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7205 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7206 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_71736_52# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7207 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7208 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7209 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7210 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7211 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7212 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7213 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7214 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7215 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R896 m1_71736_52# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R897 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R898 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R899 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7216 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7217 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7218 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7219 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7220 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7221 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7222 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7223 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7224 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7225 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7226 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7227 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7228 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7229 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7230 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7231 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7232 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7233 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7234 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7235 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7236 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7237 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7238 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7239 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R900 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R901 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R902 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R903 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7240 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7241 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7242 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7243 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7244 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7245 VDD D2 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7246 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7247 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7248 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7249 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7250 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7251 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7252 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7253 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7254 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7255 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7256 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7257 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7258 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7259 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7260 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7261 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7262 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7263 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7264 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7265 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7266 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7267 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7268 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7269 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7270 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7271 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R904 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R905 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R906 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R907 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7272 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7273 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7274 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7275 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7276 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7277 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7278 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7279 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7280 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7281 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7282 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7283 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7284 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7285 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7286 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7287 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7288 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7289 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7290 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7291 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7292 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7293 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7294 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7295 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R908 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R909 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R910 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R911 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7296 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7297 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7298 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7299 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7300 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7301 VDD D3 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7302 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7303 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7304 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7305 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7306 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7307 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7308 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7309 VDD D2 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7310 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7311 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7312 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7313 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7314 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7315 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7316 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7317 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7318 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7319 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7320 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7321 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7322 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7323 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7324 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7325 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7326 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7327 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7328 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7329 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7330 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7331 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7332 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7333 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7334 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7335 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R912 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R913 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R914 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R915 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7336 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7337 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7338 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7339 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7340 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7341 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7342 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7343 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7344 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7345 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7346 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7347 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7348 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7349 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7350 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7351 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7352 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7353 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7354 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7355 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7356 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7357 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7358 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7359 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R916 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R917 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R918 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R919 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7360 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7361 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7362 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7363 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7364 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7365 VDD D2 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7366 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7367 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7368 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7369 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7370 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7371 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7372 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7373 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7374 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7375 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7376 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7377 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7378 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7379 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7380 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7381 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7382 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7383 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7384 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7385 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7386 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7387 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7388 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7389 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7390 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7391 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R920 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R921 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R922 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R923 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7392 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7393 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7394 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7395 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7396 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7397 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7398 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7399 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7400 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7401 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7402 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7403 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7404 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7405 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7406 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7407 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7408 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7409 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7410 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7411 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7412 VDD 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7413 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7414 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7415 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R924 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R925 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R926 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R927 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7416 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7417 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7418 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7419 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7420 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7421 VDD D4 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7422 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X7423 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7424 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7425 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7426 9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7427 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7428 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7429 VDD D3 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7430 9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X7431 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7432 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7433 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7434 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7435 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7436 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7437 VDD D2 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7438 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7439 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7440 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7441 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7442 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7443 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7444 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7445 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7446 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7447 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7448 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7449 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7450 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7451 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7452 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7453 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7454 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/m1_14_20144# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7455 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7456 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7457 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7458 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7459 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7460 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7461 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7462 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7463 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R928 9good_1/8good_1/7good_1/6good_0/m1_14_20144# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R929 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R930 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R931 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7464 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7465 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7466 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7467 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7468 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7469 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7470 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7471 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7472 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7473 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7474 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7475 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7476 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7477 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7478 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7479 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7480 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7481 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7482 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7483 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7484 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7485 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7486 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7487 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R932 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R933 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R934 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R935 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7488 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7489 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7490 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7491 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7492 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7493 VDD D2 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7494 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7495 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7496 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7497 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7498 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7499 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7500 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7501 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7502 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7503 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7504 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7505 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7506 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7507 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7508 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7509 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7510 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7511 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7512 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7513 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7514 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7515 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7516 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7517 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7518 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7519 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R936 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R937 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R938 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R939 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7520 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7521 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7522 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7523 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7524 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7525 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7526 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7527 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7528 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7529 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7530 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7531 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7532 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7533 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7534 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7535 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7536 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7537 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7538 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7539 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7540 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7541 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7542 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7543 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R940 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R941 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R942 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R943 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7544 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7545 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7546 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7547 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7548 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7549 VDD D3 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7550 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7551 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7552 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7553 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7554 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7555 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7556 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7557 VDD D2 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7558 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7559 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7560 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7561 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7562 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7563 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7564 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7565 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7566 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7567 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7568 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7569 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7570 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7571 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7572 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7573 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7574 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7575 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7576 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7577 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7578 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7579 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7580 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7581 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7582 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7583 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R944 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R945 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R946 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R947 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7584 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7585 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7586 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7587 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7588 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7589 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7590 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7591 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7592 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7593 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7594 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7595 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7596 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7597 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7598 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7599 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7600 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7601 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7602 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7603 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7604 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7605 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7606 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7607 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R948 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R949 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R950 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R951 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7608 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7609 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7610 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7611 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7612 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7613 VDD D2 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7614 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7615 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7616 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7617 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7618 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7619 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7620 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7621 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7622 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7623 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7624 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7625 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7626 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7627 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7628 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7629 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7630 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7631 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7632 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7633 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7634 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7635 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7636 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7637 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7638 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7639 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R952 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R953 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R954 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R955 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7640 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7641 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7642 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7643 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7644 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7645 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7646 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7647 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7648 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7649 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7650 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7651 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7652 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7653 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7654 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7655 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7656 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7657 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7658 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7659 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7660 VDD 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7661 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7662 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7663 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R956 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R957 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R958 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_66618_22# sky130_fd_pr__res_generic_po1 w=66 l=342
R959 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7664 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# D5 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7665 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/m1_8436_40544# 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X7666 9good_1/8good_1/7good_1/m1_8436_40544# 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7667 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7668 VDD 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7669 VDD D5 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7670 9good_1/8good_1/7good_1/m1_8436_40544# 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 9good_1/8good_1/7good_1/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X7671 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/m1_8436_40544# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7672 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7673 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7674 9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7675 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7676 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7677 VDD D4 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7678 9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 9good_1/8good_1/7good_1/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X7679 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/m1_4002_19952# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7680 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7681 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7682 9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7683 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7684 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7685 VDD D3 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7686 9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X7687 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7688 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7689 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7690 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7691 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7692 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7693 VDD D2 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7694 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7695 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7696 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7697 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7698 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7699 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7700 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7701 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7702 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7703 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7704 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7705 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7706 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# m1_76798_18# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7707 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7708 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7709 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7710 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# m1_76798_18# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7711 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7712 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7713 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7714 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7715 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7716 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7717 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7718 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7719 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R960 m1_76798_18# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R961 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R962 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R963 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7720 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7721 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7722 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7723 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7724 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7725 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7726 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7727 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7728 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7729 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7730 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7731 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7732 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7733 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7734 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7735 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7736 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7737 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7738 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7739 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7740 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7741 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7742 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7743 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R964 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R965 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R966 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R967 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7744 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7745 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7746 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7747 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7748 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7749 VDD D2 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7750 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7751 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7752 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7753 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7754 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7755 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7756 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7757 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7758 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7759 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7760 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7761 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7762 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7763 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7764 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7765 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7766 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7767 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7768 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7769 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7770 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7771 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7772 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7773 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7774 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7775 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R968 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R969 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R970 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R971 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7776 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7777 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7778 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7779 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7780 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7781 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7782 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7783 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7784 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7785 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7786 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7787 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7788 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7789 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7790 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7791 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7792 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7793 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7794 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7795 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7796 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7797 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7798 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7799 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R972 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R973 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R974 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R975 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7800 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7801 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7802 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7803 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7804 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7805 VDD D3 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7806 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7807 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7808 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7809 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7810 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7811 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7812 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7813 VDD D2 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7814 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7815 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7816 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7817 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7818 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7819 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7820 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7821 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7822 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7823 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7824 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7825 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7826 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7827 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7828 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7829 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7830 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7831 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7832 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7833 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7834 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7835 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7836 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7837 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7838 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7839 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R976 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R977 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R978 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R979 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7840 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7841 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7842 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7843 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7844 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7845 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7846 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7847 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7848 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7849 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7850 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7851 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7852 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7853 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7854 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7855 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7856 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7857 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7858 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7859 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7860 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7861 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7862 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7863 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R980 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R981 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R982 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R983 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7864 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7865 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7866 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7867 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7868 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7869 VDD D2 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7870 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7871 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7872 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7873 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7874 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7875 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7876 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7877 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7878 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7879 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7880 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7881 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7882 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7883 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7884 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7885 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7886 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7887 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7888 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7889 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7890 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7891 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7892 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7893 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7894 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7895 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R984 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R985 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R986 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R987 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7896 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7897 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7898 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7899 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7900 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7901 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7902 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7903 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7904 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7905 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7906 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7907 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7908 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7909 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7910 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7911 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7912 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7913 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7914 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7915 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7916 VDD 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7917 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7918 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7919 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R988 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R989 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R990 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po1 w=66 l=342
R991 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7920 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# D4 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7921 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7922 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7923 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7924 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7925 VDD D4 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7926 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X7927 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7928 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7929 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7930 9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7931 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7932 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7933 VDD D3 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7934 9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X7935 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7936 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7937 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7938 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7939 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7940 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7941 VDD D2 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7942 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7943 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7944 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7945 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7946 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7947 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7948 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7949 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7950 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7951 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7952 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7953 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7954 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/m1_14_20144# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7955 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7956 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7957 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7958 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/m1_14_20144# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7959 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7960 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7961 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7962 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7963 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7964 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7965 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7966 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7967 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R992 9good_1/8good_1/7good_1/6good_1/m1_14_20144# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R993 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R994 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R995 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7968 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7969 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7970 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7971 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7972 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7973 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7974 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7975 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7976 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7977 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7978 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7979 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7980 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7981 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7982 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7983 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7984 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7985 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7986 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7987 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7988 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7989 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7990 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7991 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R996 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R997 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R998 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R999 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X7992 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7993 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7994 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7995 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X7996 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7997 VDD D2 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X7998 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7999 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8000 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8001 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8002 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8003 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8004 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8005 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8006 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8007 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8008 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8009 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8010 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8011 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8012 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8013 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8014 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8015 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8016 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8017 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8018 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8019 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8020 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8021 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8022 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X8023 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R1000 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R1001 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R1002 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R1003 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X8024 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8025 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8026 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8027 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8028 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8029 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8030 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8031 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8032 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8033 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8034 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8035 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8036 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8037 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8038 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8039 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8040 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8041 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8042 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8043 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8044 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8045 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8046 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8047 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R1004 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R1005 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R1006 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R1007 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X8048 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# D3 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8049 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X8050 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8051 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8052 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8053 VDD D3 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8054 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X8055 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8056 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8057 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8058 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8059 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8060 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8061 VDD D2 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8062 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X8063 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8064 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8065 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8066 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8067 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8068 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8069 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8070 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8071 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8072 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8073 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8074 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8075 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8076 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8077 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8078 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8079 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8080 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8081 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8082 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8083 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8084 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8085 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8086 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X8087 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R1008 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R1009 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R1010 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R1011 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X8088 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8089 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8090 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8091 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8092 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8093 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8094 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8095 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8096 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8097 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8098 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8099 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8100 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8101 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8102 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8103 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8104 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8105 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8106 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8107 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8108 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8109 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8110 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8111 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R1012 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R1013 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R1014 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R1015 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X8112 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# D2 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8113 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8114 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8115 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8116 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8117 VDD D2 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8118 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X8119 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8120 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8121 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8122 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8123 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8124 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8125 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8126 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8127 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8128 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8129 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8130 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8131 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8132 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8133 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8134 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8135 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8136 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8137 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8138 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8139 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8140 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8141 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8142 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X8143 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R1016 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R1017 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R1018 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# sky130_fd_pr__res_generic_po1 w=66 l=342
R1019 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X8144 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8145 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8146 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8147 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8148 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8149 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8150 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8151 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8152 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/m1_32342_44672# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8153 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8154 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8155 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8156 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8157 VDD 9good_1/m1_32342_44672# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8158 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8159 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8160 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/m1_32720_44664# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8161 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8162 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8163 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8164 VDD 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8165 VDD 9good_1/m1_32720_44664# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8166 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8167 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
R1020 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_1324# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po1 w=66 l=342
R1021 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po1 w=66 l=342
R1022 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# m1_71736_52# sky130_fd_pr__res_generic_po1 w=66 l=342
R1023 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po1 w=66 l=342
X8168 9good_1/Sw-1_0/li_29_719# D8 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8169 9good_1/m1_19068_42976# 9good_1/Sw-1_0/li_29_719# m1_78452_45530# 9good_1/m1_19068_42976# sky130_fd_pr__pfet_01v8 w=84 l=30
X8170 m1_78452_45530# 9good_1/Sw-1_0/li_29_719# 9good_1/m1_38716_44140# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8171 9good_1/Sw-1_0/li_126_470# 9good_1/Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8172 VDD 9good_1/Sw-1_0/li_29_719# 9good_1/Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8173 VDD D8 9good_1/Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8174 m1_78452_45530# 9good_1/Sw-1_0/li_126_470# 9good_1/m1_38716_44140# m1_78452_45530# sky130_fd_pr__pfet_01v8 w=84 l=30
X8175 9good_1/m1_19068_42976# 9good_1/Sw-1_0/li_126_470# m1_78452_45530# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8176 Sw-1_0/li_29_719# D9 VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8177 m1_39076_44800# Sw-1_0/li_29_719# Y m1_39076_44800# sky130_fd_pr__pfet_01v8 w=84 l=30
X8178 Y Sw-1_0/li_29_719# m1_78452_45530# VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8179 Sw-1_0/li_126_470# Sw-1_0/li_29_719# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
X8180 VDD Sw-1_0/li_29_719# Sw-1_0/li_126_470# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8181 VDD D9 Sw-1_0/li_29_719# VDD sky130_fd_pr__pfet_01v8 w=84 l=30
X8182 Y Sw-1_0/li_126_470# m1_78452_45530# Y sky130_fd_pr__pfet_01v8 w=84 l=30
X8183 m1_39076_44800# Sw-1_0/li_126_470# Y VSUBS sky130_fd_pr__nfet_01v8 w=84 l=30
C0 9good_0/8good_1/7good_1/m1_4396_20620# m1_31884_48# 2.94fF
C1 9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 3.90fF
C2 9good_1/8good_1/7good_0/m1_4396_20620# 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 3.52fF
C3 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C4 D3 9good_1/m1_32720_44664# 6.31fF
C5 GND D2 8.12fF
C6 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 2.60fF
C7 9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 2.83fF
C8 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 2.83fF
C9 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 3.90fF
C10 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 3.90fF
C11 9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 2.60fF
C12 9good_1/8good_0/7good_1/m1_8436_40544# 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 6.45fF
C13 D6 D3 2.20fF
C14 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C15 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 2.60fF
C16 9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 2.60fF
C17 9good_1/8good_1/7good_0/m1_4396_20620# m1_61528_92# 3.32fF
C18 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 2.83fF
C19 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 2.83fF
C20 D5 D0 15.72fF
C21 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 9good_0/8good_0/7good_1/m1_8436_40544# 6.45fF
C22 D3 9good_0/m1_32720_44664# 6.31fF
C23 D1 D0 84.52fF
C24 9good_1/m1_32720_44664# D2 36.73fF
C25 9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 3.90fF
C26 9good_1/8good_1/7good_0/m1_8436_40544# 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 6.45fF
C27 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 2.60fF
C28 9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 2.60fF
C29 9good_1/m1_32342_44672# D2 4.60fF
C30 9good_1/8good_1/7good_1/m1_8436_40544# 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 6.45fF
C31 D0 VDD 76.46fF
C32 9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 9good_1/8good_0/7good_0/m1_4396_20620# 3.52fF
C33 9good_0/8good_0/7good_1/m1_4396_20620# 9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 3.52fF
C34 9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 3.90fF
C35 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 3.90fF
C36 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 2.60fF
C37 9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C38 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 2.83fF
C39 D6 D8 7.17fF
C40 9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 3.90fF
C41 9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 2.60fF
C42 D5 D3 26.99fF
C43 D6 D7 45.83fF
C44 m1_36912_2# 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 4.81fF
C45 D3 D4 284.20fF
C46 m1_1684_72# D5 5.97fF
C47 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 2.60fF
C48 D1 D3 27.28fF
C49 9good_0/m1_32720_44664# D2 36.73fF
C50 9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 3.90fF
C51 9good_1/m1_32720_44664# GND 14.50fF
C52 D3 VDD 24.25fF
C53 9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 2.83fF
C54 9good_0/m1_32720_44664# 9good_0/m1_32342_44672# 17.70fF
C55 9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 2.83fF
C56 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 2.60fF
C57 9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 9good_0/8good_0/7good_0/m1_4396_20620# 3.52fF
C58 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 2.60fF
C59 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 9good_1/8good_0/7good_1/m1_4396_20620# 3.52fF
C60 m1_36912_2# 9good_0/8good_1/7good_1/m1_8436_40544# 16.29fF
C61 D5 D2 2.21fF
C62 D4 D2 48.21fF
C63 9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 2.83fF
C64 D1 D2 123.91fF
C65 D5 9good_0/m1_32342_44672# 7.88fF
C66 9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 2.83fF
C67 GND 9good_0/m1_32720_44664# 14.50fF
C68 D5 D7 14.81fF
C69 VDD D2 38.28fF
C70 9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 3.90fF
C71 9good_1/m1_32720_44664# 9good_1/m1_32342_44672# 17.70fF
C72 VDD 9good_0/m1_32342_44672# 38.23fF
C73 9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 2.83fF
C74 9good_1/8good_0/7good_1/m1_8436_40544# m1_56844_12# 22.51fF
C75 9good_0/8good_1/7good_0/m1_8436_40544# 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 6.45fF
C76 GND D4 8.37fF
C77 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 3.90fF
C78 9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 2.60fF
C79 D1 GND 29.00fF
C80 m1_51780_62# 9good_1/8good_0/7good_1/m1_4396_20620# 3.12fF
C81 m1_71736_52# 9good_1/8good_1/7good_1/m1_4396_20620# 3.17fF
C82 VDD GND 54.87fF
C83 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 2.60fF
C84 9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 2.60fF
C85 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 2.60fF
C86 9good_1/8good_1/7good_1/m1_8436_40544# m1_76798_18# 4.80fF
C87 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 2.83fF
C88 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 9good_1/8good_1/7good_1/m1_4396_20620# 3.52fF
C89 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 2.60fF
C90 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 2.83fF
C91 9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 2.60fF
C92 9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 3.90fF
C93 9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 3.90fF
C94 9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 9good_0/8good_1/7good_1/m1_8436_40544# 6.45fF
C95 D5 9good_1/m1_32342_44672# 7.88fF
C96 9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 2.60fF
C97 m1_56844_12# 9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 2.40fF
C98 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# m1_16966_2# 2.48fF
C99 9good_0/8good_1/7good_1/m1_4396_20620# 9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 3.52fF
C100 9good_1/m1_32720_44664# VDD 25.95fF
C101 9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C102 9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 9good_0/8good_0/7good_0/m1_8436_40544# 6.45fF
C103 D6 D5 70.67fF
C104 VDD 9good_1/m1_32342_44672# 38.23fF
C105 D0 D2 24.92fF
C106 D6 D4 18.95fF
C107 9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 2.60fF
C108 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 2.60fF
C109 9good_0/8good_0/7good_1/m1_4396_20620# m1_11882_62# 5.89fF
C110 m1_1684_72# 9good_0/8good_0/7good_0/m1_4396_20620# 6.48fF
C111 9good_0/8good_1/7good_0/m1_4396_20620# 9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 3.52fF
C112 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C113 9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 2.83fF
C114 VDD 9good_0/m1_32720_44664# 25.95fF
C115 9good_1/8good_0/7good_0/m1_4396_20620# m1_41532_78# 3.66fF
C116 9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 3.90fF
C117 D3 D2 301.30fF
C118 9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 2.83fF
C119 D5 m1_11882_62# 5.97fF
C120 9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 3.90fF
C121 9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C122 9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 2.83fF
C123 9good_1/m1_19068_42976# m1_39076_44800# 4.50fF
C124 D5 D4 86.18fF
C125 9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 2.60fF
C126 9good_0/8good_0/7good_1/m1_8436_40544# m1_16966_2# 26.51fF
C127 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 2.60fF
C128 D5 VDD 9.59fF
C129 9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 2.83fF
C130 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 2.60fF
C131 VDD D4 15.12fF
C132 9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 3.90fF
C133 9good_1/8good_0/7good_0/m1_8436_40544# 9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 6.45fF
C134 D1 VDD 51.90fF
C135 m1_6754_8# 9good_0/8good_0/7good_0/m1_8436_40544# 2.51fF
C136 9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 2.60fF
C137 9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C138 9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 3.90fF
C139 D3 GND 15.43fF
C140 9good_0/m1_32342_44672# D2 4.60fF
C141 m1_56844_12# 9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 2.55fF
C142 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 2.60fF
C143 D8 D7 23.76fF
C144 9good_0/8good_0/7good_1/6good_1/m1_4002_19952# m1_16966_2# 2.64fF
C145 9good_0/8good_1/7good_0/m1_4396_20620# m1_21660_68# 3.48fF
C146 Sw-1_0/li_29_719# VSUBS 2.05fF
C147 9good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C148 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C149 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C150 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C151 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C152 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C153 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C154 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C155 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C156 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C157 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C158 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C159 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C160 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C161 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C162 9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C163 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C164 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C165 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C166 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C167 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C168 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C169 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C170 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C171 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C172 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C173 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C174 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C175 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C176 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C177 9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C178 9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C179 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C180 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C181 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C182 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C183 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C184 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C185 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C186 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C187 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C188 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C189 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C190 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C191 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C192 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C193 9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C194 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C195 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C196 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C197 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C198 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C199 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C200 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C201 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C202 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C203 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C204 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C205 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C206 m1_76798_18# VSUBS 2.50fF
C207 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C208 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C209 9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C210 9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C211 9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C212 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C213 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C214 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C215 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C216 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C217 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C218 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C219 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C220 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C221 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C222 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C223 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C224 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C225 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C226 9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C227 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C228 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C229 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C230 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C231 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C232 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C233 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C234 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C235 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C236 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C237 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C238 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C239 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C240 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C241 9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C242 9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C243 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C244 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C245 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C246 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C247 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C248 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C249 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C250 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C251 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C252 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C253 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C254 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C255 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C256 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C257 9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C258 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C259 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C260 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C261 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C262 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C263 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C264 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C265 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C266 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C267 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C268 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C269 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C270 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C271 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C272 9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C273 9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C274 9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C275 9good_1/8good_1/7good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C276 9good_1/8good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C277 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C278 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C279 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C280 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C281 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C282 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C283 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C284 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C285 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C286 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C287 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C288 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C289 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C290 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C291 9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C292 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C293 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C294 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C295 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C296 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C297 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C298 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C299 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C300 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C301 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C302 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C303 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C304 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C305 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C306 9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C307 9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C308 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C309 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C310 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C311 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C312 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C313 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C314 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C315 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C316 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C317 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C318 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C319 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C320 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C321 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C322 9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C323 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C324 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C325 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C326 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C327 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C328 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C329 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C330 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C331 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C332 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C333 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C334 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C335 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C336 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C337 9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C338 9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C339 9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C340 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C341 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C342 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C343 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C344 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C345 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C346 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C347 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C348 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C349 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C350 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C351 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C352 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C353 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C354 9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C355 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C356 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C357 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C358 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C359 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C360 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C361 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C362 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C363 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C364 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C365 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C366 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C367 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C368 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C369 9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C370 9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C371 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C372 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C373 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C374 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C375 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C376 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C377 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C378 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C379 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C380 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C381 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C382 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C383 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C384 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C385 9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C386 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C387 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C388 9good_1/m1_32342_44672# VSUBS 178.26fF
C389 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C390 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C391 VDD VSUBS 1651.54fF
C392 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C393 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C394 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C395 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C396 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C397 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C398 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C399 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C400 m1_61528_92# VSUBS 2.71fF
C401 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C402 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C403 9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C404 9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C405 9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C406 9good_1/8good_1/7good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C407 9good_1/8good_1/m1_8774_43264# VSUBS 5.31fF
C408 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C409 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C410 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C411 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C412 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C413 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C414 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C415 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C416 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C417 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C418 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C419 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C420 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C421 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C422 9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C423 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C424 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C425 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C426 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C427 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C428 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C429 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C430 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C431 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C432 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C433 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C434 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C435 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C436 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C437 9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C438 9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C439 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C440 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C441 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C442 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C443 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C444 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C445 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C446 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C447 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C448 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C449 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C450 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C451 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C452 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C453 9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C454 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C455 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C456 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C457 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C458 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C459 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C460 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C461 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C462 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C463 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C464 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C465 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C466 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C467 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C468 9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C469 9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C470 9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C471 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C472 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C473 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C474 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C475 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C476 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C477 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C478 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C479 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C480 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C481 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C482 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C483 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C484 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C485 9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C486 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C487 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C488 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C489 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C490 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C491 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C492 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C493 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C494 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C495 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C496 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C497 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C498 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C499 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C500 9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C501 9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C502 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C503 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C504 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C505 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C506 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C507 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C508 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C509 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C510 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C511 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C512 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C513 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C514 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C515 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C516 9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C517 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C518 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C519 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C520 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C521 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C522 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C523 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C524 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C525 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C526 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C527 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C528 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C529 m1_51780_62# VSUBS 2.67fF
C530 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C531 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C532 9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C533 9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C534 9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C535 9good_1/8good_0/7good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C536 9good_1/8good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C537 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C538 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C539 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C540 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C541 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C542 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C543 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C544 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C545 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C546 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C547 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C548 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C549 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C550 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C551 9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C552 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C553 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C554 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C555 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C556 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C557 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C558 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C559 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C560 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C561 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C562 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C563 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C564 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C565 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C566 9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C567 9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C568 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C569 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C570 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C571 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C572 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C573 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C574 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C575 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C576 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C577 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C578 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C579 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C580 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C581 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C582 9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C583 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C584 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C585 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C586 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C587 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C588 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C589 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C590 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C591 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C592 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C593 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C594 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C595 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C596 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C597 9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C598 9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C599 9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C600 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C601 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C602 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C603 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C604 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C605 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C606 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C607 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C608 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C609 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C610 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C611 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C612 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C613 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C614 9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C615 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C616 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C617 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C618 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C619 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C620 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C621 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C622 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C623 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C624 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C625 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C626 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C627 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C628 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C629 9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C630 9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C631 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C632 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C633 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C634 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C635 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C636 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C637 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C638 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C639 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C640 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C641 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C642 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C643 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C644 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C645 9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C646 GND VSUBS 451.33fF **FLOATING
C647 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C648 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C649 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C650 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C651 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C652 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C653 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C654 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C655 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C656 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C657 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C658 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C659 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C660 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C661 9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C662 9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C663 9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C664 9good_1/8good_0/7good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C665 9good_1/8good_0/m1_8774_43264# VSUBS 5.31fF
C666 9good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C667 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C668 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C669 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C670 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C671 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C672 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C673 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C674 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C675 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C676 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C677 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C678 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C679 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C680 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C681 9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C682 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C683 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C684 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C685 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C686 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C687 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C688 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C689 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C690 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C691 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C692 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C693 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C694 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C695 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C696 9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C697 9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C698 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C699 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C700 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C701 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C702 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C703 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C704 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C705 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C706 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C707 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C708 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C709 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C710 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C711 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C712 9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C713 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C714 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C715 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C716 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C717 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C718 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C719 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C720 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C721 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C722 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C723 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C724 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C725 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C726 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C727 9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C728 9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C729 9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C730 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C731 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C732 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C733 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C734 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C735 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C736 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C737 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C738 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C739 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C740 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C741 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C742 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C743 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C744 9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C745 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C746 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C747 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C748 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C749 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C750 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C751 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C752 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C753 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C754 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C755 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C756 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C757 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C758 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C759 9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C760 9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C761 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C762 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C763 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C764 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C765 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C766 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C767 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C768 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C769 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C770 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C771 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C772 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C773 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C774 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C775 9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C776 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C777 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C778 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C779 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C780 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C781 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C782 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C783 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C784 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C785 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C786 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C787 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C788 m1_31884_48# VSUBS 2.82fF
C789 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C790 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C791 9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C792 9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C793 9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C794 9good_0/8good_1/7good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C795 9good_0/8good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C796 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C797 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C798 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C799 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C800 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C801 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C802 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C803 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C804 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C805 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C806 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C807 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C808 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C809 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C810 9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C811 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C812 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C813 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C814 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C815 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C816 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C817 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C818 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C819 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C820 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C821 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C822 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C823 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C824 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C825 9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C826 9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C827 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C828 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C829 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C830 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C831 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C832 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C833 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C834 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C835 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C836 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C837 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C838 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C839 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C840 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C841 9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C842 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C843 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C844 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C845 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C846 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C847 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C848 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C849 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C850 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C851 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C852 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C853 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C854 m1_26760_28# VSUBS 2.60fF
C855 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C856 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C857 9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C858 9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C859 9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C860 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C861 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C862 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C863 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C864 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C865 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C866 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C867 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C868 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C869 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C870 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C871 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C872 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C873 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C874 9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C875 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C876 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C877 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C878 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C879 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C880 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C881 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C882 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C883 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C884 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C885 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C886 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C887 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C888 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C889 9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C890 9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C891 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C892 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C893 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C894 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C895 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C896 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C897 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C898 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C899 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C900 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C901 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C902 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C903 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C904 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C905 9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C906 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C907 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C908 9good_0/m1_32342_44672# VSUBS 178.26fF
C909 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C910 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C911 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C912 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C913 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C914 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C915 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C916 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C917 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C918 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C919 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C920 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C921 9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C922 9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C923 9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C924 9good_0/8good_1/7good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C925 9good_0/8good_1/m1_8774_43264# VSUBS 5.31fF
C926 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C927 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C928 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C929 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C930 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C931 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C932 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C933 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C934 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C935 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C936 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C937 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C938 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C939 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C940 9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C941 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C942 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C943 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C944 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C945 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C946 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C947 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C948 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C949 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C950 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C951 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C952 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C953 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C954 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C955 9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C956 9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C957 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C958 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C959 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C960 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C961 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C962 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C963 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C964 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C965 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C966 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C967 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C968 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C969 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C970 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C971 9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C972 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C973 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C974 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C975 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C976 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C977 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C978 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C979 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C980 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C981 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C982 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C983 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C984 m1_16966_2# VSUBS 2.60fF
C985 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C986 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C987 9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C988 9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C989 9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C990 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C991 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C992 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C993 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C994 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C995 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C996 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C997 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C998 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C999 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1000 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1001 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1002 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1003 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1004 9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1005 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1006 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1007 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1008 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1009 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1010 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1011 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1012 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1013 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1014 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1015 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1016 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1017 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1018 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1019 9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1020 9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1021 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1022 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1023 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1024 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1025 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1026 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1027 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1028 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1029 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1030 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1031 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1032 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1033 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1034 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1035 9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1036 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1037 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1038 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1039 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1040 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1041 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1042 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1043 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1044 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1045 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1046 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1047 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1048 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1049 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1050 9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1051 9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1052 9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1053 9good_0/8good_0/7good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1054 9good_0/8good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1055 D7 VSUBS 29.31fF
C1056 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1057 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1058 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1059 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1060 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1061 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1062 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1063 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1064 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1065 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1066 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1067 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1068 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1069 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1070 9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1071 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1072 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1073 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1074 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1075 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1076 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1077 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1078 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1079 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1080 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1081 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1082 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1083 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1084 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1085 9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1086 9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1087 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1088 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1089 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1090 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1091 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1092 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1093 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1094 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1095 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1096 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1097 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1098 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1099 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1100 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1101 9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1102 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1103 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1104 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1105 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1106 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1107 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1108 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1109 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1110 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1111 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1112 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1113 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1114 m1_6754_8# VSUBS 2.85fF
C1115 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1116 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1117 9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1118 9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1119 9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1120 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1121 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1122 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1123 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1124 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1125 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1126 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1127 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1128 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1129 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1130 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1131 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1132 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1133 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1134 9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1135 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1136 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1137 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1138 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1139 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1140 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1141 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1142 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1143 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1144 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1145 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1146 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1147 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1148 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1149 9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1150 9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1151 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1152 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1153 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1154 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1155 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1156 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1157 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1158 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1159 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1160 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1161 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1162 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1163 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1164 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1165 9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1166 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1167 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1168 D0 VSUBS 352.22fF
C1169 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1170 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1171 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1172 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1173 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1174 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# VSUBS 2.05fF
C1175 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# VSUBS 2.05fF
C1176 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# VSUBS 2.05fF
C1177 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# VSUBS 2.05fF
C1178 D1 VSUBS 16.88fF
C1179 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# VSUBS 2.05fF
C1180 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1181 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1182 9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1183 D3 VSUBS 41.95fF
C1184 9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1185 9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1186 9good_0/8good_0/7good_0/Sw-1_0/li_29_719# VSUBS 2.05fF
C1187 9good_0/8good_0/m1_8774_43264# VSUBS 5.31fF
C1188 D6 VSUBS 13.17fF








valpha  VREF Gnd 3.3
vbeta  VDD Gnd 3.3
vzero D0 Gnd pulse(0 1.8 0.1m 60p 60p 0.1m 0.2m)
vone  D1 Gnd pulse(0 1.8 0.2m 60p 60p 0.2m 0.4m)
vtwo  D2 Gnd pulse(0 1.8 0.4m 60p 60p 0.4m 0.8m)
vthree D3 Gnd pulse(0 1.8 0.8m 60p 60p 0.8m 1.6m)
vfour D4 Gnd pulse (0 1.8 1.6m 60p 60p 1.6m 3.2m)
vfive D5 Gnd pulse (0 1.8 3.2m 60p 60p 3.2m 6.4m)
vsix D6 Gnd pulse (0 1.8 6.4m 60p 60p 6.4m 12.8m)
vseven D7 Gnd pulse (0 1.8 12.8m 60p 60p 12.8m 25.6m)
veight D8 Gnd pulse (0 1.8 25.6m 60p 60p 25.6m 51.2m)
vnine D9 Gnd pulse (0 1.8 51.2m 60p 60p 51.2m 102.4m)
.tran 0.01m 102.4m
.control
run

plot V(Y) V(D0)

.endc
.end
