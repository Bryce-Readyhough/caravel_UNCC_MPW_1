* SPICE3 file created from user_project_wrapper.ext - technology: sky130A

.option scale=0.005

* from online
* DC source for current measure
Vdd vdda1 gnd DC 0.7V
Vgnd vssa1 gnd DC 0.0V
Vth analog_io[10] gnd DC 0.1V
Vk analog_io[9] gnd DC 0.15V
Vw analog_io[11] gnd DC 0.18V
Vr analog_io[8] gnd DC 0.25V
Vau analog_io[12] gnd DC 0.7V
Vad analog_io[7] gnd DC 0.0V

Vdd_aux vdda2 gnd DC 1.8V
Ibias analog_io[6] gnd DC 1n

Vsel analog_io[19] gnd DC 1.8V
Vsyn0 analog_io[13] gnd DC 0.7V
Vsyn1 analog_io[14] gnd DC 0.426V


* Vdd VPWR gnd DC 0.7V
* Vgnd VGND gnd DC 0.0V
* Vth vth gnd DC 0.1V
* Vk vk gnd DC 0.15V
* Vw vw gnd DC 0.01V
* Vr vr gnd DC 0.37V
* Vau vau gnd DC 0.08V
* Vad vad gnd DC 0.25V

Idc vdd analog_io[24] DC 10p

.subckt sky130_fd_pr__nfet_01v8_j74adr VSUBS a_109_249# a_109_337# a_21_289#
X0 a_109_337# a_21_289# a_109_249# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_htftno VSUBS w_n187_n133# a_n184_n57# a_n87_n9# a_n87_n97#
X0 a_n87_n9# a_n184_n57# a_n87_n97# w_n187_n133# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_h5gdbm VSUBS a_n101_295# a_n13_343# a_n13_255#
X0 a_n13_343# a_n101_295# a_n13_255# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_dma3uj VSUBS a_n57_109# a_31_157# a_31_69#
X0 a_31_157# a_n57_109# a_31_69# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_hf7xew VSUBS w_n109_n123# a_n106_n47# a_n9_1# a_n9_n87#
X0 a_n9_1# a_n106_n47# a_n9_n87# w_n109_n123# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_b4l3oq VSUBS a_n11_n3# a_n11_n91# w_n111_n127# a_n108_n51#
X0 a_n11_n3# a_n108_n51# a_n11_n91# w_n111_n127# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_k0ujpa VSUBS a_n151_n105# a_n151_n17# w_n251_n141#
+ a_n248_n65#
X0 a_n151_n17# a_n248_n65# a_n151_n105# w_n251_n141# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lz0viw VSUBS a_n55_313# a_n25_343# a_n25_255#
X0 a_n25_343# a_n55_313# a_n25_255# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt Sw-1 VSUBS li_402_584# w_10_596# w_6_312# li_762_210# w_928_594# w_1442_592#
Xsky130_fd_pr__nfet_01v8_j74adr_0 VSUBS VSUBS li_29_719# li_402_584# sky130_fd_pr__nfet_01v8_j74adr
Xsky130_fd_pr__pfet_01v8_htftno_0 VSUBS w_928_594# li_29_719# w_928_594# w_1442_592#
+ sky130_fd_pr__pfet_01v8_htftno
Xsky130_fd_pr__nfet_01v8_h5gdbm_0 VSUBS li_29_719# w_1442_592# li_762_210# sky130_fd_pr__nfet_01v8_h5gdbm
Xsky130_fd_pr__nfet_01v8_dma3uj_0 VSUBS li_29_719# li_126_470# VSUBS sky130_fd_pr__nfet_01v8_dma3uj
Xsky130_fd_pr__pfet_01v8_hf7xew_0 VSUBS w_10_596# li_29_719# w_10_596# li_126_470#
+ sky130_fd_pr__pfet_01v8_hf7xew
Xsky130_fd_pr__pfet_01v8_b4l3oq_0 VSUBS w_10_596# li_29_719# w_10_596# li_402_584#
+ sky130_fd_pr__pfet_01v8_b4l3oq
Xsky130_fd_pr__pfet_01v8_k0ujpa_0 VSUBS li_762_210# w_1442_592# w_1442_592# li_126_470#
+ sky130_fd_pr__pfet_01v8_k0ujpa
Xsky130_fd_pr__nfet_01v8_lz0viw_0 VSUBS li_126_470# w_928_594# w_1442_592# sky130_fd_pr__nfet_01v8_lz0viw
.ends

.subckt sky130_fd_pr__pfet_01v8_owy61o VSUBS a_n73_n61# w_n109_n123# a_15_n61# a_n33_54#
X0 a_15_n61# a_n33_54# a_n73_n61# w_n109_n123# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_63vi9a VSUBS a_15_n11# a_n33_n99# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt one-way VSUBS li_12_16# w_n37_405# li_100_394#
Xsky130_fd_pr__pfet_01v8_owy61o_0 VSUBS li_12_16# w_n37_405# li_100_394# li_100_394#
+ sky130_fd_pr__pfet_01v8_owy61o
Xsky130_fd_pr__nfet_01v8_63vi9a_0 VSUBS li_100_394# li_12_16# li_12_16# sky130_fd_pr__nfet_01v8_63vi9a
.ends

.subckt sky130_fd_pr__nfet_01v8_8mr83b VSUBS a_n73_n42# a_n15_n68# a_15_n42#
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_ykwexw VSUBS a_n73_n42# w_n109_n104# a_n15_n68# a_15_n42#
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt inverter in out vdd vss
Xsky130_fd_pr__nfet_01v8_8mr83b_0 vss vss in out sky130_fd_pr__nfet_01v8_8mr83b
Xsky130_fd_pr__pfet_01v8_ykwexw_0 vss vdd vdd in out sky130_fd_pr__pfet_01v8_ykwexw
.ends

* .subckt sky130_fd_bs_flash__special_sonosfet_star_ocehe0 VSUBS a_15_n11# a_n33_n99#
* + dw_n429_n439# a_n73_n11#
* X0 a_15_n11# a_n33_n99# a_n73_n11# VSUBS sky130_fd_bs_flash__special_sonosfet_star w=420000u l=150000u
* .ends
* 
* .subckt T-cell gate drain source body sky130_fd_bs_flash__special_sonosfet_star_ocehe0_0/dw_n429_n439#
* Xsky130_fd_bs_flash__special_sonosfet_star_ocehe0_0 body source gate sky130_fd_bs_flash__special_sonosfet_star_ocehe0_0/dw_n429_n439#
* + drain sky130_fd_bs_flash__special_sonosfet_star_ocehe0
* .ends
* 
* .subckt x2-array WL0 WL1 BL0 SL0 BL1 SL1 body nwell body SL1 BL1 BL0 SL0 SL1 body
* + BL1 SL0 body BL0
* X1T-cell_0[0|0] WL1 BL0 SL0 body nwell T-cell
* X1T-cell_0[1|0] WL0 BL0 SL0 body nwell T-cell
* X1T-cell_0[0|1] WL1 BL1 SL1 body nwell T-cell
* X1T-cell_0[1|1] WL0 BL1 SL1 body nwell T-cell
* .ends

.subckt sky130_fd_pr__nfet_01v8_r0atdz VSUBS a_n40_n107# a_n98_n81# a_40_n81#
X0 a_40_n81# a_n40_n107# a_n98_n81# VSUBS sky130_fd_pr__nfet_01v8 w=500000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4pknhj VSUBS a_n98_n86# w_n134_n148# a_40_n86# a_n40_n112#
X0 a_40_n86# a_n40_n112# a_n98_n86# w_n134_n148# sky130_fd_pr__pfet_01v8 w=500000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4ujh9u VSUBS w_n144_n198# a_n50_n162# a_n108_n136#
+ a_50_n136#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_01v8 w=1e+06u l=500000u
.ends

.subckt pmos-diff-amp in_1 in_2 out i_bias vdd vss
Xsky130_fd_pr__nfet_01v8_r0atdz_0 vss m1_91_n137# m1_91_n137# vss sky130_fd_pr__nfet_01v8_r0atdz
Xsky130_fd_pr__nfet_01v8_r0atdz_1 vss m1_91_n137# vss out sky130_fd_pr__nfet_01v8_r0atdz
Xsky130_fd_pr__pfet_01v8_4pknhj_0 vss m1_91_n137# vdd li_184_186# in_1 sky130_fd_pr__pfet_01v8_4pknhj
Xsky130_fd_pr__pfet_01v8_4ujh9u_0 vss vdd i_bias li_184_186# vdd sky130_fd_pr__pfet_01v8_4ujh9u
Xsky130_fd_pr__pfet_01v8_4pknhj_1 vss li_184_186# vdd out in_2 sky130_fd_pr__pfet_01v8_4pknhj
Xsky130_fd_pr__pfet_01v8_4ujh9u_1 vss vdd i_bias vdd i_bias sky130_fd_pr__pfet_01v8_4ujh9u
.ends

.subckt sky130_fd_pr__nfet_01v8_dlksd1 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_s3efqo VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lca7f7 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_u061qr VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_h2n75u VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_zt2j7p VSUBS a_n98_n120# a_n40_n146# a_40_n120# w_n134_n182#
X0 a_40_n120# a_n40_n146# a_n98_n120# w_n134_n182# sky130_fd_pr__pfet_01v8 w=1.2e+06u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ckptud VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_2vaynq VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_wpylm8 VSUBS a_n388_n400# a_n330_n426# a_330_n400#
X0 a_330_n400# a_n330_n426# a_n388_n400# VSUBS sky130_fd_pr__nfet_01v8 w=4e+06u l=3.3e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_9i6r5e VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_9hqhhq VSUBS a_n498_n500# a_n440_n526# a_440_n500#
X0 a_440_n500# a_n440_n526# a_n498_n500# VSUBS sky130_fd_pr__nfet_01v8 w=5e+06u l=4.4e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_h43ndc VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_6z4qh8 VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_tb02ql VSUBS a_n618_n800# a_n560_n826# a_560_n800#
X0 a_560_n800# a_n560_n826# a_n618_n800# VSUBS sky130_fd_pr__nfet_01v8 w=8e+06u l=5.6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_zgaw3c VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt neuron-labeled VPWR VGND vth vk vw vr vau vad v u# a# axon
XM10 VGND VGND vad a# sky130_fd_pr__nfet_01v8_dlksd1
XM11 VGND v a# VGND sky130_fd_pr__nfet_01v8_s3efqo
XM1 VGND a_35_1497# v vth sky130_fd_pr__nfet_01v8_lca7f7
XM2 VGND a_35_1497# VPWR VPWR a_35_1497# sky130_fd_pr__pfet_01v8_u061qr
XM3 VGND a_35_1497# VPWR VPWR v sky130_fd_pr__pfet_01v8_h2n75u
XM4 VGND VPWR a_35_1497# axon VPWR sky130_fd_pr__pfet_01v8_zt2j7p
XM5 VGND VGND a_35_1497# axon sky130_fd_pr__nfet_01v8_ckptud
XM6 VGND vw axon VPWR u# sky130_fd_pr__pfet_01v8_2vaynq
XCu VGND VGND u# VGND sky130_fd_pr__nfet_01v8_wpylm8
XM7 VGND VGND vr u# sky130_fd_pr__nfet_01v8_9i6r5e
XCv VGND VGND v VGND sky130_fd_pr__nfet_01v8_9hqhhq
XM8 VGND v u# VGND sky130_fd_pr__nfet_01v8_h43ndc
XM9 VGND vau axon VPWR a# sky130_fd_pr__pfet_01v8_6z4qh8
XCa VGND VGND a# VGND sky130_fd_pr__nfet_01v8_tb02ql
XMk VGND v vk VGND sky130_fd_pr__nfet_01v8_zgaw3c
.ends

.subckt neuron-labeled-extended-opamp v u a vau vw vth vk vr vad vdd vss axon i_bias
+ v_buff u_buff a_buff axon_buff vdd_aux vss vdd v vss
Xpmos-diff-amp_0 v v_buff v_buff i_bias vdd_aux vss pmos-diff-amp
Xpmos-diff-amp_1 u u_buff u_buff i_bias vdd_aux vss pmos-diff-amp
Xpmos-diff-amp_2 a a_buff a_buff i_bias vdd_aux vss pmos-diff-amp
Xpmos-diff-amp_3 axon axon_buff axon_buff i_bias vdd_aux vss pmos-diff-amp
Xneuron-labeled_0 vdd vss vth vk vw vr vau vad v u a axon neuron-labeled
.ends

.subckt sky130_fd_pr__nfet_01v8_5mkfxl VSUBS a_n73_n42# a_15_n42# a_n33_n130#
X0 a_15_n42# a_n33_n130# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_pa2hmj VSUBS a_n33_n177# a_15_n80# w_n109_n180# a_n73_n80#
X0 a_15_n80# a_n33_n177# a_n73_n80# w_n109_n180# sky130_fd_pr__pfet_01v8 w=800000u l=150000u
.ends

.subckt pass-gate clk clk_bar v_in v_out v_newll v_sub v_out
Xsky130_fd_pr__nfet_01v8_5mkfxl_0 v_sub v_out v_in clk sky130_fd_pr__nfet_01v8_5mkfxl
Xsky130_fd_pr__pfet_01v8_pa2hmj_0 v_sub clk_bar v_out v_newll v_in sky130_fd_pr__pfet_01v8_pa2hmj
.ends

.subckt pass-gate-inv-2 in_1 in_2 clk clk_bar out vdd vss vss vdd clk out in_1 clk
+ vss vss
Xinverter_0 clk clk_bar vdd vss inverter
Xpass-gate_0 clk clk_bar in_1 out vdd vss out pass-gate
Xpass-gate_1 clk_bar clk in_2 out vdd vss out pass-gate
.ends

.subckt chip-w-opamp i_bias vad vr vk vth vw vau vsyn0 vsyn1 vdd vss vdd_aux sel v_syn
+ u_syn a_syn axon_syn v_buff u_buff a_buff axon_buff WL0 WL1 BL0 SL0 BL1 SL1 i_in
+ nwell vdd_aux vss BL0 BL1 SL0 vdd_aux BL0 vdd_aux BL1 WL0 BL0 SL1 SL0 BL1 SL1
Xone-way_0 vss inverter_0/out vdd neuron-labeled-extended-opamp_0/v one-way
Xone-way_1 vss inverter_1/out vdd neuron-labeled-extended-opamp_1/v one-way
Xinverter_0 vsyn0 inverter_0/out vdd vss inverter
Xinverter_1 vsyn1 inverter_1/out vdd vss inverter
* X2x2-array_0 WL0 WL1 BL0 SL0 BL1 SL1 vss nwell vss SL1 BL1 BL0 SL0 SL1 vss BL1 SL0
* + vss BL0 x2-array
Xneuron-labeled-extended-opamp_0 neuron-labeled-extended-opamp_0/v neuron-labeled-extended-opamp_0/u
+ neuron-labeled-extended-opamp_0/a vau vw vth vk vr vad vdd vss neuron-labeled-extended-opamp_0/axon
+ i_bias pass-gate-inv-2_0/in_2 pass-gate-inv-2_1/in_2 pass-gate-inv-2_2/in_2 pass-gate-inv-2_3/in_2
+ vdd_aux vss vdd neuron-labeled-extended-opamp_0/v vss neuron-labeled-extended-opamp
Xneuron-labeled-extended-opamp_1 neuron-labeled-extended-opamp_1/v neuron-labeled-extended-opamp_1/u
+ neuron-labeled-extended-opamp_1/a vau vw vth vk vr vad vdd vss neuron-labeled-extended-opamp_1/axon
+ i_bias pass-gate-inv-2_0/in_1 pass-gate-inv-2_1/in_1 pass-gate-inv-2_2/in_1 pass-gate-inv-2_3/in_1
+ vdd_aux vss vdd neuron-labeled-extended-opamp_1/v vss neuron-labeled-extended-opamp
Xneuron-labeled-extended-opamp_2 i_in neuron-labeled-extended-opamp_2/u neuron-labeled-extended-opamp_2/a
+ vau vw vth vk vr vad vdd vss neuron-labeled-extended-opamp_2/axon i_bias v_buff
+ u_buff a_buff axon_buff vdd_aux vss vdd i_in vss neuron-labeled-extended-opamp
Xpass-gate-inv-2_0 pass-gate-inv-2_0/in_1 pass-gate-inv-2_0/in_2 sel pass-gate-inv-2_0/clk_bar
+ v_syn vdd_aux vss vss vdd_aux sel v_syn pass-gate-inv-2_0/in_1 sel vss vss pass-gate-inv-2
Xpass-gate-inv-2_1 pass-gate-inv-2_1/in_1 pass-gate-inv-2_1/in_2 sel pass-gate-inv-2_1/clk_bar
+ u_syn vdd_aux vss vss vdd_aux sel u_syn pass-gate-inv-2_1/in_1 sel vss vss pass-gate-inv-2
Xpass-gate-inv-2_2 pass-gate-inv-2_2/in_1 pass-gate-inv-2_2/in_2 sel pass-gate-inv-2_2/clk_bar
+ a_syn vdd_aux vss vss vdd_aux sel a_syn pass-gate-inv-2_2/in_1 sel vss vss pass-gate-inv-2
Xpass-gate-inv-2_3 pass-gate-inv-2_3/in_1 pass-gate-inv-2_3/in_2 sel pass-gate-inv-2_3/clk_bar
+ axon_syn vdd_aux vss vss vdd_aux sel axon_syn pass-gate-inv-2_3/in_1 sel vss vss
+ pass-gate-inv-2
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[29]
+ analog_io[2] analog_io[30] analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7]
+ analog_io[8] analog_io[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] user_clock2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2
X0 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5 vdda1 io_in[5] 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X7 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X9 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X10 10good_0/9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X11 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X12 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X13 vdda1 io_in[4] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X14 10good_0/9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X15 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X16 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X17 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X18 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X19 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X20 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X21 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X22 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X23 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X24 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X25 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X26 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X27 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X28 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X29 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X30 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X31 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X32 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X33 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X34 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X35 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X36 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X37 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X38 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X39 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X40 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X41 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X42 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X43 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X44 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X45 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X46 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X47 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X48 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X49 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X50 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X51 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X52 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X53 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X54 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X55 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R0 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R2 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R3 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X56 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X57 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X58 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X59 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X60 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X61 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X62 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X63 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X64 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X65 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X66 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X67 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X68 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X69 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X70 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X71 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X72 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X73 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X74 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X75 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X76 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X77 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X78 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X79 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R4 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R5 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R6 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R7 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X80 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X81 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X82 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X83 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X84 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X85 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X86 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X87 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X88 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X89 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X90 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_1684_72# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X91 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X92 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X93 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X94 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_1684_72# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X95 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X96 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X97 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X98 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X99 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X100 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X101 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X102 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X103 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X104 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X105 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X106 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X107 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X108 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X109 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X110 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X111 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R8 10good_0/m1_1684_72# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R9 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R10 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R11 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X112 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X113 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X114 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X115 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X116 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X117 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X118 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X119 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X120 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X121 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X122 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X123 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X124 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X125 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X126 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X127 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X128 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X129 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X130 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X131 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X132 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X133 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X134 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X135 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R12 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R13 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R14 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R15 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X136 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X137 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X138 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X139 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X140 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X141 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X142 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X143 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X144 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X145 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X146 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X147 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X148 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X149 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X150 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X151 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X152 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X153 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X154 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X155 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X156 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X157 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X158 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X159 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X160 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X161 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X162 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X163 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X164 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X165 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X166 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X167 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X168 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X169 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X170 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X171 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X172 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X173 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X174 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X175 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R16 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R17 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R18 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R19 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X176 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X177 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X178 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X179 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X180 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X181 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X182 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X183 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X184 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X185 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X186 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X187 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X188 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X189 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X190 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X191 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X192 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X193 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X194 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X195 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X196 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X197 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X198 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X199 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R20 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R21 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R22 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R23 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X200 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X201 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X202 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X203 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X204 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X205 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X206 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X207 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X208 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X209 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X210 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X211 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X212 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X213 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X214 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X215 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X216 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X217 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X218 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X219 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X220 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X221 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X222 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X223 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X224 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X225 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X226 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X227 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X228 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X229 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X230 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X231 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R24 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R25 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R26 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R27 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X232 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X233 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X234 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X235 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X236 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X237 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X238 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X239 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X240 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X241 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X242 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X243 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X244 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X245 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X246 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X247 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X248 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X249 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X250 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X251 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X252 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X253 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X254 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X255 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R28 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R29 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R30 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R31 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X256 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X257 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X258 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X259 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X260 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X261 vdda1 io_in[4] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X262 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X263 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X264 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X265 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X266 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X267 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X268 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X269 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X270 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X271 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X272 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X273 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X274 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X275 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X276 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X277 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X278 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X279 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X280 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X281 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X282 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X283 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X284 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X285 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X286 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X287 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X288 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X289 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X290 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X291 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X292 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X293 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X294 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X295 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X296 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X297 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X298 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X299 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X300 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X301 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X302 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X303 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R32 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R33 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R34 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R35 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X304 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X305 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X306 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X307 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X308 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X309 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X310 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X311 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X312 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X313 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X314 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X315 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X316 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X317 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X318 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X319 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X320 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X321 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X322 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X323 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X324 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X325 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X326 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X327 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R36 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R37 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R38 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R39 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X328 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X329 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X330 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X331 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X332 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X333 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X334 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X335 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X336 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X337 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X338 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X339 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X340 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X341 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X342 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/m1_14_20144# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X343 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X344 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X345 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X346 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X347 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X348 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X349 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X350 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X351 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X352 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X353 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X354 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X355 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X356 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X357 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X358 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X359 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R40 10good_0/9good_0/8good_0/7good_0/6good_0/m1_14_20144# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R41 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R42 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R43 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X360 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X361 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X362 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X363 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X364 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X365 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X366 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X367 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X368 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X369 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X370 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X371 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X372 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X373 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X374 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X375 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X376 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X377 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X378 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X379 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X380 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X381 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X382 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X383 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R44 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R45 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R46 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R47 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X384 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X385 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X386 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X387 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X388 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X389 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X390 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X391 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X392 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X393 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X394 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X395 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X396 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X397 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X398 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X399 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X400 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X401 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X402 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X403 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X404 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X405 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X406 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X407 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X408 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X409 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X410 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X411 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X412 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X413 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X414 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X415 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X416 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X417 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X418 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X419 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X420 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X421 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X422 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X423 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R48 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R49 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R50 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R51 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X424 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X425 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X426 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X427 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X428 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X429 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X430 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X431 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X432 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X433 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X434 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X435 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X436 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X437 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X438 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X439 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X440 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X441 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X442 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X443 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X444 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X445 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X446 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X447 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R52 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R53 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R54 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# vdda1 sky130_fd_pr__res_generic_po w=66 l=342
R55 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X448 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X449 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X450 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X451 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X452 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X453 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X454 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X455 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X456 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X457 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X458 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X459 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X460 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X461 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X462 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X463 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X464 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X465 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X466 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X467 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X468 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X469 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X470 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X471 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X472 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X473 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X474 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X475 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X476 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X477 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X478 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X479 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R56 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R57 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R58 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R59 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X480 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X481 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X482 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X483 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X484 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X485 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X486 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X487 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X488 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X489 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X490 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X491 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X492 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X493 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X494 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X495 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X496 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X497 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X498 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X499 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X500 vdda1 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X501 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X502 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X503 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R60 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R61 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R62 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R63 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X504 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_29_719# io_in[6] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X505 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/m1_8774_43264# 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X506 10good_0/9good_0/8good_0/m1_8774_43264# 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X507 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X508 vdda1 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X509 vdda1 io_in[6] 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X510 10good_0/9good_0/8good_0/m1_8774_43264# 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# 10good_0/9good_0/8good_0/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X511 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# 10good_0/9good_0/8good_0/7good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/m1_8774_43264# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X512 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X513 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X514 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X515 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X516 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X517 vdda1 io_in[5] 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X518 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X519 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X520 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X521 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X522 10good_0/9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X523 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X524 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X525 vdda1 io_in[4] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X526 10good_0/9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X527 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X528 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X529 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X530 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X531 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X532 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X533 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X534 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X535 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X536 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X537 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X538 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X539 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X540 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X541 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X542 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X543 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X544 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X545 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X546 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X547 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X548 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X549 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X550 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X551 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X552 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X553 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X554 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X555 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X556 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X557 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X558 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X559 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X560 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X561 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X562 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X563 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X564 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X565 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X566 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X567 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R64 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R65 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R66 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R67 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X568 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X569 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X570 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X571 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X572 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X573 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X574 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X575 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X576 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X577 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X578 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X579 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X580 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X581 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X582 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X583 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X584 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X585 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X586 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X587 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X588 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X589 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X590 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X591 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R68 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R69 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R70 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R71 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X592 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X593 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X594 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X595 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X596 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X597 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X598 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X599 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X600 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X601 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X602 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_6754_8# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X603 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X604 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X605 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X606 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_6754_8# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X607 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X608 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X609 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X610 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X611 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X612 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X613 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X614 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X615 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X616 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X617 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X618 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X619 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X620 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X621 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X622 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X623 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R72 10good_0/m1_6754_8# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R73 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R74 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R75 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X624 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X625 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X626 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X627 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X628 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X629 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X630 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X631 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X632 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X633 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X634 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X635 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X636 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X637 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X638 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X639 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X640 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X641 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X642 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X643 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X644 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X645 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X646 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X647 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R76 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R77 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R78 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R79 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X648 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X649 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X650 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X651 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X652 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X653 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X654 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X655 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X656 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X657 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X658 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X659 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X660 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X661 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X662 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X663 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X664 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X665 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X666 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X667 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X668 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X669 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X670 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X671 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X672 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X673 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X674 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X675 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X676 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X677 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X678 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X679 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X680 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X681 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X682 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X683 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X684 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X685 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X686 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X687 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R80 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R81 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R82 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R83 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X688 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X689 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X690 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X691 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X692 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X693 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X694 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X695 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X696 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X697 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X698 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X699 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X700 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X701 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X702 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X703 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X704 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X705 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X706 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X707 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X708 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X709 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X710 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X711 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R84 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R85 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R86 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R87 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X712 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X713 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X714 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X715 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X716 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X717 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X718 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X719 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X720 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X721 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X722 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X723 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X724 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X725 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X726 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X727 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X728 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X729 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X730 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X731 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X732 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X733 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X734 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X735 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X736 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X737 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X738 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X739 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X740 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X741 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X742 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X743 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R88 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R89 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R90 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R91 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X744 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X745 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X746 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X747 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X748 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X749 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X750 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X751 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X752 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X753 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X754 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X755 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X756 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X757 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X758 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X759 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X760 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X761 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X762 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X763 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X764 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X765 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X766 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X767 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R92 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R93 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R94 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R95 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X768 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X769 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X770 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X771 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X772 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X773 vdda1 io_in[4] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X774 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X775 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X776 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X777 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X778 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X779 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X780 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X781 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X782 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X783 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X784 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X785 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X786 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X787 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X788 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X789 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X790 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X791 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X792 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X793 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X794 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X795 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X796 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X797 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X798 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X799 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X800 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X801 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X802 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X803 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X804 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X805 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X806 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X807 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X808 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X809 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X810 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X811 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X812 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X813 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X814 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X815 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R96 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R97 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R98 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R99 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X816 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X817 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X818 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X819 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X820 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X821 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X822 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X823 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X824 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X825 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X826 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X827 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X828 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X829 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X830 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X831 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X832 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X833 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X834 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X835 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X836 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X837 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X838 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X839 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R100 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R101 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R102 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R103 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X840 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X841 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X842 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X843 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X844 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X845 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X846 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X847 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X848 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X849 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X850 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X851 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X852 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X853 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X854 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/m1_14_20144# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X855 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X856 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X857 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X858 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X859 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X860 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X861 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X862 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X863 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X864 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X865 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X866 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X867 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X868 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X869 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X870 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X871 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R104 10good_0/9good_0/8good_0/7good_0/6good_1/m1_14_20144# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R105 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R106 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R107 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X872 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X873 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X874 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X875 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X876 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X877 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X878 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X879 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X880 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X881 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X882 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X883 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X884 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X885 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X886 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X887 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X888 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X889 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X890 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X891 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X892 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X893 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X894 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X895 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R108 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R109 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R110 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R111 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X896 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X897 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X898 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X899 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X900 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X901 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X902 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X903 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X904 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X905 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X906 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X907 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X908 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X909 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X910 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X911 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X912 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X913 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X914 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X915 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X916 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X917 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X918 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X919 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X920 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X921 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X922 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X923 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X924 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X925 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X926 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X927 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X928 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X929 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X930 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X931 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X932 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X933 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X934 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X935 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R112 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R113 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R114 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R115 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X936 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X937 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X938 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X939 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X940 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X941 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X942 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X943 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X944 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X945 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X946 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X947 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X948 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X949 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X950 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X951 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X952 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X953 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X954 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X955 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X956 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X957 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X958 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X959 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R116 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R117 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R118 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_1684_72# sky130_fd_pr__res_generic_po w=66 l=342
R119 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X960 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X961 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X962 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X963 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X964 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X965 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X966 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X967 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X968 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X969 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X970 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X971 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X972 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X973 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X974 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X975 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X976 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X977 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X978 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X979 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X980 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X981 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X982 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X983 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X984 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X985 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X986 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X987 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X988 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X989 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X990 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X991 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R120 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R121 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R122 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R123 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X992 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X993 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X994 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X995 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X996 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X997 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X998 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X999 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1000 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1001 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1002 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1003 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1004 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1005 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1006 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1007 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1008 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1009 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1010 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1011 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1012 vdda1 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1013 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1014 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1015 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R124 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R125 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R126 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R127 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1016 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1017 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X1018 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1019 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1020 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1021 vdda1 io_in[5] 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1022 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X1023 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1024 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1025 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1026 10good_0/9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1027 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1028 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1029 vdda1 io_in[4] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1030 10good_0/9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X1031 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1032 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1033 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1034 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1035 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1036 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1037 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1038 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X1039 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1040 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1041 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1042 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1043 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1044 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1045 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1046 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1047 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1048 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1049 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1050 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1051 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1052 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1053 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1054 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1055 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1056 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1057 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1058 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1059 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1060 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1061 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1062 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1063 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1064 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1065 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1066 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1067 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1068 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1069 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1070 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1071 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R128 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R129 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R130 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R131 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1072 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1073 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1074 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1075 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1076 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1077 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1078 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1079 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1080 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1081 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1082 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1083 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1084 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1085 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1086 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1087 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1088 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1089 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1090 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1091 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1092 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1093 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1094 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1095 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R132 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R133 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R134 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R135 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1096 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1097 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1098 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1099 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1100 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1101 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1102 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1103 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1104 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1105 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1106 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_11882_62# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1107 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1108 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1109 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1110 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_11882_62# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1111 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1112 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1113 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1114 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1115 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1116 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1117 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1118 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1119 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1120 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1121 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1122 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1123 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1124 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1125 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1126 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1127 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R136 10good_0/m1_11882_62# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R137 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R138 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R139 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1128 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1129 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1130 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1131 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1132 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1133 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1134 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1135 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1136 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1137 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1138 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1139 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1140 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1141 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1142 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1143 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1144 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1145 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1146 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1147 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1148 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1149 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1150 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1151 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R140 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R141 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R142 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R143 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1152 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1153 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1154 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1155 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1156 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1157 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1158 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1159 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1160 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1161 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1162 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1163 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1164 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1165 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1166 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1167 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1168 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1169 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1170 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1171 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1172 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1173 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1174 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1175 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1176 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1177 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1178 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1179 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1180 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1181 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1182 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1183 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1184 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1185 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1186 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1187 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1188 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1189 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1190 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1191 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R144 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R145 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R146 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R147 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1192 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1193 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1194 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1195 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1196 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1197 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1198 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1199 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1200 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1201 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1202 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1203 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1204 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1205 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1206 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1207 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1208 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1209 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1210 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1211 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1212 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1213 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1214 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1215 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R148 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R149 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R150 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R151 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1216 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1217 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1218 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1219 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1220 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1221 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1222 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1223 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1224 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1225 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1226 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1227 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1228 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1229 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1230 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1231 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1232 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1233 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1234 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1235 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1236 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1237 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1238 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1239 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1240 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1241 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1242 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1243 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1244 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1245 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1246 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1247 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R152 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R153 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R154 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R155 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1248 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1249 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1250 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1251 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1252 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1253 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1254 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1255 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1256 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1257 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1258 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1259 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1260 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1261 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1262 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1263 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1264 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1265 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1266 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1267 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1268 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1269 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1270 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1271 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R156 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R157 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R158 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R159 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1272 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1273 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1274 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1275 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1276 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1277 vdda1 io_in[4] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1278 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X1279 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1280 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1281 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1282 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1283 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1284 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1285 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1286 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X1287 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1288 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1289 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1290 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1291 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1292 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1293 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1294 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1295 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1296 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1297 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1298 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1299 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1300 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1301 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1302 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1303 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1304 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1305 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1306 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1307 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1308 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1309 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1310 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1311 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1312 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1313 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1314 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1315 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1316 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1317 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1318 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1319 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R160 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R161 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R162 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R163 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1320 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1321 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1322 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1323 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1324 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1325 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1326 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1327 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1328 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1329 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1330 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1331 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1332 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1333 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1334 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1335 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1336 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1337 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1338 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1339 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1340 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1341 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1342 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1343 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R164 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R165 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R166 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R167 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1344 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1345 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1346 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1347 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1348 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1349 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1350 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1351 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1352 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1353 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1354 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1355 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1356 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1357 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1358 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_14_20144# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1359 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1360 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1361 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1362 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1363 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1364 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1365 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1366 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1367 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1368 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1369 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1370 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1371 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1372 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1373 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1374 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1375 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R168 10good_0/9good_0/8good_0/7good_1/6good_0/m1_14_20144# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R169 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R170 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R171 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1376 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1377 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1378 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1379 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1380 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1381 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1382 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1383 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1384 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1385 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1386 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1387 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1388 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1389 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1390 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1391 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1392 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1393 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1394 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1395 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1396 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1397 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1398 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1399 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R172 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R173 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R174 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R175 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1400 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1401 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1402 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1403 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1404 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1405 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1406 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1407 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1408 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1409 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1410 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1411 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1412 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1413 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1414 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1415 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1416 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1417 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1418 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1419 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1420 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1421 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1422 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1423 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1424 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1425 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1426 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1427 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1428 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1429 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1430 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1431 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1432 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1433 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1434 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1435 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1436 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1437 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1438 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1439 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R176 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R177 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R178 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R179 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1440 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1441 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1442 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1443 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1444 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1445 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1446 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1447 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1448 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1449 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1450 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1451 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1452 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1453 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1454 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1455 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1456 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1457 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1458 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1459 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1460 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1461 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1462 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1463 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R180 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R181 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R182 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_6754_8# sky130_fd_pr__res_generic_po w=66 l=342
R183 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1464 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1465 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1466 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1467 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1468 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1469 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1470 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1471 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1472 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1473 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1474 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1475 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1476 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1477 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1478 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1479 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1480 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1481 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1482 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1483 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1484 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1485 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1486 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1487 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1488 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1489 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1490 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1491 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1492 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1493 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1494 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1495 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R184 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R185 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R186 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R187 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1496 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1497 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1498 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1499 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1500 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1501 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1502 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1503 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1504 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1505 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1506 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1507 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1508 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1509 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1510 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1511 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1512 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1513 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1514 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1515 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1516 vdda1 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1517 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1518 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1519 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R188 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R189 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R190 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R191 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1520 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_29_719# io_in[6] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1521 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/m1_18694_42308# 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X1522 10good_0/9good_0/8good_0/m1_18694_42308# 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1523 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1524 vdda1 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1525 vdda1 io_in[6] 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1526 10good_0/9good_0/8good_0/m1_18694_42308# 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# 10good_0/9good_0/8good_0/m1_18694_42308# sky130_fd_pr__pfet_01v8 w=84 l=30
X1527 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# 10good_0/9good_0/8good_0/7good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/m1_18694_42308# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1528 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1529 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X1530 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1531 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1532 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1533 vdda1 io_in[5] 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1534 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X1535 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1536 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1537 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1538 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1539 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1540 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1541 vdda1 io_in[4] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1542 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X1543 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1544 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1545 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1546 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1547 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1548 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1549 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1550 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X1551 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1552 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1553 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1554 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1555 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1556 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1557 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1558 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1559 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1560 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1561 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1562 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1563 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1564 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1565 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1566 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1567 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1568 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1569 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1570 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1571 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1572 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1573 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1574 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1575 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1576 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1577 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1578 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1579 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1580 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1581 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1582 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1583 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R192 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R193 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R194 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R195 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1584 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1585 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1586 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1587 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1588 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1589 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1590 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1591 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1592 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1593 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1594 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1595 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1596 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1597 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1598 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1599 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1600 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1601 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1602 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1603 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1604 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1605 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1606 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1607 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R196 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R197 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R198 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R199 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1608 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1609 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1610 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1611 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1612 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1613 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1614 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1615 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1616 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1617 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1618 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_16966_2# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1619 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1620 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1621 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1622 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_16966_2# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1623 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1624 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1625 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1626 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1627 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1628 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1629 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1630 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1631 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1632 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1633 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1634 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1635 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1636 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1637 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1638 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1639 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R200 10good_0/m1_16966_2# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R201 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R202 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R203 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1640 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1641 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1642 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1643 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1644 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1645 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1646 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1647 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1648 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1649 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1650 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1651 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1652 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1653 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1654 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1655 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1656 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1657 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1658 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1659 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1660 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1661 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1662 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1663 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R204 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R205 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R206 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R207 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1664 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1665 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1666 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1667 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1668 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1669 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1670 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1671 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1672 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1673 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1674 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1675 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1676 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1677 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1678 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1679 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1680 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1681 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1682 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1683 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1684 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1685 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1686 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1687 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1688 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1689 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1690 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1691 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1692 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1693 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1694 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1695 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1696 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1697 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1698 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1699 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1700 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1701 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1702 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1703 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R208 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R209 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R210 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R211 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1704 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1705 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1706 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1707 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1708 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1709 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1710 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1711 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1712 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1713 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1714 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1715 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1716 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1717 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1718 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1719 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1720 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1721 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1722 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1723 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1724 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1725 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1726 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1727 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R212 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R213 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R214 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R215 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1728 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1729 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1730 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1731 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1732 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1733 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1734 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1735 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1736 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1737 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1738 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1739 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1740 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1741 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1742 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1743 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1744 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1745 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1746 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1747 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1748 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1749 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1750 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1751 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1752 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1753 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1754 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1755 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1756 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1757 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1758 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1759 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R216 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R217 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R218 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R219 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1760 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1761 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1762 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1763 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1764 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1765 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1766 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1767 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1768 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1769 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1770 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1771 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1772 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1773 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1774 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1775 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1776 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1777 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1778 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1779 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1780 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1781 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1782 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1783 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R220 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R221 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R222 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R223 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1784 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1785 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1786 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1787 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1788 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1789 vdda1 io_in[4] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1790 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X1791 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1792 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1793 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1794 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1795 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1796 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1797 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1798 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X1799 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1800 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1801 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1802 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1803 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1804 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1805 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1806 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1807 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1808 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1809 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1810 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1811 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1812 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1813 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1814 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1815 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1816 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1817 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1818 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1819 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1820 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1821 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1822 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1823 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1824 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1825 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1826 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1827 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1828 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1829 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1830 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1831 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R224 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R225 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R226 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R227 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1832 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1833 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1834 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1835 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1836 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1837 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1838 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1839 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1840 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1841 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1842 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1843 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1844 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1845 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1846 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1847 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1848 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1849 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1850 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1851 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1852 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1853 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1854 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1855 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R228 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R229 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R230 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R231 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1856 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1857 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1858 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1859 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1860 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1861 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1862 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1863 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1864 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1865 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1866 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1867 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1868 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1869 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1870 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_14_20144# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1871 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1872 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1873 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1874 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1875 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1876 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1877 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1878 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1879 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1880 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1881 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1882 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1883 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1884 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1885 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1886 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1887 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R232 10good_0/9good_0/8good_0/7good_1/6good_1/m1_14_20144# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R233 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R234 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R235 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1888 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1889 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1890 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1891 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1892 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1893 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1894 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1895 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1896 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1897 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1898 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1899 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1900 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1901 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1902 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1903 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1904 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1905 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1906 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1907 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1908 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1909 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1910 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1911 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R236 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R237 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R238 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R239 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1912 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1913 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1914 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1915 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1916 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1917 vdda1 io_in[3] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1918 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X1919 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1920 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1921 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1922 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1923 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1924 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1925 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1926 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X1927 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1928 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1929 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1930 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1931 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1932 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1933 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1934 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1935 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1936 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1937 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1938 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1939 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1940 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1941 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1942 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1943 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1944 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1945 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1946 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1947 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1948 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1949 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1950 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X1951 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R240 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R241 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R242 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R243 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1952 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1953 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1954 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1955 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1956 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1957 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1958 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1959 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1960 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1961 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1962 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1963 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1964 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1965 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1966 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1967 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1968 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1969 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1970 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1971 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1972 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1973 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1974 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1975 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R244 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R245 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R246 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_11882_62# sky130_fd_pr__res_generic_po w=66 l=342
R247 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X1976 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1977 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X1978 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1979 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1980 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1981 vdda1 io_in[2] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1982 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X1983 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1984 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1985 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X1986 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1987 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1988 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1989 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1990 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X1991 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1992 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1993 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X1994 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1995 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X1996 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1997 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X1998 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X1999 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2000 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2001 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2002 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2003 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2004 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2005 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2006 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2007 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R248 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R249 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R250 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R251 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2008 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2009 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2010 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2011 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2012 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2013 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2014 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2015 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2016 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2017 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2018 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2019 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2020 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2021 vdda1 io_in[0] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2022 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2023 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2024 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2025 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2026 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2027 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2028 vdda1 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2029 vdda1 io_in[1] 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2030 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2031 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R252 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R253 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R254 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R255 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2032 10good_0/9good_0/8good_0/Sw-1_0/li_29_719# io_in[7] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2033 10good_0/9good_0/8good_0/m1_8774_43264# 10good_0/9good_0/8good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_19068_42976# 10good_0/9good_0/8good_0/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X2034 10good_0/9good_0/m1_19068_42976# 10good_0/9good_0/8good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/m1_18694_42308# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2035 10good_0/9good_0/8good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2036 vdda1 10good_0/9good_0/8good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2037 vdda1 io_in[7] 10good_0/9good_0/8good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2038 10good_0/9good_0/m1_19068_42976# 10good_0/9good_0/8good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_0/m1_18694_42308# 10good_0/9good_0/m1_19068_42976# sky130_fd_pr__pfet_01v8 w=84 l=30
X2039 10good_0/9good_0/8good_0/m1_8774_43264# 10good_0/9good_0/8good_0/Sw-1_0/li_126_470# 10good_0/9good_0/m1_19068_42976# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2040 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2041 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2042 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2043 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2044 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2045 vdda1 io_in[5] 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2046 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X2047 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2048 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2049 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2050 10good_0/9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2051 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2052 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2053 vdda1 io_in[4] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2054 10good_0/9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X2055 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2056 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2057 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2058 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2059 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2060 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2061 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2062 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X2063 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2064 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2065 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2066 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2067 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2068 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2069 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2070 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2071 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2072 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2073 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2074 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2075 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2076 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2077 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2078 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2079 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2080 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2081 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2082 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2083 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2084 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2085 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2086 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2087 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2088 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2089 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2090 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2091 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2092 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2093 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2094 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2095 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R256 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R257 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R258 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R259 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2096 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2097 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2098 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2099 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2100 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2101 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2102 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2103 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2104 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2105 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2106 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2107 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2108 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2109 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2110 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2111 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2112 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2113 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2114 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2115 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2116 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2117 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2118 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2119 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R260 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R261 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R262 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R263 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2120 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2121 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2122 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2123 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2124 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2125 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2126 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2127 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2128 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2129 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2130 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_21660_68# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2131 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2132 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2133 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2134 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_21660_68# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2135 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2136 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2137 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2138 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2139 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2140 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2141 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2142 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2143 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2144 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2145 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2146 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2147 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2148 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2149 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2150 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2151 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R264 10good_0/m1_21660_68# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R265 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R266 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R267 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2152 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2153 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2154 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2155 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2156 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2157 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2158 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2159 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2160 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2161 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2162 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2163 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2164 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2165 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2166 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2167 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2168 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2169 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2170 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2171 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2172 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2173 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2174 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2175 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R268 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R269 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R270 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R271 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2176 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2177 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2178 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2179 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2180 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2181 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2182 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2183 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2184 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2185 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2186 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2187 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2188 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2189 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2190 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2191 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2192 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2193 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2194 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2195 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2196 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2197 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2198 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2199 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2200 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2201 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2202 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2203 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2204 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2205 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2206 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2207 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2208 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2209 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2210 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2211 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2212 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2213 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2214 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2215 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R272 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R273 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R274 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R275 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2216 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2217 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2218 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2219 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2220 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2221 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2222 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2223 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2224 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2225 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2226 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2227 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2228 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2229 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2230 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2231 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2232 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2233 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2234 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2235 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2236 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2237 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2238 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2239 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R276 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R277 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R278 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R279 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2240 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2241 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2242 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2243 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2244 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2245 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2246 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2247 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2248 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2249 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2250 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2251 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2252 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2253 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2254 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2255 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2256 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2257 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2258 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2259 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2260 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2261 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2262 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2263 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2264 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2265 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2266 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2267 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2268 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2269 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2270 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2271 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R280 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R281 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R282 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R283 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2272 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2273 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2274 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2275 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2276 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2277 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2278 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2279 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2280 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2281 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2282 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2283 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2284 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2285 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2286 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2287 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2288 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2289 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2290 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2291 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2292 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2293 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2294 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2295 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R284 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R285 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R286 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R287 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2296 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2297 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2298 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2299 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2300 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2301 vdda1 io_in[4] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2302 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2303 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2304 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2305 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2306 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2307 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2308 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2309 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2310 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X2311 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2312 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2313 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2314 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2315 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2316 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2317 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2318 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2319 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2320 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2321 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2322 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2323 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2324 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2325 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2326 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2327 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2328 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2329 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2330 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2331 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2332 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2333 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2334 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2335 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2336 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2337 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2338 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2339 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2340 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2341 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2342 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2343 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R288 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R289 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R290 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R291 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2344 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2345 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2346 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2347 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2348 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2349 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2350 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2351 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2352 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2353 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2354 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2355 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2356 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2357 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2358 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2359 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2360 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2361 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2362 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2363 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2364 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2365 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2366 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2367 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R292 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R293 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R294 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R295 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2368 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2369 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2370 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2371 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2372 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2373 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2374 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2375 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2376 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2377 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2378 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2379 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2380 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2381 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2382 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_14_20144# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2383 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2384 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2385 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2386 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2387 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2388 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2389 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2390 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2391 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2392 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2393 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2394 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2395 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2396 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2397 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2398 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2399 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R296 10good_0/9good_0/8good_1/7good_0/6good_0/m1_14_20144# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R297 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R298 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R299 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2400 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2401 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2402 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2403 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2404 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2405 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2406 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2407 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2408 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2409 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2410 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2411 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2412 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2413 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2414 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2415 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2416 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2417 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2418 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2419 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2420 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2421 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2422 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2423 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R300 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R301 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R302 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R303 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2424 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2425 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2426 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2427 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2428 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2429 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2430 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2431 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2432 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2433 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2434 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2435 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2436 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2437 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2438 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2439 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2440 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2441 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2442 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2443 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2444 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2445 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2446 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2447 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2448 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2449 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2450 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2451 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2452 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2453 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2454 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2455 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2456 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2457 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2458 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2459 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2460 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2461 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2462 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2463 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R304 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R305 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R306 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R307 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2464 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2465 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2466 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2467 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2468 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2469 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2470 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2471 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2472 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2473 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2474 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2475 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2476 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2477 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2478 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2479 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2480 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2481 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2482 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2483 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2484 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2485 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2486 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2487 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R308 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R309 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R310 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_16966_2# sky130_fd_pr__res_generic_po w=66 l=342
R311 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2488 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2489 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2490 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2491 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2492 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2493 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2494 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2495 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2496 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2497 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2498 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2499 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2500 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2501 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2502 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2503 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2504 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2505 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2506 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2507 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2508 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2509 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2510 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2511 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2512 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2513 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2514 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2515 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2516 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2517 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2518 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2519 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R312 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R313 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R314 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R315 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2520 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2521 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2522 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2523 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2524 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2525 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2526 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2527 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2528 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2529 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2530 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2531 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2532 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2533 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2534 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2535 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2536 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2537 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2538 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2539 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2540 vdda1 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2541 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2542 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2543 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R316 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R317 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R318 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R319 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2544 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_29_719# io_in[6] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2545 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/m1_8774_43264# 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X2546 10good_0/9good_0/8good_1/m1_8774_43264# 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2547 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2548 vdda1 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2549 vdda1 io_in[6] 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2550 10good_0/9good_0/8good_1/m1_8774_43264# 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/m1_8436_40544# 10good_0/9good_0/8good_1/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X2551 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# 10good_0/9good_0/8good_1/7good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/m1_8774_43264# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2552 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2553 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/m1_8436_40544# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2554 10good_0/9good_0/8good_1/7good_0/m1_8436_40544# 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2555 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2556 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2557 vdda1 io_in[5] 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2558 10good_0/9good_0/8good_1/7good_0/m1_8436_40544# 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X2559 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2560 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2561 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2562 10good_0/9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2563 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2564 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2565 vdda1 io_in[4] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2566 10good_0/9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X2567 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2568 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2569 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2570 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2571 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2572 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2573 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2574 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X2575 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2576 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2577 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2578 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2579 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2580 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2581 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2582 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2583 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2584 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2585 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2586 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2587 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2588 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2589 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2590 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2591 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2592 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2593 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2594 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2595 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2596 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2597 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2598 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2599 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2600 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2601 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2602 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2603 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2604 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2605 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2606 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2607 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R320 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R321 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R322 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R323 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2608 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2609 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2610 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2611 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2612 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2613 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2614 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2615 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2616 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2617 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2618 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2619 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2620 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2621 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2622 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2623 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2624 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2625 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2626 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2627 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2628 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2629 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2630 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2631 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R324 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R325 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R326 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R327 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2632 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2633 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2634 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2635 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2636 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2637 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2638 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2639 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2640 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2641 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2642 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_26760_28# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2643 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2644 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2645 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2646 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_26760_28# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2647 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2648 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2649 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2650 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2651 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2652 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2653 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2654 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2655 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2656 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2657 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2658 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2659 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2660 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2661 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2662 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2663 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R328 10good_0/m1_26760_28# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R329 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R330 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R331 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2664 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2665 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2666 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2667 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2668 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2669 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2670 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2671 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2672 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2673 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2674 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2675 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2676 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2677 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2678 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2679 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2680 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2681 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2682 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2683 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2684 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2685 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2686 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2687 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R332 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R333 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R334 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R335 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2688 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2689 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2690 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2691 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2692 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2693 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2694 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2695 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2696 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2697 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2698 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2699 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2700 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2701 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2702 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2703 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2704 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2705 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2706 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2707 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2708 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2709 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2710 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2711 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2712 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2713 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2714 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2715 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2716 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2717 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2718 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2719 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2720 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2721 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2722 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2723 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2724 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2725 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2726 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2727 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R336 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R337 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R338 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R339 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2728 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2729 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2730 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2731 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2732 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2733 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2734 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2735 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2736 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2737 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2738 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2739 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2740 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2741 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2742 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2743 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2744 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2745 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2746 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2747 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2748 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2749 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2750 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2751 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R340 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R341 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R342 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R343 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2752 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2753 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2754 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2755 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2756 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2757 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2758 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2759 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2760 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2761 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2762 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2763 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2764 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2765 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2766 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2767 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2768 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2769 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2770 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2771 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2772 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2773 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2774 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2775 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2776 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2777 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2778 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2779 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2780 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2781 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2782 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2783 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R344 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R345 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R346 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R347 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2784 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2785 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2786 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2787 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2788 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2789 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2790 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2791 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2792 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2793 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2794 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2795 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2796 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2797 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2798 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2799 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2800 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2801 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2802 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2803 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2804 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2805 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2806 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2807 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R348 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R349 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R350 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R351 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2808 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2809 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2810 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2811 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2812 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2813 vdda1 io_in[4] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2814 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X2815 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2816 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2817 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2818 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2819 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2820 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2821 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2822 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X2823 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2824 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2825 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2826 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2827 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2828 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2829 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2830 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2831 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2832 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2833 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2834 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2835 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2836 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2837 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2838 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2839 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2840 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2841 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2842 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2843 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2844 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2845 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2846 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2847 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2848 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2849 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2850 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2851 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2852 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2853 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2854 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2855 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R352 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R353 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R354 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R355 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2856 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2857 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2858 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2859 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2860 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2861 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2862 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2863 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2864 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2865 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2866 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2867 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2868 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2869 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2870 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2871 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2872 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2873 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2874 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2875 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2876 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2877 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2878 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2879 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R356 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R357 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R358 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R359 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2880 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2881 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2882 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2883 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2884 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2885 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2886 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X2887 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2888 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2889 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2890 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2891 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2892 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2893 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2894 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_14_20144# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2895 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2896 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2897 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2898 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2899 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2900 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2901 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2902 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2903 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2904 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2905 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2906 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2907 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2908 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2909 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2910 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2911 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R360 10good_0/9good_0/8good_1/7good_0/6good_1/m1_14_20144# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R361 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R362 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R363 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2912 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2913 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2914 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2915 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2916 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2917 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2918 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2919 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2920 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2921 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2922 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2923 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2924 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2925 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2926 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2927 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2928 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2929 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2930 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2931 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2932 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2933 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2934 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2935 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R364 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R365 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R366 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R367 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2936 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2937 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2938 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2939 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2940 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2941 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2942 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X2943 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2944 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2945 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2946 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2947 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2948 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2949 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2950 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X2951 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2952 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2953 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2954 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2955 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2956 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2957 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2958 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2959 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2960 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2961 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2962 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2963 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2964 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2965 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2966 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2967 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2968 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2969 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2970 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2971 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2972 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2973 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2974 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X2975 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R368 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R369 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R370 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R371 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X2976 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2977 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X2978 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2979 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2980 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2981 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2982 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X2983 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2984 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2985 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X2986 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2987 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2988 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2989 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2990 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2991 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2992 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2993 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X2994 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2995 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X2996 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2997 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X2998 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X2999 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R372 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R373 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R374 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_21660_68# sky130_fd_pr__res_generic_po w=66 l=342
R375 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3000 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3001 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3002 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3003 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3004 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3005 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3006 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3007 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3008 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3009 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3010 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3011 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3012 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3013 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3014 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3015 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3016 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3017 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3018 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3019 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3020 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3021 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3022 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3023 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3024 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3025 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3026 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3027 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3028 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3029 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3030 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3031 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R376 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R377 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R378 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R379 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3032 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3033 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3034 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3035 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3036 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3037 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3038 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3039 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3040 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3041 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3042 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3043 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3044 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3045 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3046 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3047 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3048 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3049 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3050 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3051 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3052 vdda1 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3053 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3054 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3055 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R380 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R381 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R382 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R383 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3056 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3057 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X3058 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3059 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3060 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3061 vdda1 io_in[5] 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3062 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X3063 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3064 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3065 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3066 10good_0/9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3067 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3068 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3069 vdda1 io_in[4] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3070 10good_0/9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X3071 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3072 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3073 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3074 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3075 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3076 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3077 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3078 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X3079 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3080 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3081 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3082 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3083 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3084 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3085 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3086 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3087 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3088 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3089 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3090 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3091 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3092 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3093 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3094 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3095 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3096 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3097 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3098 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3099 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3100 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3101 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3102 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3103 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3104 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3105 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3106 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3107 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3108 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3109 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3110 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3111 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R384 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R385 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R386 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R387 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3112 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3113 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3114 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3115 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3116 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3117 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3118 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3119 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3120 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3121 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3122 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3123 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3124 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3125 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3126 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3127 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3128 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3129 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3130 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3131 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3132 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3133 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3134 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3135 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R388 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R389 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R390 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R391 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3136 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3137 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3138 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3139 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3140 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3141 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3142 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3143 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3144 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3145 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3146 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_31884_48# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3147 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3148 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3149 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3150 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_31884_48# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3151 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3152 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3153 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3154 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3155 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3156 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3157 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3158 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3159 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3160 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3161 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3162 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3163 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3164 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3165 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3166 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3167 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R392 10good_0/m1_31884_48# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R393 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R394 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R395 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3168 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3169 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3170 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3171 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3172 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3173 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3174 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3175 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3176 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3177 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3178 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3179 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3180 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3181 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3182 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3183 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3184 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3185 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3186 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3187 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3188 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3189 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3190 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3191 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R396 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R397 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R398 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R399 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3192 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3193 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3194 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3195 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3196 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3197 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3198 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3199 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3200 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3201 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3202 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3203 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3204 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3205 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3206 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3207 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3208 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3209 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3210 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3211 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3212 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3213 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3214 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3215 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3216 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3217 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3218 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3219 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3220 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3221 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3222 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3223 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3224 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3225 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3226 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3227 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3228 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3229 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3230 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3231 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R400 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R401 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R402 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R403 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3232 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3233 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3234 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3235 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3236 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3237 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3238 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3239 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3240 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3241 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3242 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3243 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3244 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3245 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3246 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3247 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3248 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3249 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3250 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3251 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3252 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3253 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3254 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3255 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R404 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R405 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R406 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R407 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3256 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3257 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3258 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3259 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3260 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3261 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3262 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3263 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3264 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3265 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3266 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3267 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3268 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3269 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3270 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3271 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3272 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3273 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3274 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3275 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3276 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3277 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3278 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3279 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3280 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3281 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3282 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3283 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3284 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3285 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3286 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3287 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R408 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R409 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R410 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R411 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3288 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3289 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3290 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3291 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3292 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3293 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3294 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3295 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3296 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3297 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3298 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3299 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3300 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3301 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3302 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3303 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3304 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3305 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3306 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3307 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3308 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3309 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3310 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3311 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R412 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R413 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R414 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R415 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3312 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3313 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3314 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3315 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3316 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3317 vdda1 io_in[4] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3318 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X3319 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3320 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3321 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3322 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3323 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3324 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3325 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3326 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X3327 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3328 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3329 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3330 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3331 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3332 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3333 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3334 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3335 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3336 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3337 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3338 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3339 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3340 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3341 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3342 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3343 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3344 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3345 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3346 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3347 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3348 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3349 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3350 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3351 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3352 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3353 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3354 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3355 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3356 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3357 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3358 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3359 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R416 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R417 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R418 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R419 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3360 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3361 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3362 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3363 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3364 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3365 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3366 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3367 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3368 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3369 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3370 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3371 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3372 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3373 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3374 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3375 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3376 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3377 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3378 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3379 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3380 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3381 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3382 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3383 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R420 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R421 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R422 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R423 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3384 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3385 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3386 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3387 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3388 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3389 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3390 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3391 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3392 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3393 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3394 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3395 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3396 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3397 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3398 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/m1_14_20144# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3399 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3400 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3401 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3402 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3403 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3404 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3405 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3406 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3407 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3408 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3409 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3410 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3411 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3412 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3413 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3414 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3415 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R424 10good_0/9good_0/8good_1/7good_1/6good_0/m1_14_20144# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R425 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R426 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R427 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3416 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3417 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3418 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3419 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3420 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3421 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3422 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3423 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3424 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3425 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3426 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3427 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3428 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3429 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3430 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3431 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3432 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3433 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3434 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3435 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3436 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3437 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3438 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3439 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R428 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R429 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R430 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R431 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3440 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3441 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3442 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3443 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3444 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3445 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3446 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3447 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3448 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3449 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3450 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3451 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3452 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3453 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3454 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3455 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3456 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3457 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3458 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3459 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3460 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3461 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3462 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3463 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3464 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3465 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3466 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3467 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3468 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3469 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3470 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3471 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3472 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3473 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3474 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3475 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3476 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3477 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3478 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3479 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R432 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R433 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R434 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R435 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3480 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3481 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3482 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3483 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3484 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3485 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3486 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3487 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3488 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3489 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3490 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3491 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3492 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3493 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3494 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3495 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3496 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3497 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3498 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3499 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3500 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3501 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3502 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3503 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R436 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R437 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R438 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_26760_28# sky130_fd_pr__res_generic_po w=66 l=342
R439 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3504 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3505 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3506 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3507 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3508 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3509 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3510 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3511 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3512 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3513 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3514 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3515 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3516 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3517 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3518 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3519 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3520 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3521 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3522 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3523 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3524 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3525 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3526 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3527 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3528 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3529 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3530 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3531 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3532 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3533 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3534 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3535 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R440 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R441 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R442 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R443 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3536 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3537 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3538 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3539 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3540 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3541 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3542 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3543 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3544 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3545 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3546 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3547 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3548 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3549 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3550 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3551 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3552 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3553 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3554 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3555 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3556 vdda1 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3557 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3558 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3559 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R444 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R445 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R446 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R447 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3560 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_29_719# io_in[6] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3561 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/m1_18694_42308# 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X3562 10good_0/9good_0/8good_1/m1_18694_42308# 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3563 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3564 vdda1 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3565 vdda1 io_in[6] 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3566 10good_0/9good_0/8good_1/m1_18694_42308# 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# 10good_0/9good_0/8good_1/m1_18694_42308# sky130_fd_pr__pfet_01v8 w=84 l=30
X3567 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# 10good_0/9good_0/8good_1/7good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/m1_18694_42308# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3568 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3569 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X3570 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3571 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3572 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3573 vdda1 io_in[5] 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3574 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X3575 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3576 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3577 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3578 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3579 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3580 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3581 vdda1 io_in[4] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3582 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X3583 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3584 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3585 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3586 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3587 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3588 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3589 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3590 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X3591 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3592 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3593 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3594 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3595 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3596 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3597 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3598 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3599 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3600 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3601 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3602 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3603 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3604 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3605 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3606 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3607 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3608 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3609 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3610 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3611 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3612 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3613 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3614 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3615 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3616 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3617 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3618 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3619 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3620 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3621 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3622 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3623 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R448 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R449 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R450 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R451 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3624 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3625 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3626 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3627 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3628 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3629 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3630 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3631 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3632 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3633 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3634 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3635 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3636 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3637 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3638 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3639 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3640 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3641 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3642 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3643 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3644 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3645 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3646 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3647 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R452 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R453 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R454 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R455 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3648 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3649 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3650 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3651 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3652 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3653 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3654 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3655 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3656 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3657 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3658 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_36912_2# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3659 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3660 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3661 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3662 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_36912_2# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3663 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3664 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3665 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3666 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3667 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3668 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3669 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3670 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3671 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3672 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3673 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3674 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3675 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3676 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3677 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3678 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3679 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R456 10good_0/m1_36912_2# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R457 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R458 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R459 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3680 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3681 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3682 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3683 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3684 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3685 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3686 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3687 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3688 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3689 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3690 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3691 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3692 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3693 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3694 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3695 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3696 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3697 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3698 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3699 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3700 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3701 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3702 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3703 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R460 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R461 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R462 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R463 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3704 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3705 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3706 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3707 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3708 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3709 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3710 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3711 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3712 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3713 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3714 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3715 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3716 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3717 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3718 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3719 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3720 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3721 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3722 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3723 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3724 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3725 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3726 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3727 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3728 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3729 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3730 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3731 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3732 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3733 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3734 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3735 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3736 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3737 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3738 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3739 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3740 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3741 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3742 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3743 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R464 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R465 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R466 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R467 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3744 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3745 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3746 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3747 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3748 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3749 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3750 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3751 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3752 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3753 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3754 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3755 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3756 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3757 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3758 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3759 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3760 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3761 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3762 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3763 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3764 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3765 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3766 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3767 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R468 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R469 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R470 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R471 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3768 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3769 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3770 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3771 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3772 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3773 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3774 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3775 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3776 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3777 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3778 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3779 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3780 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3781 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3782 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3783 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3784 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3785 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3786 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3787 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3788 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3789 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3790 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3791 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3792 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3793 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3794 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3795 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3796 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3797 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3798 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3799 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R472 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R473 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R474 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R475 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3800 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3801 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3802 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3803 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3804 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3805 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3806 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3807 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3808 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3809 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3810 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3811 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3812 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3813 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3814 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3815 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3816 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3817 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3818 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3819 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3820 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3821 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3822 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3823 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R476 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R477 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R478 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R479 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3824 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3825 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3826 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3827 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3828 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3829 vdda1 io_in[4] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3830 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X3831 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3832 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3833 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3834 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3835 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3836 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3837 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3838 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X3839 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3840 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3841 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3842 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3843 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3844 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3845 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3846 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3847 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3848 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3849 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3850 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3851 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3852 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3853 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3854 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3855 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3856 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3857 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3858 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3859 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3860 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3861 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3862 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3863 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3864 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3865 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3866 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3867 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3868 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3869 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3870 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3871 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R480 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R481 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R482 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R483 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3872 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3873 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3874 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3875 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3876 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3877 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3878 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3879 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3880 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3881 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3882 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3883 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3884 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3885 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3886 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3887 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3888 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3889 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3890 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3891 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3892 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3893 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3894 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3895 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R484 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R485 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R486 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R487 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3896 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3897 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3898 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3899 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3900 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3901 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3902 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X3903 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3904 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3905 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3906 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3907 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3908 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3909 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3910 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_14_20144# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3911 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3912 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3913 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3914 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3915 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3916 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3917 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3918 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3919 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3920 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3921 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3922 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3923 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3924 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3925 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3926 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3927 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R488 10good_0/9good_0/8good_1/7good_1/6good_1/m1_14_20144# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R489 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R490 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R491 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3928 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3929 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3930 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3931 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3932 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3933 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3934 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3935 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3936 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3937 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3938 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3939 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3940 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3941 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3942 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3943 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3944 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3945 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3946 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3947 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3948 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3949 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3950 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3951 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R492 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R493 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R494 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R495 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3952 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3953 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3954 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3955 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3956 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3957 vdda1 io_in[3] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3958 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X3959 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3960 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3961 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X3962 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3963 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3964 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3965 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3966 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X3967 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3968 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3969 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3970 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3971 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3972 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3973 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3974 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3975 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3976 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3977 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X3978 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3979 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3980 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3981 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3982 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3983 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3984 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3985 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X3986 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3987 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3988 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3989 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3990 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X3991 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R496 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R497 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R498 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R499 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X3992 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3993 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X3994 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3995 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X3996 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3997 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X3998 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X3999 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4000 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4001 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4002 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4003 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4004 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4005 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4006 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4007 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4008 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4009 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4010 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4011 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4012 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4013 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4014 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4015 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R500 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R501 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R502 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_31884_48# sky130_fd_pr__res_generic_po w=66 l=342
R503 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4016 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4017 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4018 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4019 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4020 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4021 vdda1 io_in[2] 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4022 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4023 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4024 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4025 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4026 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4027 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4028 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4029 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4030 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4031 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4032 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4033 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4034 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4035 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4036 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4037 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4038 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4039 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4040 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4041 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4042 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4043 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4044 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4045 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4046 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4047 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R504 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R505 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R506 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R507 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4048 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4049 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4050 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4051 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4052 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4053 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4054 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4055 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4056 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4057 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4058 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4059 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4060 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4061 vdda1 10good_0/9good_0/m1_32342_44672# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4062 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4063 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4064 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4065 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4066 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4067 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4068 vdda1 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4069 vdda1 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4070 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4071 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R508 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R509 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R510 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R511 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4072 10good_0/9good_0/8good_1/Sw-1_0/li_29_719# io_in[7] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4073 10good_0/9good_0/8good_1/m1_8774_43264# 10good_0/9good_0/8good_1/Sw-1_0/li_29_719# 10good_0/9good_0/m1_38716_44140# 10good_0/9good_0/8good_1/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X4074 10good_0/9good_0/m1_38716_44140# 10good_0/9good_0/8good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/m1_18694_42308# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4075 10good_0/9good_0/8good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4076 vdda1 10good_0/9good_0/8good_1/Sw-1_0/li_29_719# 10good_0/9good_0/8good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4077 vdda1 io_in[7] 10good_0/9good_0/8good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4078 10good_0/9good_0/m1_38716_44140# 10good_0/9good_0/8good_1/Sw-1_0/li_126_470# 10good_0/9good_0/8good_1/m1_18694_42308# 10good_0/9good_0/m1_38716_44140# sky130_fd_pr__pfet_01v8 w=84 l=30
X4079 10good_0/9good_0/8good_1/m1_8774_43264# 10good_0/9good_0/8good_1/Sw-1_0/li_126_470# 10good_0/9good_0/m1_38716_44140# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4080 10good_0/9good_0/Sw-1_0/li_29_719# io_in[8] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4081 10good_0/9good_0/m1_19068_42976# 10good_0/9good_0/Sw-1_0/li_29_719# 10good_0/m1_39076_44800# 10good_0/9good_0/m1_19068_42976# sky130_fd_pr__pfet_01v8 w=84 l=30
X4082 10good_0/m1_39076_44800# 10good_0/9good_0/Sw-1_0/li_29_719# 10good_0/9good_0/m1_38716_44140# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4083 10good_0/9good_0/Sw-1_0/li_126_470# 10good_0/9good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4084 vdda1 10good_0/9good_0/Sw-1_0/li_29_719# 10good_0/9good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4085 vdda1 io_in[8] 10good_0/9good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4086 10good_0/m1_39076_44800# 10good_0/9good_0/Sw-1_0/li_126_470# 10good_0/9good_0/m1_38716_44140# 10good_0/m1_39076_44800# sky130_fd_pr__pfet_01v8 w=84 l=30
X4087 10good_0/9good_0/m1_19068_42976# 10good_0/9good_0/Sw-1_0/li_126_470# 10good_0/m1_39076_44800# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4088 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4089 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X4090 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4091 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4092 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4093 vdda1 io_in[5] 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4094 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X4095 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4096 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4097 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4098 10good_0/9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4099 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4100 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4101 vdda1 io_in[4] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4102 10good_0/9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X4103 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4104 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4105 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4106 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4107 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4108 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4109 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4110 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X4111 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4112 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4113 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4114 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4115 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4116 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4117 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4118 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4119 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4120 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4121 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4122 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4123 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4124 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4125 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4126 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4127 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4128 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4129 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4130 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4131 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4132 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4133 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4134 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4135 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4136 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4137 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4138 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4139 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4140 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4141 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4142 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4143 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R512 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R513 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R514 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R515 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4144 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4145 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4146 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4147 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4148 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4149 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4150 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4151 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4152 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4153 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4154 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4155 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4156 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4157 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4158 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4159 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4160 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4161 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4162 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4163 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4164 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4165 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4166 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4167 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R516 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R517 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R518 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R519 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4168 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4169 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4170 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4171 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4172 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4173 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4174 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4175 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4176 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4177 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4178 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_41532_78# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4179 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4180 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4181 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4182 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_41532_78# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4183 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4184 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4185 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4186 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4187 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4188 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4189 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4190 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4191 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4192 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4193 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4194 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4195 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4196 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4197 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4198 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4199 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R520 10good_0/m1_41532_78# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R521 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R522 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R523 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4200 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4201 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4202 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4203 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4204 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4205 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4206 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4207 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4208 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4209 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4210 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4211 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4212 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4213 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4214 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4215 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4216 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4217 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4218 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4219 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4220 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4221 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4222 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4223 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R524 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R525 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R526 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R527 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4224 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4225 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4226 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4227 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4228 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4229 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4230 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4231 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4232 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4233 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4234 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4235 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4236 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4237 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4238 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4239 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4240 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4241 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4242 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4243 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4244 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4245 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4246 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4247 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4248 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4249 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4250 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4251 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4252 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4253 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4254 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4255 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4256 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4257 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4258 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4259 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4260 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4261 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4262 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4263 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R528 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R529 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R530 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R531 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4264 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4265 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4266 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4267 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4268 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4269 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4270 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4271 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4272 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4273 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4274 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4275 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4276 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4277 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4278 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4279 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4280 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4281 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4282 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4283 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4284 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4285 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4286 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4287 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R532 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R533 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R534 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R535 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4288 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4289 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4290 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4291 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4292 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4293 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4294 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4295 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4296 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4297 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4298 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4299 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4300 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4301 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4302 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4303 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4304 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4305 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4306 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4307 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4308 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4309 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4310 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4311 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4312 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4313 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4314 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4315 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4316 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4317 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4318 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4319 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R536 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R537 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R538 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R539 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4320 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4321 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4322 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4323 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4324 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4325 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4326 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4327 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4328 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4329 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4330 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4331 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4332 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4333 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4334 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4335 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4336 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4337 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4338 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4339 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4340 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4341 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4342 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4343 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R540 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R541 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R542 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R543 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4344 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4345 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4346 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4347 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4348 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4349 vdda1 io_in[4] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4350 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X4351 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4352 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4353 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4354 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4355 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4356 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4357 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4358 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X4359 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4360 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4361 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4362 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4363 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4364 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4365 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4366 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4367 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4368 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4369 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4370 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4371 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4372 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4373 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4374 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4375 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4376 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4377 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4378 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4379 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4380 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4381 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4382 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4383 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4384 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4385 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4386 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4387 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4388 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4389 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4390 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4391 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R544 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R545 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R546 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R547 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4392 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4393 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4394 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4395 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4396 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4397 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4398 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4399 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4400 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4401 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4402 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4403 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4404 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4405 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4406 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4407 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4408 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4409 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4410 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4411 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4412 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4413 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4414 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4415 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R548 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R549 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R550 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R551 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4416 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4417 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4418 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4419 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4420 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4421 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4422 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4423 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4424 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4425 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4426 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4427 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4428 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4429 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4430 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_14_20144# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4431 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4432 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4433 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4434 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4435 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4436 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4437 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4438 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4439 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4440 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4441 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4442 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4443 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4444 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4445 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4446 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4447 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R552 10good_0/9good_1/8good_0/7good_0/6good_0/m1_14_20144# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R553 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R554 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R555 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4448 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4449 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4450 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4451 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4452 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4453 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4454 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4455 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4456 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4457 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4458 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4459 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4460 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4461 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4462 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4463 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4464 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4465 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4466 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4467 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4468 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4469 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4470 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4471 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R556 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R557 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R558 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R559 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4472 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4473 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4474 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4475 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4476 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4477 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4478 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4479 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4480 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4481 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4482 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4483 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4484 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4485 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4486 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4487 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4488 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4489 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4490 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4491 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4492 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4493 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4494 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4495 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4496 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4497 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4498 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4499 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4500 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4501 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4502 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4503 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4504 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4505 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4506 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4507 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4508 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4509 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4510 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4511 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R560 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R561 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R562 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R563 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4512 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4513 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4514 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4515 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4516 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4517 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4518 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4519 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4520 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4521 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4522 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4523 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4524 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4525 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4526 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4527 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4528 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4529 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4530 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4531 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4532 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4533 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4534 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4535 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R564 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R565 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R566 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_36912_2# sky130_fd_pr__res_generic_po w=66 l=342
R567 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4536 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4537 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4538 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4539 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4540 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4541 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4542 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4543 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4544 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4545 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4546 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4547 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4548 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4549 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4550 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4551 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4552 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4553 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4554 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4555 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4556 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4557 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4558 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4559 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4560 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4561 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4562 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4563 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4564 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4565 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4566 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4567 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R568 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R569 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R570 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R571 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4568 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4569 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4570 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4571 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4572 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4573 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4574 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4575 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4576 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4577 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4578 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4579 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4580 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4581 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4582 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4583 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4584 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4585 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4586 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4587 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4588 vdda1 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4589 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4590 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4591 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R572 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R573 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R574 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R575 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4592 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_29_719# io_in[6] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4593 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/m1_8774_43264# 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X4594 10good_0/9good_1/8good_0/m1_8774_43264# 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4595 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4596 vdda1 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4597 vdda1 io_in[6] 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4598 10good_0/9good_1/8good_0/m1_8774_43264# 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/m1_8436_40544# 10good_0/9good_1/8good_0/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X4599 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# 10good_0/9good_1/8good_0/7good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/m1_8774_43264# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4600 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4601 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/m1_8436_40544# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X4602 10good_0/9good_1/8good_0/7good_0/m1_8436_40544# 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4603 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4604 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4605 vdda1 io_in[5] 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4606 10good_0/9good_1/8good_0/7good_0/m1_8436_40544# 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X4607 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4608 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4609 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4610 10good_0/9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4611 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4612 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4613 vdda1 io_in[4] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4614 10good_0/9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X4615 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4616 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4617 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4618 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4619 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4620 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4621 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4622 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X4623 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4624 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4625 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4626 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4627 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4628 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4629 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4630 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4631 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4632 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4633 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4634 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4635 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4636 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4637 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4638 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4639 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4640 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4641 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4642 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4643 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4644 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4645 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4646 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4647 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4648 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4649 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4650 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4651 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4652 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4653 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4654 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4655 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R576 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R577 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R578 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R579 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4656 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4657 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4658 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4659 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4660 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4661 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4662 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4663 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4664 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4665 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4666 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4667 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4668 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4669 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4670 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4671 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4672 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4673 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4674 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4675 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4676 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4677 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4678 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4679 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R580 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R581 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R582 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R583 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4680 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4681 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4682 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4683 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4684 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4685 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4686 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4687 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4688 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4689 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4690 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_46616_8# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4691 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4692 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4693 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4694 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_46616_8# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4695 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4696 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4697 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4698 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4699 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4700 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4701 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4702 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4703 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4704 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4705 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4706 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4707 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4708 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4709 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4710 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4711 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R584 10good_0/m1_46616_8# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R585 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R586 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R587 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4712 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4713 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4714 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4715 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4716 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4717 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4718 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4719 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4720 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4721 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4722 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4723 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4724 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4725 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4726 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4727 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4728 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4729 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4730 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4731 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4732 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4733 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4734 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4735 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R588 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R589 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R590 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R591 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4736 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4737 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4738 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4739 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4740 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4741 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4742 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4743 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4744 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4745 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4746 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4747 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4748 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4749 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4750 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4751 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4752 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4753 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4754 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4755 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4756 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4757 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4758 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4759 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4760 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4761 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4762 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4763 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4764 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4765 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4766 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4767 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4768 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4769 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4770 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4771 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4772 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4773 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4774 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4775 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R592 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R593 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R594 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R595 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4776 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4777 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4778 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4779 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4780 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4781 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4782 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4783 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4784 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4785 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4786 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4787 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4788 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4789 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4790 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4791 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4792 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4793 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4794 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4795 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4796 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4797 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4798 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4799 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R596 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R597 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R598 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R599 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4800 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4801 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4802 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4803 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4804 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4805 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4806 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4807 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4808 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4809 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4810 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4811 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4812 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4813 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4814 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4815 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4816 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4817 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4818 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4819 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4820 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4821 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4822 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4823 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4824 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4825 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4826 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4827 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4828 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4829 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4830 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4831 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R600 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R601 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R602 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R603 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4832 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4833 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4834 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4835 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4836 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4837 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4838 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4839 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4840 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4841 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4842 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4843 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4844 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4845 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4846 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4847 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4848 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4849 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4850 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4851 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4852 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4853 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4854 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4855 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R604 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R605 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R606 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R607 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4856 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4857 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4858 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4859 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4860 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4861 vdda1 io_in[4] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4862 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X4863 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4864 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4865 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4866 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4867 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4868 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4869 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4870 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X4871 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4872 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4873 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4874 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4875 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4876 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4877 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4878 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4879 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4880 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4881 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4882 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4883 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4884 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4885 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4886 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4887 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4888 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4889 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4890 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4891 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4892 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4893 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4894 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4895 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4896 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4897 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4898 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4899 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4900 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4901 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4902 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4903 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R608 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R609 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R610 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R611 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4904 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4905 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4906 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4907 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4908 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4909 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4910 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4911 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4912 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4913 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4914 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4915 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4916 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4917 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4918 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4919 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4920 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4921 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4922 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4923 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4924 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4925 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4926 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4927 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R612 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R613 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R614 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R615 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4928 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4929 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4930 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4931 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4932 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4933 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4934 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X4935 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4936 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4937 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4938 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4939 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4940 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4941 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4942 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/m1_14_20144# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4943 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4944 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4945 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4946 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4947 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4948 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4949 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4950 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4951 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4952 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4953 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4954 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4955 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4956 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4957 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4958 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X4959 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R616 10good_0/9good_1/8good_0/7good_0/6good_1/m1_14_20144# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R617 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R618 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R619 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4960 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4961 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X4962 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4963 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4964 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4965 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4966 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X4967 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4968 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4969 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X4970 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4971 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4972 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4973 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4974 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4975 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4976 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4977 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X4978 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4979 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4980 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4981 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4982 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4983 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R620 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R621 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R622 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R623 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X4984 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4985 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4986 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4987 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4988 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4989 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4990 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X4991 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4992 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4993 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X4994 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4995 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X4996 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4997 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X4998 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X4999 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5000 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5001 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5002 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5003 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5004 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5005 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5006 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5007 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5008 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5009 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5010 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5011 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5012 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5013 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5014 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5015 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5016 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5017 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5018 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5019 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5020 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5021 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5022 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5023 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R624 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R625 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R626 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R627 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5024 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5025 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5026 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5027 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5028 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5029 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5030 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5031 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5032 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5033 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5034 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5035 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5036 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5037 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5038 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5039 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5040 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5041 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5042 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5043 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5044 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5045 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5046 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5047 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R628 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R629 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R630 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_41532_78# sky130_fd_pr__res_generic_po w=66 l=342
R631 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5048 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5049 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5050 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5051 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5052 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5053 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5054 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5055 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5056 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5057 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5058 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5059 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5060 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5061 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5062 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5063 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5064 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5065 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5066 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5067 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5068 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5069 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5070 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5071 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5072 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5073 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5074 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5075 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5076 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5077 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5078 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5079 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R632 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R633 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R634 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R635 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5080 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5081 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5082 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5083 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5084 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5085 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5086 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5087 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5088 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5089 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5090 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5091 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5092 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5093 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5094 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5095 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5096 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5097 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5098 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5099 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5100 vdda1 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5101 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5102 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5103 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R636 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R637 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R638 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R639 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5104 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5105 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X5106 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5107 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5108 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5109 vdda1 io_in[5] 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5110 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X5111 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5112 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5113 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5114 10good_0/9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5115 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5116 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5117 vdda1 io_in[4] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5118 10good_0/9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X5119 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5120 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5121 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5122 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5123 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5124 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5125 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5126 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X5127 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5128 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5129 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5130 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5131 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5132 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5133 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5134 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5135 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5136 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5137 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5138 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5139 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5140 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5141 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5142 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5143 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5144 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5145 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5146 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5147 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5148 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5149 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5150 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5151 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5152 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5153 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5154 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5155 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5156 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5157 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5158 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5159 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R640 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R641 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R642 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R643 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5160 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5161 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5162 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5163 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5164 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5165 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5166 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5167 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5168 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5169 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5170 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5171 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5172 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5173 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5174 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5175 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5176 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5177 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5178 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5179 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5180 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5181 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5182 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5183 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R644 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R645 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R646 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R647 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5184 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5185 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5186 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5187 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5188 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5189 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5190 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5191 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5192 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5193 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5194 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_51780_62# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5195 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5196 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5197 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5198 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_51780_62# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5199 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5200 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5201 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5202 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5203 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5204 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5205 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5206 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5207 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5208 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5209 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5210 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5211 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5212 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5213 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5214 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5215 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R648 10good_0/m1_51780_62# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R649 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R650 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R651 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5216 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5217 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5218 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5219 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5220 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5221 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5222 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5223 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5224 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5225 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5226 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5227 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5228 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5229 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5230 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5231 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5232 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5233 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5234 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5235 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5236 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5237 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5238 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5239 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R652 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R653 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R654 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R655 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5240 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5241 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5242 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5243 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5244 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5245 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5246 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5247 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5248 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5249 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5250 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5251 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5252 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5253 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5254 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5255 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5256 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5257 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5258 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5259 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5260 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5261 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5262 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5263 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5264 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5265 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5266 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5267 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5268 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5269 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5270 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5271 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5272 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5273 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5274 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5275 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5276 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5277 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5278 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5279 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R656 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R657 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R658 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R659 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5280 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5281 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5282 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5283 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5284 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5285 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5286 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5287 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5288 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5289 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5290 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5291 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5292 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5293 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5294 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5295 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5296 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5297 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5298 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5299 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5300 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5301 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5302 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5303 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R660 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R661 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R662 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R663 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5304 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5305 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5306 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5307 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5308 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5309 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5310 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5311 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5312 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5313 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5314 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5315 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5316 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5317 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5318 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5319 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5320 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5321 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5322 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5323 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5324 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5325 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5326 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5327 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5328 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5329 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5330 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5331 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5332 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5333 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5334 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5335 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R664 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R665 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R666 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R667 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5336 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5337 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5338 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5339 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5340 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5341 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5342 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5343 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5344 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5345 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5346 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5347 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5348 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5349 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5350 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5351 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5352 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5353 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5354 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5355 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5356 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5357 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5358 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5359 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R668 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R669 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R670 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R671 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5360 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5361 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5362 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5363 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5364 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5365 vdda1 io_in[4] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5366 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X5367 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5368 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5369 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5370 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5371 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5372 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5373 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5374 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X5375 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5376 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5377 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5378 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5379 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5380 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5381 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5382 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5383 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5384 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5385 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5386 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5387 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5388 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5389 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5390 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5391 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5392 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5393 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5394 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5395 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5396 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5397 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5398 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5399 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5400 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5401 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5402 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5403 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5404 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5405 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5406 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5407 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R672 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R673 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R674 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R675 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5408 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5409 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5410 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5411 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5412 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5413 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5414 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5415 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5416 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5417 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5418 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5419 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5420 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5421 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5422 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5423 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5424 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5425 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5426 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5427 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5428 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5429 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5430 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5431 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R676 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R677 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R678 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R679 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5432 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5433 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5434 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5435 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5436 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5437 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5438 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5439 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5440 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5441 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5442 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5443 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5444 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5445 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5446 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/m1_14_20144# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5447 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5448 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5449 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5450 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5451 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5452 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5453 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5454 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5455 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5456 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5457 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5458 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5459 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5460 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5461 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5462 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5463 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R680 10good_0/9good_1/8good_0/7good_1/6good_0/m1_14_20144# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R681 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R682 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R683 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5464 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5465 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5466 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5467 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5468 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5469 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5470 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5471 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5472 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5473 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5474 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5475 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5476 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5477 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5478 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5479 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5480 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5481 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5482 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5483 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5484 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5485 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5486 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5487 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R684 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R685 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R686 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R687 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5488 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5489 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5490 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5491 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5492 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5493 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5494 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5495 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5496 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5497 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5498 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5499 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5500 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5501 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5502 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5503 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5504 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5505 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5506 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5507 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5508 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5509 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5510 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5511 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5512 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5513 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5514 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5515 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5516 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5517 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5518 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5519 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5520 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5521 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5522 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5523 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5524 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5525 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5526 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5527 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R688 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R689 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R690 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R691 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5528 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5529 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5530 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5531 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5532 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5533 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5534 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5535 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5536 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5537 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5538 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5539 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5540 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5541 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5542 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5543 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5544 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5545 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5546 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5547 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5548 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5549 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5550 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5551 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R692 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R693 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R694 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_46616_8# sky130_fd_pr__res_generic_po w=66 l=342
R695 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5552 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5553 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5554 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5555 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5556 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5557 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5558 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5559 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5560 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5561 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5562 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5563 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5564 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5565 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5566 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5567 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5568 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5569 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5570 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5571 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5572 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5573 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5574 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5575 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5576 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5577 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5578 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5579 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5580 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5581 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5582 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5583 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R696 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R697 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R698 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R699 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5584 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5585 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5586 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5587 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5588 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5589 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5590 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5591 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5592 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5593 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5594 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5595 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5596 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5597 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5598 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5599 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5600 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5601 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5602 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5603 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5604 vdda1 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5605 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5606 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5607 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R700 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R701 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R702 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R703 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5608 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_29_719# io_in[6] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5609 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/m1_18694_42308# 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X5610 10good_0/9good_1/8good_0/m1_18694_42308# 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5611 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5612 vdda1 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5613 vdda1 io_in[6] 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5614 10good_0/9good_1/8good_0/m1_18694_42308# 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# 10good_0/9good_1/8good_0/m1_18694_42308# sky130_fd_pr__pfet_01v8 w=84 l=30
X5615 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# 10good_0/9good_1/8good_0/7good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/m1_18694_42308# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5616 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5617 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X5618 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5619 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5620 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5621 vdda1 io_in[5] 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5622 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X5623 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5624 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5625 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5626 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5627 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5628 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5629 vdda1 io_in[4] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5630 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X5631 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5632 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5633 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5634 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5635 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5636 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5637 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5638 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X5639 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5640 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5641 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5642 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5643 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5644 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5645 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5646 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5647 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5648 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5649 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5650 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5651 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5652 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5653 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5654 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5655 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5656 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5657 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5658 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5659 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5660 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5661 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5662 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5663 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5664 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5665 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5666 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5667 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5668 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5669 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5670 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5671 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R704 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R705 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R706 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R707 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5672 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5673 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5674 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5675 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5676 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5677 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5678 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5679 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5680 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5681 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5682 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5683 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5684 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5685 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5686 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5687 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5688 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5689 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5690 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5691 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5692 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5693 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5694 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5695 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R708 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R709 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R710 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R711 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5696 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5697 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5698 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5699 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5700 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5701 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5702 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5703 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5704 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5705 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5706 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_56844_12# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5707 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5708 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5709 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5710 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_56844_12# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5711 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5712 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5713 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5714 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5715 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5716 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5717 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5718 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5719 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5720 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5721 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5722 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5723 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5724 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5725 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5726 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5727 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R712 10good_0/m1_56844_12# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R713 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R714 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R715 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5728 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5729 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5730 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5731 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5732 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5733 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5734 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5735 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5736 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5737 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5738 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5739 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5740 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5741 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5742 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5743 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5744 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5745 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5746 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5747 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5748 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5749 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5750 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5751 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R716 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R717 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R718 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R719 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5752 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5753 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5754 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5755 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5756 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5757 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5758 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5759 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5760 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5761 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5762 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5763 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5764 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5765 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5766 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5767 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5768 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5769 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5770 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5771 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5772 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5773 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5774 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5775 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5776 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5777 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5778 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5779 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5780 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5781 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5782 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5783 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5784 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5785 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5786 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5787 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5788 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5789 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5790 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5791 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R720 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R721 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R722 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R723 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5792 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5793 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5794 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5795 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5796 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5797 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5798 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5799 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5800 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5801 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5802 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5803 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5804 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5805 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5806 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5807 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5808 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5809 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5810 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5811 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5812 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5813 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5814 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5815 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R724 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R725 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R726 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R727 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5816 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5817 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5818 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5819 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5820 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5821 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5822 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5823 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5824 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5825 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5826 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5827 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5828 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5829 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5830 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5831 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5832 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5833 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5834 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5835 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5836 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5837 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5838 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5839 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5840 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5841 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5842 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5843 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5844 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5845 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5846 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5847 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R728 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R729 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R730 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R731 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5848 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5849 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5850 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5851 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5852 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5853 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5854 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5855 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5856 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5857 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5858 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5859 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5860 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5861 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5862 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5863 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5864 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5865 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5866 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5867 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5868 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5869 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5870 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5871 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R732 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R733 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R734 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R735 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5872 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5873 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X5874 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5875 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5876 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5877 vdda1 io_in[4] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5878 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X5879 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5880 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5881 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5882 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5883 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5884 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5885 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5886 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X5887 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5888 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5889 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5890 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5891 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5892 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5893 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5894 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X5895 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5896 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5897 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5898 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5899 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5900 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5901 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5902 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5903 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5904 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5905 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5906 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5907 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5908 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5909 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5910 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5911 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5912 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5913 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5914 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5915 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5916 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5917 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5918 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5919 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R736 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R737 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R738 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R739 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5920 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5921 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5922 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5923 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5924 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5925 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5926 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5927 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5928 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5929 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5930 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5931 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5932 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5933 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5934 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5935 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5936 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5937 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5938 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5939 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5940 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5941 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5942 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5943 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R740 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R741 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R742 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R743 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5944 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5945 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5946 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5947 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5948 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5949 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5950 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X5951 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5952 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5953 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5954 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5955 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5956 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5957 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5958 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_14_20144# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5959 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5960 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5961 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5962 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5963 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5964 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5965 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5966 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5967 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5968 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5969 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5970 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5971 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5972 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5973 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5974 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X5975 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R744 10good_0/9good_1/8good_0/7good_1/6good_1/m1_14_20144# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R745 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R746 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R747 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X5976 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5977 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X5978 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5979 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5980 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5981 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5982 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X5983 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5984 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5985 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X5986 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5987 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5988 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5989 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5990 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5991 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5992 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5993 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X5994 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5995 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X5996 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5997 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X5998 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X5999 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R748 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R749 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R750 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R751 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6000 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6001 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6002 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6003 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6004 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6005 vdda1 io_in[3] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6006 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6007 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6008 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6009 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6010 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6011 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6012 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6013 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6014 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6015 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6016 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6017 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6018 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6019 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6020 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6021 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6022 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6023 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6024 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6025 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6026 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6027 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6028 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6029 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6030 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6031 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6032 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6033 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6034 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6035 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6036 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6037 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6038 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6039 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R752 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R753 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R754 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R755 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6040 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6041 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6042 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6043 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6044 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6045 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6046 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6047 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6048 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6049 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6050 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6051 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6052 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6053 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6054 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6055 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6056 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6057 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6058 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6059 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6060 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6061 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6062 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6063 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R756 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R757 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R758 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_51780_62# sky130_fd_pr__res_generic_po w=66 l=342
R759 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6064 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6065 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6066 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6067 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6068 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6069 vdda1 io_in[2] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6070 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6071 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6072 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6073 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6074 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6075 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6076 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6077 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6078 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6079 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6080 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6081 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6082 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6083 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6084 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6085 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6086 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6087 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6088 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6089 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6090 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6091 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6092 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6093 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6094 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6095 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R760 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R761 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R762 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R763 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6096 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6097 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6098 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6099 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6100 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6101 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6102 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6103 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6104 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# io_in[0] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6105 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6106 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6107 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6108 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6109 vdda1 io_in[0] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6110 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6111 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6112 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# io_in[1] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6113 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6114 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6115 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6116 vdda1 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6117 vdda1 io_in[1] 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6118 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6119 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R764 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R765 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R766 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R767 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6120 10good_0/9good_1/8good_0/Sw-1_0/li_29_719# io_in[7] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6121 10good_0/9good_1/8good_0/m1_8774_43264# 10good_0/9good_1/8good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_19068_42976# 10good_0/9good_1/8good_0/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X6122 10good_0/9good_1/m1_19068_42976# 10good_0/9good_1/8good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/m1_18694_42308# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6123 10good_0/9good_1/8good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6124 vdda1 10good_0/9good_1/8good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6125 vdda1 io_in[7] 10good_0/9good_1/8good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6126 10good_0/9good_1/m1_19068_42976# 10good_0/9good_1/8good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_0/m1_18694_42308# 10good_0/9good_1/m1_19068_42976# sky130_fd_pr__pfet_01v8 w=84 l=30
X6127 10good_0/9good_1/8good_0/m1_8774_43264# 10good_0/9good_1/8good_0/Sw-1_0/li_126_470# 10good_0/9good_1/m1_19068_42976# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6128 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6129 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X6130 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6131 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6132 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6133 vdda1 io_in[5] 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6134 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X6135 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6136 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6137 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6138 10good_0/9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6139 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6140 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6141 vdda1 io_in[4] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6142 10good_0/9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X6143 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6144 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6145 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6146 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6147 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6148 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6149 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6150 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X6151 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6152 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6153 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6154 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6155 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6156 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6157 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6158 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6159 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6160 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6161 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6162 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6163 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6164 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6165 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6166 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6167 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6168 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6169 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6170 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6171 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6172 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6173 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6174 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6175 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6176 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6177 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6178 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6179 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6180 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6181 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6182 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6183 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R768 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R769 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R770 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R771 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6184 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6185 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6186 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6187 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6188 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6189 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6190 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6191 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6192 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6193 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6194 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6195 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6196 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6197 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6198 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6199 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6200 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6201 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6202 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6203 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6204 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6205 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6206 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6207 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R772 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R773 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R774 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R775 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6208 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6209 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6210 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6211 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6212 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6213 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6214 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6215 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6216 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6217 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6218 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_61528_92# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6219 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6220 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6221 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6222 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_61528_92# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6223 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6224 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6225 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6226 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6227 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6228 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6229 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6230 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6231 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6232 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6233 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6234 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6235 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6236 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6237 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6238 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6239 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R776 10good_0/m1_61528_92# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R777 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R778 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R779 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6240 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6241 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6242 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6243 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6244 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6245 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6246 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6247 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6248 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6249 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6250 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6251 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6252 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6253 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6254 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6255 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6256 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6257 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6258 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6259 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6260 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6261 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6262 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6263 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R780 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R781 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R782 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R783 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6264 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6265 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6266 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6267 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6268 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6269 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6270 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6271 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6272 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6273 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6274 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6275 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6276 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6277 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6278 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6279 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6280 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6281 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6282 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6283 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6284 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6285 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6286 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6287 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6288 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6289 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6290 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6291 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6292 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6293 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6294 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6295 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6296 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6297 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6298 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6299 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6300 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6301 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6302 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6303 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R784 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R785 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R786 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R787 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6304 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6305 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6306 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6307 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6308 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6309 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6310 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6311 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6312 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6313 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6314 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6315 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6316 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6317 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6318 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6319 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6320 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6321 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6322 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6323 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6324 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6325 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6326 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6327 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R788 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R789 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R790 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R791 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6328 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6329 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6330 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6331 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6332 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6333 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6334 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6335 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6336 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6337 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6338 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6339 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6340 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6341 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6342 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6343 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6344 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6345 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6346 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6347 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6348 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6349 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6350 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6351 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6352 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6353 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6354 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6355 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6356 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6357 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6358 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6359 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R792 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R793 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R794 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R795 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6360 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6361 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6362 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6363 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6364 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6365 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6366 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6367 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6368 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6369 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6370 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6371 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6372 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6373 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6374 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6375 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6376 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6377 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6378 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6379 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6380 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6381 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6382 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6383 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R796 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R797 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R798 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R799 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6384 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6385 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6386 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6387 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6388 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6389 vdda1 io_in[4] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6390 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X6391 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6392 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6393 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6394 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6395 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6396 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6397 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6398 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X6399 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6400 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6401 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6402 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6403 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6404 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6405 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6406 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6407 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6408 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6409 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6410 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6411 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6412 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6413 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6414 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6415 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6416 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6417 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6418 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6419 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6420 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6421 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6422 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6423 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6424 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6425 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6426 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6427 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6428 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6429 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6430 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6431 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R800 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R801 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R802 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R803 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6432 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6433 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6434 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6435 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6436 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6437 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6438 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6439 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6440 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6441 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6442 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6443 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6444 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6445 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6446 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6447 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6448 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6449 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6450 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6451 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6452 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6453 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6454 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6455 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R804 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R805 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R806 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R807 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6456 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6457 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6458 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6459 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6460 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6461 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6462 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6463 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6464 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6465 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6466 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6467 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6468 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6469 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6470 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_14_20144# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6471 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6472 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6473 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6474 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6475 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6476 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6477 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6478 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6479 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6480 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6481 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6482 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6483 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6484 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6485 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6486 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6487 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R808 10good_0/9good_1/8good_1/7good_0/6good_0/m1_14_20144# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R809 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R810 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R811 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6488 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6489 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6490 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6491 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6492 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6493 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6494 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6495 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6496 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6497 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6498 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6499 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6500 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6501 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6502 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6503 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6504 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6505 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6506 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6507 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6508 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6509 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6510 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6511 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R812 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R813 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R814 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R815 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6512 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6513 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6514 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6515 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6516 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6517 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6518 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6519 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6520 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6521 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6522 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6523 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6524 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6525 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6526 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6527 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6528 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6529 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6530 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6531 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6532 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6533 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6534 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6535 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6536 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6537 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6538 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6539 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6540 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6541 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6542 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6543 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6544 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6545 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6546 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6547 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6548 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6549 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6550 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6551 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R816 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R817 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R818 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R819 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6552 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6553 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6554 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6555 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6556 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6557 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6558 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6559 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6560 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6561 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6562 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6563 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6564 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6565 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6566 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6567 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6568 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6569 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6570 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6571 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6572 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6573 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6574 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6575 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R820 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R821 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R822 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_56844_12# sky130_fd_pr__res_generic_po w=66 l=342
R823 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6576 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6577 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6578 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6579 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6580 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6581 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6582 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6583 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6584 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6585 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6586 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6587 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6588 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6589 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6590 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6591 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6592 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6593 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6594 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6595 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6596 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6597 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6598 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6599 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6600 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6601 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6602 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6603 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6604 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6605 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6606 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6607 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R824 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R825 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R826 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R827 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6608 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6609 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6610 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6611 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6612 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6613 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6614 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6615 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6616 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6617 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6618 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6619 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6620 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6621 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6622 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6623 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6624 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6625 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6626 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6627 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6628 vdda1 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6629 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6630 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6631 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R828 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R829 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R830 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R831 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6632 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_29_719# io_in[6] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6633 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/m1_8774_43264# 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X6634 10good_0/9good_1/8good_1/m1_8774_43264# 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6635 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6636 vdda1 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6637 vdda1 io_in[6] 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6638 10good_0/9good_1/8good_1/m1_8774_43264# 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/m1_8436_40544# 10good_0/9good_1/8good_1/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X6639 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# 10good_0/9good_1/8good_1/7good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/m1_8774_43264# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6640 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6641 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/m1_8436_40544# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X6642 10good_0/9good_1/8good_1/7good_0/m1_8436_40544# 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6643 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6644 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6645 vdda1 io_in[5] 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6646 10good_0/9good_1/8good_1/7good_0/m1_8436_40544# 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X6647 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6648 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6649 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6650 10good_0/9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6651 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6652 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6653 vdda1 io_in[4] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6654 10good_0/9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X6655 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6656 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6657 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6658 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6659 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6660 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6661 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6662 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X6663 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6664 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6665 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6666 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6667 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6668 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6669 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6670 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6671 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6672 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6673 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6674 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6675 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6676 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6677 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6678 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6679 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6680 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6681 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6682 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6683 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6684 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6685 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6686 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6687 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6688 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6689 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6690 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6691 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6692 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6693 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6694 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6695 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R832 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R833 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R834 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R835 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6696 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6697 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6698 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6699 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6700 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6701 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6702 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6703 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6704 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6705 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6706 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6707 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6708 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6709 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6710 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6711 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6712 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6713 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6714 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6715 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6716 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6717 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6718 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6719 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R836 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R837 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R838 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R839 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6720 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6721 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6722 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6723 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6724 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6725 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6726 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6727 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6728 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6729 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6730 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_66618_22# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6731 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6732 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6733 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6734 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_66618_22# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6735 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6736 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6737 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6738 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6739 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6740 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6741 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6742 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6743 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6744 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6745 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6746 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6747 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6748 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6749 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6750 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6751 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R840 10good_0/m1_66618_22# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R841 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R842 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R843 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6752 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6753 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6754 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6755 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6756 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6757 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6758 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6759 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6760 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6761 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6762 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6763 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6764 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6765 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6766 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6767 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6768 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6769 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6770 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6771 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6772 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6773 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6774 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6775 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R844 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R845 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R846 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R847 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6776 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6777 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6778 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6779 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6780 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6781 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6782 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6783 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6784 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6785 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6786 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6787 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6788 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6789 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6790 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6791 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6792 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6793 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6794 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6795 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6796 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6797 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6798 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6799 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6800 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6801 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6802 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6803 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6804 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6805 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6806 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6807 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6808 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6809 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6810 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6811 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6812 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6813 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6814 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6815 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R848 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R849 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R850 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R851 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6816 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6817 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6818 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6819 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6820 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6821 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6822 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6823 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6824 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6825 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6826 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6827 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6828 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6829 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6830 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6831 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6832 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6833 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6834 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6835 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6836 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6837 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6838 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6839 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R852 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R853 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R854 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R855 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6840 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6841 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6842 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6843 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6844 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6845 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6846 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6847 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6848 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6849 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6850 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6851 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6852 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6853 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6854 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6855 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6856 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6857 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6858 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6859 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6860 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6861 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6862 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6863 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6864 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6865 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6866 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6867 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6868 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6869 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6870 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6871 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R856 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R857 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R858 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R859 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6872 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6873 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6874 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6875 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6876 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6877 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6878 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6879 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6880 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6881 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6882 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6883 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6884 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6885 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6886 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6887 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6888 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6889 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6890 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6891 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6892 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6893 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6894 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6895 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R860 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R861 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R862 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R863 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6896 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6897 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X6898 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6899 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6900 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6901 vdda1 io_in[4] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6902 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X6903 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6904 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6905 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6906 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6907 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6908 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6909 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6910 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X6911 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6912 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6913 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6914 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6915 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6916 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6917 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6918 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X6919 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6920 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6921 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6922 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6923 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6924 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6925 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6926 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6927 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6928 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6929 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6930 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6931 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6932 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6933 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6934 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6935 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6936 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6937 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6938 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6939 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6940 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6941 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6942 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6943 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R864 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R865 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R866 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R867 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6944 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6945 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6946 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6947 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6948 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6949 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6950 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6951 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6952 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6953 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6954 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6955 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6956 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6957 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6958 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6959 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6960 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6961 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6962 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6963 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6964 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6965 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6966 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6967 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R868 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R869 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R870 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R871 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X6968 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6969 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X6970 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6971 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6972 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6973 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6974 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X6975 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6976 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6977 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X6978 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6979 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6980 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6981 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6982 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/m1_14_20144# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X6983 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6984 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6985 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X6986 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6987 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6988 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6989 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6990 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6991 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6992 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6993 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X6994 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6995 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X6996 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6997 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X6998 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X6999 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R872 10good_0/9good_1/8good_1/7good_0/6good_1/m1_14_20144# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R873 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R874 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R875 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7000 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7001 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7002 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7003 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7004 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7005 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7006 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7007 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7008 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7009 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7010 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7011 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7012 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7013 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7014 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7015 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7016 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7017 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7018 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7019 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7020 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7021 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7022 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7023 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R876 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R877 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R878 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R879 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7024 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7025 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7026 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7027 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7028 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7029 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7030 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7031 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7032 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7033 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7034 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7035 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7036 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7037 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7038 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7039 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7040 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7041 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7042 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7043 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7044 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7045 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7046 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7047 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7048 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7049 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7050 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7051 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7052 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7053 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7054 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7055 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7056 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7057 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7058 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7059 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7060 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7061 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7062 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7063 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R880 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R881 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R882 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R883 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7064 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7065 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7066 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7067 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7068 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7069 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7070 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7071 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7072 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7073 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7074 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7075 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7076 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7077 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7078 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7079 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7080 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7081 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7082 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7083 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7084 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7085 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7086 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7087 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R884 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R885 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R886 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_61528_92# sky130_fd_pr__res_generic_po w=66 l=342
R887 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7088 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7089 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7090 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7091 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7092 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7093 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7094 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7095 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7096 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7097 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7098 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7099 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7100 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7101 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7102 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7103 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7104 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7105 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7106 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7107 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7108 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7109 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7110 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7111 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7112 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7113 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7114 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7115 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7116 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7117 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7118 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7119 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R888 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R889 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R890 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R891 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7120 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7121 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7122 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7123 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7124 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7125 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7126 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7127 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7128 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7129 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7130 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7131 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7132 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7133 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7134 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7135 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7136 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7137 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7138 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7139 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7140 vdda1 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7141 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7142 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7143 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R892 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R893 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R894 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R895 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7144 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7145 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X7146 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7147 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7148 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7149 vdda1 io_in[5] 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7150 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X7151 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7152 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7153 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7154 10good_0/9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7155 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7156 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7157 vdda1 io_in[4] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7158 10good_0/9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X7159 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7160 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7161 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7162 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7163 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7164 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7165 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7166 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X7167 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7168 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7169 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7170 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7171 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7172 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7173 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7174 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7175 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7176 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7177 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7178 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7179 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7180 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7181 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7182 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7183 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7184 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7185 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7186 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7187 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7188 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7189 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7190 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7191 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7192 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7193 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7194 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7195 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7196 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7197 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7198 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7199 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R896 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R897 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R898 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R899 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7200 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7201 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7202 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7203 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7204 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7205 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7206 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7207 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7208 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7209 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7210 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7211 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7212 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7213 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7214 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7215 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7216 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7217 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7218 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7219 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7220 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7221 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7222 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7223 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R900 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R901 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R902 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R903 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7224 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7225 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7226 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7227 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7228 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7229 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7230 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7231 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7232 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7233 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7234 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_71736_52# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7235 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7236 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7237 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7238 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_71736_52# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7239 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7240 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7241 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7242 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7243 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7244 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7245 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7246 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7247 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7248 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7249 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7250 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7251 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7252 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7253 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7254 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7255 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R904 10good_0/m1_71736_52# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R905 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R906 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R907 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7256 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7257 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7258 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7259 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7260 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7261 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7262 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7263 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7264 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7265 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7266 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7267 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7268 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7269 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7270 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7271 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7272 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7273 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7274 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7275 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7276 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7277 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7278 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7279 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R908 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R909 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R910 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R911 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7280 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7281 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7282 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7283 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7284 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7285 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7286 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7287 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7288 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7289 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7290 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7291 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7292 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7293 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7294 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7295 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7296 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7297 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7298 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7299 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7300 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7301 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7302 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7303 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7304 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7305 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7306 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7307 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7308 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7309 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7310 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7311 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7312 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7313 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7314 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7315 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7316 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7317 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7318 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7319 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R912 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R913 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R914 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R915 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7320 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7321 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7322 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7323 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7324 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7325 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7326 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7327 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7328 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7329 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7330 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7331 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7332 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7333 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7334 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7335 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7336 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7337 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7338 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7339 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7340 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7341 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7342 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7343 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R916 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R917 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R918 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R919 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7344 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7345 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7346 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7347 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7348 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7349 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7350 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7351 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7352 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7353 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7354 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7355 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7356 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7357 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7358 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7359 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7360 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7361 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7362 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7363 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7364 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7365 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7366 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7367 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7368 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7369 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7370 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7371 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7372 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7373 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7374 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7375 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R920 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R921 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R922 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R923 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7376 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7377 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7378 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7379 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7380 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7381 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7382 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7383 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7384 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7385 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7386 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7387 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7388 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7389 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7390 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7391 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7392 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7393 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7394 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7395 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7396 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7397 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7398 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7399 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R924 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R925 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R926 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R927 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7400 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7401 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7402 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7403 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7404 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7405 vdda1 io_in[4] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7406 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X7407 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7408 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7409 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7410 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7411 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7412 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7413 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7414 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X7415 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7416 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7417 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7418 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7419 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7420 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7421 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7422 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7423 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7424 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7425 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7426 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7427 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7428 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7429 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7430 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7431 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7432 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7433 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7434 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7435 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7436 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7437 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7438 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7439 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7440 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7441 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7442 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7443 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7444 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7445 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7446 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7447 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R928 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R929 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R930 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R931 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7448 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7449 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7450 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7451 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7452 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7453 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7454 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7455 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7456 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7457 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7458 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7459 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7460 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7461 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7462 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7463 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7464 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7465 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7466 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7467 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7468 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7469 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7470 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7471 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R932 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R933 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R934 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R935 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7472 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7473 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7474 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7475 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7476 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7477 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7478 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7479 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7480 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7481 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7482 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7483 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7484 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7485 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7486 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/m1_14_20144# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7487 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7488 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7489 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7490 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7491 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7492 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7493 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7494 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7495 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7496 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7497 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7498 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7499 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7500 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7501 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7502 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7503 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R936 10good_0/9good_1/8good_1/7good_1/6good_0/m1_14_20144# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R937 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R938 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R939 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7504 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7505 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7506 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7507 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7508 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7509 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7510 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7511 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7512 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7513 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7514 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7515 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7516 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7517 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7518 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7519 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7520 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7521 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7522 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7523 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7524 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7525 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7526 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7527 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R940 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R941 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R942 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R943 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7528 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7529 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7530 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7531 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7532 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7533 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7534 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7535 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7536 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7537 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7538 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7539 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7540 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7541 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7542 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7543 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7544 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7545 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7546 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7547 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7548 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7549 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7550 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7551 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7552 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7553 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7554 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7555 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7556 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7557 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7558 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7559 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7560 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7561 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7562 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7563 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7564 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7565 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7566 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7567 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R944 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R945 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R946 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R947 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7568 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7569 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7570 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7571 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7572 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7573 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7574 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7575 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7576 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7577 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7578 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7579 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7580 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7581 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7582 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7583 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7584 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7585 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7586 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7587 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7588 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7589 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7590 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7591 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R948 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R949 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R950 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_66618_22# sky130_fd_pr__res_generic_po w=66 l=342
R951 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7592 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7593 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7594 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7595 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7596 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7597 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7598 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7599 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7600 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7601 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7602 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7603 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7604 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7605 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7606 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7607 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7608 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7609 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7610 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7611 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7612 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7613 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7614 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7615 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7616 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7617 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7618 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7619 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7620 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7621 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7622 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7623 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R952 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R953 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R954 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R955 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7624 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7625 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7626 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7627 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7628 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7629 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7630 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7631 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7632 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7633 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7634 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7635 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7636 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7637 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7638 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7639 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7640 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7641 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7642 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7643 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7644 vdda1 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7645 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7646 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7647 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R956 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R957 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R958 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R959 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7648 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_29_719# io_in[6] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7649 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/m1_18694_42308# 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# sky130_fd_pr__pfet_01v8 w=84 l=30
X7650 10good_0/9good_1/8good_1/m1_18694_42308# 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7651 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7652 vdda1 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7653 vdda1 io_in[6] 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7654 10good_0/9good_1/8good_1/m1_18694_42308# 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# 10good_0/9good_1/8good_1/m1_18694_42308# sky130_fd_pr__pfet_01v8 w=84 l=30
X7655 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# 10good_0/9good_1/8good_1/7good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/m1_18694_42308# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7656 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# io_in[5] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7657 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X7658 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7659 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7660 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7661 vdda1 io_in[5] 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7662 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# sky130_fd_pr__pfet_01v8 w=84 l=30
X7663 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7664 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7665 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7666 10good_0/9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7667 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7668 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7669 vdda1 io_in[4] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7670 10good_0/9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_4002_19952# sky130_fd_pr__pfet_01v8 w=84 l=30
X7671 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_4002_19952# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7672 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7673 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7674 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7675 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7676 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7677 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7678 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X7679 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7680 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7681 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7682 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7683 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7684 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7685 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7686 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7687 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7688 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7689 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7690 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7691 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7692 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7693 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7694 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7695 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7696 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7697 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7698 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7699 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7700 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7701 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7702 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7703 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7704 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7705 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7706 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7707 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7708 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7709 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7710 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7711 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R960 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R961 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R962 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R963 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7712 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7713 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7714 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7715 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7716 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7717 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7718 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7719 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7720 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7721 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7722 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7723 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7724 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7725 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7726 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7727 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7728 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7729 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7730 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7731 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7732 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7733 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7734 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7735 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R964 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R965 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R966 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R967 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7736 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7737 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7738 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7739 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7740 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7741 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7742 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7743 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7744 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7745 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7746 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/m1_76798_18# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7747 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7748 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7749 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7750 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/m1_76798_18# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7751 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7752 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7753 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7754 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7755 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7756 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7757 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7758 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7759 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7760 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7761 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7762 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7763 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7764 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7765 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7766 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7767 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R968 10good_0/m1_76798_18# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R969 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R970 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R971 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7768 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7769 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7770 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7771 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7772 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7773 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7774 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7775 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7776 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7777 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7778 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7779 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7780 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7781 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7782 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7783 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7784 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7785 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7786 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7787 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7788 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7789 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7790 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7791 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R972 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R973 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R974 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R975 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7792 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7793 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7794 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7795 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7796 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7797 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7798 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7799 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7800 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7801 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7802 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7803 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7804 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7805 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7806 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7807 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7808 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7809 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7810 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7811 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7812 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7813 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7814 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7815 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7816 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7817 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7818 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7819 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7820 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7821 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7822 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7823 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7824 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7825 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7826 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7827 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7828 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7829 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7830 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7831 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R976 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R977 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R978 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R979 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7832 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7833 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7834 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7835 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7836 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7837 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7838 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7839 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7840 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7841 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7842 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7843 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7844 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7845 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7846 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7847 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7848 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7849 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7850 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7851 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7852 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7853 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7854 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7855 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R980 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R981 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R982 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_14_20144# sky130_fd_pr__res_generic_po w=66 l=342
R983 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7856 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7857 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7858 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7859 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7860 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7861 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7862 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7863 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7864 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7865 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7866 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7867 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7868 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7869 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7870 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7871 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7872 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7873 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7874 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7875 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7876 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7877 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7878 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7879 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7880 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7881 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7882 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7883 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7884 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7885 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7886 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7887 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R984 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R985 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R986 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R987 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7888 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7889 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7890 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7891 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7892 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7893 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7894 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7895 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7896 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7897 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7898 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7899 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7900 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7901 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7902 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7903 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7904 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7905 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7906 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7907 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7908 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7909 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7910 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7911 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R988 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R989 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R990 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R991 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7912 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# io_in[4] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7913 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X7914 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7915 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7916 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7917 vdda1 io_in[4] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7918 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# sky130_fd_pr__pfet_01v8 w=84 l=30
X7919 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7920 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7921 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7922 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7923 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7924 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7925 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7926 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# sky130_fd_pr__pfet_01v8 w=84 l=30
X7927 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7928 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7929 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7930 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7931 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7932 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7933 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7934 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X7935 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7936 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7937 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7938 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7939 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7940 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7941 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7942 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7943 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7944 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7945 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7946 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7947 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7948 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7949 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7950 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7951 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7952 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7953 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7954 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7955 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7956 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7957 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7958 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X7959 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R992 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R993 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R994 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R995 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7960 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7961 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7962 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7963 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7964 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7965 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7966 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7967 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7968 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7969 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X7970 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7971 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7972 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7973 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7974 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7975 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7976 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7977 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X7978 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7979 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7980 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7981 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7982 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7983 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R996 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R997 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R998 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R999 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X7984 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7985 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X7986 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7987 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7988 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7989 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7990 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X7991 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7992 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7993 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X7994 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_14_20144# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7995 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X7996 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7997 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X7998 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_14_20144# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X7999 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8000 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8001 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8002 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8003 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8004 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8005 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8006 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8007 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8008 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8009 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8010 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8011 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8012 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8013 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8014 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X8015 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R1000 10good_0/9good_1/8good_1/7good_1/6good_1/m1_14_20144# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R1001 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R1002 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R1003 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X8016 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8017 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8018 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8019 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8020 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8021 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8022 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8023 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8024 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8025 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8026 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8027 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8028 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8029 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8030 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8031 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8032 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8033 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8034 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8035 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8036 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8037 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8038 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8039 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R1004 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R1005 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R1006 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R1007 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_0/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X8040 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# io_in[3] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8041 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X8042 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8043 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8044 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8045 vdda1 io_in[3] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8046 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# sky130_fd_pr__pfet_01v8 w=84 l=30
X8047 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8048 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8049 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8050 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8051 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8052 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8053 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8054 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# sky130_fd_pr__pfet_01v8 w=84 l=30
X8055 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3500_5610# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8056 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8057 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8058 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8059 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8060 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8061 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8062 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8063 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8064 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8065 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8066 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8067 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8068 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8069 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8070 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8071 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8072 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8073 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8074 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8075 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8076 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8077 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8078 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X8079 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R1008 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R1009 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R1010 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R1011 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X8080 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8081 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8082 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8083 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8084 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8085 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8086 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8087 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8088 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8089 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8090 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8091 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8092 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8093 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8094 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8095 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8096 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8097 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8098 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8099 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8100 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8101 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8102 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8103 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R1012 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R1013 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R1014 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_700# 10good_0/m1_71736_52# sky130_fd_pr__res_generic_po w=66 l=342
R1015 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X8104 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# io_in[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8105 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8106 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8107 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8108 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8109 vdda1 io_in[2] 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8110 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# sky130_fd_pr__pfet_01v8 w=84 l=30
X8111 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8112 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8113 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8114 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8115 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8116 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8117 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8118 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8119 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8120 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8121 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8122 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8123 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8124 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8125 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8126 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8127 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8128 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8129 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8130 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8131 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8132 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8133 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8134 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# sky130_fd_pr__pfet_01v8 w=84 l=30
X8135 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3752_2110# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R1016 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R1017 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R1018 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R1019 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_0/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X8136 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8137 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__pfet_01v8 w=84 l=30
X8138 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8139 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8140 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8141 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8142 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# sky130_fd_pr__pfet_01v8 w=84 l=30
X8143 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_1/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8144 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_32342_44672# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8145 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__pfet_01v8 w=84 l=30
X8146 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8147 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8148 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8149 vdda1 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8150 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8151 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8152 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/m1_32720_44664# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8153 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# sky130_fd_pr__pfet_01v8 w=84 l=30
X8154 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8155 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8156 vdda1 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8157 vdda1 10good_0/9good_1/m1_32720_44664# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8158 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1880_n536# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# sky130_fd_pr__pfet_01v8 w=84 l=30
X8159 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/m1_1892_666# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/Sw-1_2/li_126_470# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/m1_3532_3020# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
R1020 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n930# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# sky130_fd_pr__res_generic_po w=66 l=342
R1021 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# sky130_fd_pr__res_generic_po w=66 l=342
R1022 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_700# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_1/2good_0/li_n184_n930# sky130_fd_pr__res_generic_po w=66 l=342
R1023 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n184_n588# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/3good_0/2good_1/li_n188_368# sky130_fd_pr__res_generic_po w=66 l=342
X8160 10good_0/9good_1/8good_1/Sw-1_0/li_29_719# io_in[7] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8161 10good_0/9good_1/8good_1/m1_8774_43264# 10good_0/9good_1/8good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_38716_44140# 10good_0/9good_1/8good_1/m1_8774_43264# sky130_fd_pr__pfet_01v8 w=84 l=30
X8162 10good_0/9good_1/m1_38716_44140# 10good_0/9good_1/8good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/m1_18694_42308# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8163 10good_0/9good_1/8good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8164 vdda1 10good_0/9good_1/8good_1/Sw-1_0/li_29_719# 10good_0/9good_1/8good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8165 vdda1 io_in[7] 10good_0/9good_1/8good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8166 10good_0/9good_1/m1_38716_44140# 10good_0/9good_1/8good_1/Sw-1_0/li_126_470# 10good_0/9good_1/8good_1/m1_18694_42308# 10good_0/9good_1/m1_38716_44140# sky130_fd_pr__pfet_01v8 w=84 l=30
X8167 10good_0/9good_1/8good_1/m1_8774_43264# 10good_0/9good_1/8good_1/Sw-1_0/li_126_470# 10good_0/9good_1/m1_38716_44140# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8168 10good_0/9good_1/Sw-1_0/li_29_719# io_in[8] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8169 10good_0/9good_1/m1_19068_42976# 10good_0/9good_1/Sw-1_0/li_29_719# 10good_0/m1_78452_45530# 10good_0/9good_1/m1_19068_42976# sky130_fd_pr__pfet_01v8 w=84 l=30
X8170 10good_0/m1_78452_45530# 10good_0/9good_1/Sw-1_0/li_29_719# 10good_0/9good_1/m1_38716_44140# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8171 10good_0/9good_1/Sw-1_0/li_126_470# 10good_0/9good_1/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8172 vdda1 10good_0/9good_1/Sw-1_0/li_29_719# 10good_0/9good_1/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8173 vdda1 io_in[8] 10good_0/9good_1/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8174 10good_0/m1_78452_45530# 10good_0/9good_1/Sw-1_0/li_126_470# 10good_0/9good_1/m1_38716_44140# 10good_0/m1_78452_45530# sky130_fd_pr__pfet_01v8 w=84 l=30
X8175 10good_0/9good_1/m1_19068_42976# 10good_0/9good_1/Sw-1_0/li_126_470# 10good_0/m1_78452_45530# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8176 10good_0/Sw-1_0/li_29_719# io_in[9] vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8177 10good_0/m1_39076_44800# 10good_0/Sw-1_0/li_29_719# 10good_0/Sw-1_0/w_1442_592# 10good_0/m1_39076_44800# sky130_fd_pr__pfet_01v8 w=84 l=30
X8178 10good_0/Sw-1_0/w_1442_592# 10good_0/Sw-1_0/li_29_719# 10good_0/m1_78452_45530# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8179 10good_0/Sw-1_0/li_126_470# 10good_0/Sw-1_0/li_29_719# vssa1 vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
X8180 vdda1 10good_0/Sw-1_0/li_29_719# 10good_0/Sw-1_0/li_126_470# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8181 vdda1 io_in[9] 10good_0/Sw-1_0/li_29_719# vdda1 sky130_fd_pr__pfet_01v8 w=84 l=30
X8182 10good_0/Sw-1_0/w_1442_592# 10good_0/Sw-1_0/li_126_470# 10good_0/m1_78452_45530# 10good_0/Sw-1_0/w_1442_592# sky130_fd_pr__pfet_01v8 w=84 l=30
X8183 10good_0/m1_39076_44800# 10good_0/Sw-1_0/li_126_470# 10good_0/Sw-1_0/w_1442_592# vssa1 sky130_fd_pr__nfet_01v8 w=84 l=30
C0 10good_0/9good_1/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 3.90fF
C1 vdda1 10good_0/9good_0/m1_32720_44664# 25.95fF
C2 io_in[3] io_in[5] 27.75fF
C3 10good_0/9good_1/8good_0/7good_1/6good_0/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 3.90fF
C4 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 2.83fF
C5 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# 3.52fF
C6 vdda2 vssd1 100.22fF
C7 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# 10good_0/m1_51780_62# 3.12fF
C8 io_in[5] io_in[4] 180.16fF
C9 10good_0/9good_0/8good_0/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 3.90fF
C10 chip-w-opamp_0/pass-gate-inv-2_1/in_2 chip-w-opamp_0/pass-gate-inv-2_2/in_2 2.03fF
C11 io_in[3] io_in[1] 28.04fF
C12 10good_0/m1_61528_92# 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# 3.32fF
C13 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 2.60fF
C14 10good_0/9good_0/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 3.90fF
C15 analog_io[6] analog_io[11] 2.35fF
C16 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 2.60fF
C17 analog_io[6] analog_io[10] 2.31fF
C18 io_in[3] io_in[4] 376.65fF
C19 10good_0/9good_1/m1_32342_44672# io_in[5] 7.88fF
C20 vssa2 vssd1 97.44fF
C21 vssd2 vccd2 908.10fF
C22 analog_io[12] chip-w-opamp_0/neuron-labeled-extended-opamp_1/v 3.62fF
C23 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 2.60fF
C24 10good_0/m1_56844_12# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 2.55fF
C25 vdda2 vccd1 100.22fF
C26 io_in[5] io_in[2] 2.97fF
C27 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# 6.45fF
C28 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 3.52fF
C29 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 2.83fF
C30 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_4002_19952# 3.90fF
C31 analog_io[7] analog_io[9] 8.69fF
C32 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 3.90fF
C33 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 2.60fF
C34 10good_0/9good_0/m1_32720_44664# 10good_0/9good_0/m1_32342_44672# 17.70fF
C35 io_in[3] io_in[2] 367.30fF
C36 io_in[1] io_in[2] 167.69fF
C37 10good_0/9good_0/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 3.90fF
C38 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# 6.45fF
C39 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/m1_8436_40544# 6.45fF
C40 chip-w-opamp_0/neuron-labeled-extended-opamp_1/v chip-w-opamp_0/neuron-labeled-extended-opamp_1/u 3.65fF
C41 vssa2 vccd1 97.44fF
C42 vssd2 vssd1 97.44fF
C43 analog_io[10] analog_io[11] 25.85fF
C44 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 2.60fF
C45 vdda1 io_in[5] 10.31fF
C46 analog_io[6] analog_io[24] 4.70fF
C47 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C48 io_in[4] io_in[2] 48.97fF
C49 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 2.60fF
C50 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# 10good_0/m1_41532_78# 3.66fF
C51 analog_io[3] analog_io[4] 54.94fF
C52 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 2.60fF
C53 chip-w-opamp_0/pass-gate-inv-2_3/in_2 chip-w-opamp_0/pass-gate-inv-2_3/in_1 3.93fF
C54 analog_io[15] analog_io[16] 22.83fF
C55 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# 3.52fF
C56 10good_0/m1_56844_12# 10good_0/9good_1/8good_0/7good_1/m1_8436_40544# 22.51fF
C57 10good_0/9good_1/m1_19068_42976# 10good_0/m1_39076_44800# 4.50fF
C58 vdda1 io_in[3] 24.98fF
C59 vdda1 io_in[1] 52.64fF
C60 10good_0/9good_1/m1_32342_44672# io_in[2] 4.60fF
C61 analog_io[6] chip-w-opamp_0/neuron-labeled-extended-opamp_2/u 4.86fF
C62 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 2.83fF
C63 vdda1 io_in[4] 15.84fF
C64 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 2.83fF
C65 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_0/5good_1/m1_3814_11892# 2.60fF
C66 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 2.60fF
C67 vccd2 vssd1 822.62fF
C68 vssd2 vccd1 97.44fF
C69 io_in[8] io_in[9] 76.50fF
C70 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/m1_4396_20620# 3.52fF
C71 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 2.60fF
C72 analog_io[11] analog_io[24] 3.17fF
C73 analog_io[10] vdda1 7.65fF
C74 10good_0/9good_0/8good_1/7good_0/m1_8436_40544# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 6.45fF
C75 10good_0/9good_1/m1_32342_44672# vdda1 38.23fF
C76 10good_0/9good_0/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 2.83fF
C77 10good_0/9good_0/8good_1/7good_0/m1_4396_20620# 10good_0/m1_21660_68# 3.48fF
C78 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 2.60fF
C79 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 2.83fF
C80 analog_io[6] vdda2 4.22fF
C81 io_in[5] 10good_0/9good_0/m1_32342_44672# 7.88fF
C82 vdda1 io_in[2] 39.01fF
C83 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# 10good_0/m1_31884_48# 2.94fF
C84 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C85 vccd2 vccd1 103.01fF
C86 10good_0/m1_16966_2# 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# 26.51fF
C87 chip-w-opamp_0/pass-gate-inv-2_0/in_1 chip-w-opamp_0/pass-gate-inv-2_1/in_1 2.37fF
C88 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/m1_4396_20620# 3.52fF
C89 io_in[7] io_in[6] 93.18fF
C90 10good_0/m1_11882_62# 10good_0/9good_0/8good_0/7good_1/m1_4396_20620# 5.89fF
C91 10good_0/9good_1/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_0/5good_1/m1_4054_10970# 2.83fF
C92 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C93 chip-w-opamp_0/pass-gate-inv-2_1/in_1 chip-w-opamp_0/pass-gate-inv-2_2/in_1 2.08fF
C94 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_0/7good_1/m1_8436_40544# 6.45fF
C95 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C96 10good_0/m1_1684_72# 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# 6.48fF
C97 10good_0/m1_56844_12# 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 2.40fF
C98 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_0/m1_3768_20868# 2.83fF
C99 analog_io[3] analog_io[2] 59.93fF
C100 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_4054_10970# 2.83fF
C101 chip-w-opamp_0/neuron-labeled-extended-opamp_0/v analog_io[12] 3.62fF
C102 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 2.60fF
C103 vssd1 vccd1 903.80fF
C104 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 2.60fF
C105 analog_io[24] chip-w-opamp_0/neuron-labeled-extended-opamp_2/u 3.65fF
C106 10good_0/m1_16966_2# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 2.64fF
C107 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 2.60fF
C108 io_in[2] 10good_0/9good_0/m1_32342_44672# 4.60fF
C109 chip-w-opamp_0/pass-gate-inv-2_0/in_1 chip-w-opamp_0/pass-gate-inv-2_0/in_2 3.22fF
C110 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_3814_11892# 2.60fF
C111 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# 10good_0/m1_76798_18# 4.80fF
C112 analog_io[8] analog_io[9] 44.93fF
C113 10good_0/9good_1/8good_0/7good_0/6good_0/5good_0/m1_3814_11892# 10good_0/9good_1/8good_0/7good_0/6good_0/m1_4002_19952# 3.90fF
C114 analog_io[21] analog_io[22] 21.25fF
C115 analog_io[6] analog_io[12] 2.35fF
C116 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_3814_11892# 2.60fF
C117 10good_0/9good_1/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 2.83fF
C118 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 2.60fF
C119 10good_0/m1_11882_62# io_in[5] 5.97fF
C120 analog_io[6] chip-w-opamp_0/neuron-labeled-extended-opamp_1/v 2.91fF
C121 vdda2 vdda1 100.22fF
C122 vdda1 10good_0/9good_0/m1_32342_44672# 38.23fF
C123 analog_io[10] analog_io[9] 14.58fF
C124 io_in[5] io_in[0] 16.07fF
C125 chip-w-opamp_0/pass-gate-inv-2_1/in_2 chip-w-opamp_0/pass-gate-inv-2_1/in_1 2.93fF
C126 10good_0/9good_0/8good_0/7good_0/6good_0/m1_3768_20868# 10good_0/9good_0/8good_0/7good_0/m1_4396_20620# 3.52fF
C127 analog_io[6] chip-w-opamp_0/neuron-labeled-extended-opamp_1/u 4.86fF
C128 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/4good_1/m1_3686_4442# 2.60fF
C129 vssa2 vdda1 97.44fF
C130 io_in[1] io_in[0] 153.04fF
C131 analog_io[11] analog_io[12] 26.86fF
C132 analog_io[10] analog_io[12] 8.51fF
C133 io_in[6] io_in[5] 159.58fF
C134 10good_0/9good_1/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 3.90fF
C135 analog_io[13] analog_io[12] 7.36fF
C136 analog_io[13] analog_io[14] 14.22fF
C137 10good_0/9good_1/8good_0/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_1/m1_4054_10970# 2.83fF
C138 io_in[6] io_in[3] 2.97fF
C139 analog_io[7] analog_io[8] 45.66fF
C140 10good_0/9good_1/8good_1/7good_0/6good_1/m1_3768_20868# 10good_0/9good_1/8good_1/7good_0/m1_8436_40544# 6.45fF
C141 10good_0/9good_1/8good_1/7good_1/m1_8436_40544# 10good_0/9good_1/8good_1/7good_1/6good_1/m1_3768_20868# 6.45fF
C142 chip-w-opamp_0/pass-gate-inv-2_0/in_2 chip-w-opamp_0/pass-gate-inv-2_1/in_2 2.49fF
C143 vssd2 vdda1 824.12fF
C144 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 2.60fF
C145 analog_io[16] analog_io[17] 24.92fF
C146 io_in[6] io_in[4] 19.71fF
C147 io_in[7] io_in[5] 15.58fF
C148 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 2.60fF
C149 io_in[2] io_in[0] 25.27fF
C150 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_3814_11892# 2.60fF
C151 analog_io[12] analog_io[24] 7.53fF
C152 vdda2 vssa2 914.39fF
C153 10good_0/9good_1/8good_0/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 3.90fF
C154 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_0/4good_1/m1_3686_4442# 2.60fF
C155 io_in[6] io_in[8] 7.93fF
C156 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/4good_1/m1_3686_4442# 10good_0/9good_0/8good_0/7good_0/6good_1/5good_0/m1_3814_11892# 2.60fF
C157 10good_0/9good_1/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_0/m1_3814_11892# 3.90fF
C158 vccd2 vdda1 100.22fF
C159 vdda1 io_in[0] 77.13fF
C160 10good_0/9good_1/m1_32720_44664# io_in[3] 6.31fF
C161 10good_0/9good_0/8good_1/7good_0/6good_1/5good_1/m1_4054_10970# 10good_0/9good_0/8good_1/7good_0/6good_1/m1_3768_20868# 2.83fF
C162 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# 10good_0/m1_36912_2# 16.29fF
C163 10good_0/9good_0/8good_0/7good_1/6good_0/5good_0/m1_3814_11892# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_4002_19952# 3.90fF
C164 io_in[3] 10good_0/9good_0/m1_32720_44664# 6.31fF
C165 io_in[7] io_in[8] 129.27fF
C166 vdda2 vssd2 100.22fF
C167 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/4good_1/m1_3686_4442# 2.60fF
C168 10good_0/m1_71736_52# 10good_0/9good_1/8good_1/7good_1/m1_4396_20620# 3.17fF
C169 10good_0/9good_0/8good_1/7good_1/6good_1/m1_4002_19952# 10good_0/m1_36912_2# 4.81fF
C170 vdda1 io_in[6] 2.63fF
C171 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/m1_4396_20620# 3.52fF
C172 10good_0/9good_0/8good_1/7good_1/6good_1/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/m1_8436_40544# 6.45fF
C173 chip-w-opamp_0/pass-gate-inv-2_2/in_2 chip-w-opamp_0/pass-gate-inv-2_2/in_1 2.94fF
C174 10good_0/9good_1/m1_32342_44672# 10good_0/9good_1/m1_32720_44664# 17.70fF
C175 vssd1 vdda1 100.22fF
C176 chip-w-opamp_0/neuron-labeled-extended-opamp_0/v chip-w-opamp_0/neuron-labeled-extended-opamp_0/u 3.65fF
C177 10good_0/9good_1/8good_0/7good_1/6good_0/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 2.83fF
C178 analog_io[6] chip-w-opamp_0/neuron-labeled-extended-opamp_0/v 2.91fF
C179 10good_0/9good_1/8good_1/7good_0/6good_0/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/6good_0/5good_0/m1_3814_11892# 3.90fF
C180 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 2.60fF
C181 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/m1_3814_11892# 10good_0/9good_0/8good_1/7good_0/6good_0/5good_1/4good_1/m1_3686_4442# 2.60fF
C182 10good_0/9good_1/m1_32720_44664# io_in[2] 36.73fF
C183 vssa2 vssd2 97.44fF
C184 10good_0/9good_0/8good_0/7good_0/m1_8436_40544# 10good_0/m1_6754_8# 2.51fF
C185 10good_0/9good_0/8good_1/7good_1/6good_0/m1_4002_19952# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_0/m1_3814_11892# 3.90fF
C186 10good_0/9good_0/8good_0/7good_1/6good_1/m1_4002_19952# 10good_0/9good_0/8good_0/7good_1/6good_1/5good_0/m1_3814_11892# 3.90fF
C187 10good_0/9good_0/8good_0/7good_1/6good_0/5good_1/m1_4054_10970# 10good_0/9good_0/8good_0/7good_1/6good_0/m1_3768_20868# 2.83fF
C188 10good_0/9good_1/8good_1/7good_0/6good_1/m1_4002_19952# 10good_0/9good_1/8good_1/7good_0/6good_1/5good_0/m1_3814_11892# 3.90fF
C189 analog_io[4] analog_io[5] 46.24fF
C190 vdda2 vccd2 100.22fF
C191 io_in[7] vdda1 2.27fF
C192 io_in[2] 10good_0/9good_0/m1_32720_44664# 36.73fF
C193 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_3814_11892# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 2.60fF
C194 analog_io[6] chip-w-opamp_0/neuron-labeled-extended-opamp_0/u 4.86fF
C195 10good_0/9good_1/m1_32720_44664# vdda1 25.95fF
C196 vccd1 vdda1 100.22fF
C197 10good_0/9good_0/8good_1/7good_1/6good_0/m1_3768_20868# 10good_0/9good_0/8good_1/7good_1/6good_0/5good_1/m1_4054_10970# 2.83fF
C198 analog_io[17] analog_io[18] 27.18fF
C199 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/4good_1/m1_3686_4442# 10good_0/9good_0/8good_1/7good_1/6good_1/5good_1/m1_3814_11892# 2.60fF
C200 10good_0/m1_16966_2# 10good_0/9good_0/8good_0/7good_1/6good_1/m1_3768_20868# 2.48fF
C201 10good_0/m1_1684_72# io_in[5] 5.97fF
C202 vssa2 vccd2 97.44fF
C203 10good_0/9good_1/8good_0/7good_1/6good_1/m1_3768_20868# 10good_0/9good_1/8good_0/7good_1/6good_1/5good_1/m1_4054_10970# 2.83fF
C204 10good_0/9good_1/8good_1/7good_0/m1_4396_20620# 10good_0/9good_1/8good_1/7good_0/6good_0/m1_3768_20868# 3.52fF
Xchip-w-opamp_0 analog_io[6] analog_io[7] analog_io[8] analog_io[9] analog_io[10]
+ analog_io[11] analog_io[12] analog_io[13] analog_io[14] vdda1 vssa1 vdda2 analog_io[19]
+ analog_io[20] analog_io[21] analog_io[22] analog_io[23] analog_io[15] analog_io[16]
+ analog_io[17] analog_io[18] analog_io[1] analog_io[0] analog_io[2] analog_io[3]
+ analog_io[4] analog_io[5] analog_io[24] analog_io[26] chip-w-opamp
C205 chip-w-opamp_0/neuron-labeled-extended-opamp_2/u vssa1 2.23fF
C206 chip-w-opamp_0/neuron-labeled-extended-opamp_1/u vssa1 2.23fF
C207 chip-w-opamp_0/neuron-labeled-extended-opamp_1/v vssa1 3.05fF
C208 chip-w-opamp_0/neuron-labeled-extended-opamp_0/u vssa1 2.24fF
C209 chip-w-opamp_0/neuron-labeled-extended-opamp_0/v vssa1 4.44fF
C210 10good_0/9good_1/8good_1/m1_8774_43264# vssa1 3.98fF **FLOATING
C211 10good_0/9good_1/m1_32342_44672# vssa1 136.89fF **FLOATING
C212 10good_0/9good_1/8good_0/m1_8774_43264# vssa1 3.98fF **FLOATING
C213 10good_0/9good_0/8good_1/m1_8774_43264# vssa1 3.98fF **FLOATING
C214 10good_0/9good_0/m1_32342_44672# vssa1 136.87fF **FLOATING
C215 10good_0/9good_0/8good_0/m1_8774_43264# vssa1 3.98fF **FLOATING
.ends
