magic
tech sky130A
timestamp 1604306825
<< nwell >>
rect -67 -55 67 55
<< pmos >>
rect -20 -24 20 24
<< pdiff >>
rect -49 18 -20 24
rect -49 -18 -43 18
rect -26 -18 -20 18
rect -49 -24 -20 -18
rect 20 18 49 24
rect 20 -18 26 18
rect 43 -18 49 18
rect 20 -24 49 -18
<< pdiffc >>
rect -43 -18 -26 18
rect 26 -18 43 18
<< poly >>
rect -20 24 20 37
rect -20 -37 20 -24
<< locali >>
rect -43 18 -26 26
rect -43 -26 -26 -18
rect 26 18 43 26
rect 26 -26 43 -18
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.48 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0
string library sky130
<< end >>
