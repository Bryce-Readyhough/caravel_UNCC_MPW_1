magic
tech sky130A
timestamp 1608004133
<< metal1 >>
rect 4387 21952 4421 21979
rect 5884 21966 6423 21971
rect 5884 21960 6630 21966
rect 5821 21952 6630 21960
rect 7147 21952 7220 21965
rect 4387 21936 7220 21952
rect 4387 21915 5894 21936
rect 6383 21928 7220 21936
rect 6404 21915 7220 21928
rect 4387 21632 4421 21915
rect 6204 21896 6260 21899
rect 6204 21864 6209 21896
rect 6256 21864 6260 21896
rect 7147 21892 7220 21915
rect 6204 21856 6260 21864
rect 4394 21576 4421 21632
rect 4394 20634 4427 21576
rect 6225 21200 6255 21856
rect 6417 21825 6476 21830
rect 6417 21787 6421 21825
rect 6471 21787 6476 21825
rect 6417 21782 6476 21787
rect 6202 21190 6286 21200
rect 6429 21198 6467 21782
rect 6597 21746 6654 21751
rect 6597 21706 6603 21746
rect 6648 21706 6654 21746
rect 6597 21699 6654 21706
rect 6202 21127 6210 21190
rect 6278 21127 6286 21190
rect 6202 21121 6286 21127
rect 6408 21191 6489 21198
rect 6614 21194 6649 21699
rect 7183 21666 7206 21892
rect 6776 21647 6844 21654
rect 6776 21612 6783 21647
rect 6837 21612 6844 21647
rect 7183 21652 7383 21666
rect 7183 21622 8807 21652
rect 6776 21605 6844 21612
rect 7196 21609 7383 21622
rect 6790 21258 6822 21605
rect 6961 21552 7023 21558
rect 6961 21515 6964 21552
rect 7018 21515 7023 21552
rect 6961 21507 7023 21515
rect 6408 21130 6415 21191
rect 6482 21130 6489 21191
rect 6595 21188 6664 21194
rect 6786 21193 6827 21258
rect 6986 21217 7011 21507
rect 7140 21286 7191 21291
rect 7140 21241 7144 21286
rect 7186 21277 7191 21286
rect 7343 21289 7391 21293
rect 7343 21277 7348 21289
rect 7186 21253 7348 21277
rect 7186 21241 7191 21253
rect 7140 21236 7191 21241
rect 7343 21243 7348 21253
rect 7386 21243 7391 21289
rect 7343 21240 7391 21243
rect 6595 21135 6601 21188
rect 6658 21135 6664 21188
rect 6595 21130 6664 21135
rect 6761 21188 6849 21193
rect 6408 21123 6489 21130
rect 6761 21125 6770 21188
rect 6840 21125 6849 21188
rect 6941 21181 7018 21217
rect 6941 21133 6948 21181
rect 7010 21133 7018 21181
rect 9347 21185 9618 21192
rect 9347 21154 9621 21185
rect 6941 21125 7018 21133
rect 6761 21119 6849 21125
rect 9585 20641 9621 21154
rect 9521 20626 9626 20641
rect 9585 20625 9621 20626
<< via1 >>
rect 6209 21864 6256 21896
rect 6421 21787 6471 21825
rect 6603 21706 6648 21746
rect 6210 21127 6278 21190
rect 6783 21612 6837 21647
rect 6964 21515 7018 21552
rect 6415 21130 6482 21191
rect 7144 21241 7186 21286
rect 7348 21243 7386 21289
rect 6601 21135 6658 21188
rect 6770 21125 6840 21188
rect 6948 21133 7010 21181
<< metal2 >>
rect 6204 21897 6262 21902
rect 6204 21896 6211 21897
rect 6255 21896 6262 21897
rect 6204 21864 6209 21896
rect 6256 21864 6262 21896
rect 6204 21861 6262 21864
rect 6417 21825 6476 21830
rect 6417 21787 6421 21825
rect 6471 21787 6476 21825
rect 6417 21784 6476 21787
rect 6597 21748 6658 21753
rect 6597 21746 6604 21748
rect 6597 21706 6603 21746
rect 6649 21708 6658 21748
rect 6648 21706 6658 21708
rect 6597 21700 6658 21706
rect 6775 21649 6841 21656
rect 6775 21612 6783 21649
rect 6833 21647 6841 21649
rect 6837 21612 6841 21647
rect 6775 21604 6841 21612
rect 8463 21602 8822 21613
rect 8462 21582 8822 21602
rect 6960 21552 7023 21557
rect 6960 21515 6964 21552
rect 7018 21515 7023 21552
rect 6960 21509 7023 21515
rect 7138 21286 7192 21293
rect 7138 21241 7144 21286
rect 7186 21241 7192 21286
rect 7138 21235 7192 21241
rect 7341 21291 7407 21300
rect 7341 21289 7349 21291
rect 7341 21243 7348 21289
rect 7341 21239 7349 21243
rect 7398 21239 7407 21291
rect 7341 21233 7407 21239
rect 6196 21190 6292 21200
rect 6196 21188 6210 21190
rect 6278 21188 6292 21190
rect 6196 21118 6205 21188
rect 6282 21118 6292 21188
rect 6196 21111 6292 21118
rect 6410 21191 6489 21198
rect 6410 21130 6415 21191
rect 6482 21130 6489 21191
rect 6410 21123 6416 21130
rect 6478 21123 6489 21130
rect 6593 21188 6668 21193
rect 6593 21131 6601 21188
rect 6658 21185 6668 21188
rect 6659 21131 6668 21185
rect 6593 21124 6668 21131
rect 6761 21188 6850 21195
rect 6410 21117 6489 21123
rect 6761 21121 6770 21188
rect 6840 21184 6850 21188
rect 6843 21121 6850 21184
rect 6942 21181 7015 21186
rect 6942 21133 6948 21181
rect 7010 21133 7015 21181
rect 6942 21131 6950 21133
rect 7009 21131 7015 21133
rect 6942 21125 7015 21131
rect 6761 21114 6850 21121
rect 3652 20812 5376 20849
rect 8462 20821 8504 21582
<< via2 >>
rect 6211 21896 6255 21897
rect 6211 21867 6255 21896
rect 6423 21790 6469 21824
rect 6604 21746 6649 21748
rect 6604 21708 6648 21746
rect 6648 21708 6649 21746
rect 6783 21647 6833 21649
rect 6783 21612 6833 21647
rect 6967 21517 7016 21551
rect 7144 21241 7185 21286
rect 7349 21289 7398 21291
rect 7349 21243 7386 21289
rect 7386 21243 7398 21289
rect 7349 21239 7398 21243
rect 6205 21127 6210 21188
rect 6210 21127 6278 21188
rect 6278 21127 6282 21188
rect 6205 21118 6282 21127
rect 6416 21130 6478 21186
rect 6416 21123 6478 21130
rect 6601 21135 6658 21185
rect 6658 21135 6659 21185
rect 6601 21131 6659 21135
rect 6770 21125 6840 21184
rect 6840 21125 6843 21184
rect 6770 21121 6843 21125
rect 6950 21133 7009 21176
rect 6950 21131 7009 21133
<< metal3 >>
rect 1306 21894 1361 21906
rect 6206 21897 6261 21902
rect 6206 21894 6211 21897
rect 1306 21867 6211 21894
rect 6255 21867 6261 21897
rect 1306 21863 6261 21867
rect 737 20627 786 20628
rect 1306 20627 1361 21863
rect 1447 21824 6475 21829
rect 1447 21821 6423 21824
rect 737 20600 1361 20627
rect 1419 21790 6423 21821
rect 6469 21790 6475 21824
rect 1419 21787 6475 21790
rect 737 20577 1355 20600
rect 737 20220 786 20577
rect 1419 20479 1476 21787
rect 1575 21748 6658 21755
rect 1575 21741 6604 21748
rect 888 20458 1476 20479
rect 1546 21708 6604 21741
rect 6649 21708 6658 21748
rect 1546 21701 6658 21708
rect 888 20424 1461 20458
rect 888 20340 946 20424
rect 1546 20393 1598 21701
rect 1681 21649 6837 21653
rect 1681 21628 6783 21649
rect 1667 21612 6783 21628
rect 6833 21612 6837 21649
rect 1667 21608 6837 21612
rect 1667 20471 1735 21608
rect 1792 21557 3822 21559
rect 1792 21555 5794 21557
rect 1792 21551 7023 21555
rect 1792 21517 6967 21551
rect 7016 21517 7023 21551
rect 1792 21512 7023 21517
rect 1792 20551 1859 21512
rect 3792 21510 5794 21512
rect 1946 21431 4923 21437
rect 1946 21410 7160 21431
rect 7252 21410 7310 21430
rect 1946 21358 7310 21410
rect 1946 21355 7160 21358
rect 1952 20657 2031 21355
rect 4183 21349 7160 21355
rect 7060 21346 7139 21349
rect 6970 21290 7158 21291
rect 3360 21286 7190 21290
rect 3357 21241 7144 21286
rect 7185 21241 7190 21286
rect 3357 21237 7190 21241
rect 3357 20601 3407 21237
rect 7002 21236 7190 21237
rect 6193 21188 6294 21200
rect 6193 21118 6205 21188
rect 6282 21118 6294 21188
rect 6193 21100 6294 21118
rect 6405 21186 6490 21197
rect 6405 21123 6416 21186
rect 6478 21123 6490 21186
rect 6405 21103 6490 21123
rect 6588 21185 6669 21193
rect 6588 21131 6601 21185
rect 6659 21146 6669 21185
rect 6761 21184 6853 21197
rect 6659 21131 6692 21146
rect 6208 20630 6279 21100
rect 3357 20561 3491 20601
rect 5746 20598 6289 20630
rect 3359 20554 3491 20561
rect 5739 20573 6289 20598
rect 5739 20219 5803 20573
rect 6426 20506 6483 21103
rect 6588 21089 6692 21131
rect 6761 21121 6770 21184
rect 6843 21121 6853 21184
rect 6761 21107 6853 21121
rect 6938 21176 7019 21182
rect 6938 21131 6950 21176
rect 7009 21131 7019 21176
rect 6938 21116 7019 21131
rect 6651 20717 6692 21089
rect 6785 21069 6846 21107
rect 6784 21060 6846 21069
rect 6908 21078 7019 21116
rect 6784 20918 6837 21060
rect 6651 20664 6710 20717
rect 6009 20491 6486 20506
rect 5994 20465 6486 20491
rect 5994 20454 6051 20465
rect 5986 20426 6051 20454
rect 5986 20371 6047 20426
rect 6665 20390 6710 20664
rect 6784 20491 6839 20918
rect 6908 20587 6990 21078
rect 7252 20875 7310 21358
rect 7343 21296 7413 21303
rect 7487 21296 7539 21303
rect 7343 21291 7539 21296
rect 7343 21239 7349 21291
rect 7398 21239 7539 21291
rect 7343 21233 7413 21239
rect 7064 20860 7315 20875
rect 7060 20807 7315 20860
rect 7060 20671 7139 20807
rect 7487 20703 7539 21239
rect 7487 20654 8610 20703
rect 8558 20549 8604 20654
<< metal4 >>
rect 8921 20343 8970 21232
rect 3803 20291 5579 20343
rect 8913 20329 8970 20343
rect 8913 20262 8956 20329
use 7good  7good_0
timestamp 1608004133
transform 1 0 0 0 1 28
box -1 -28 4820 20841
use 7good  7good_1
timestamp 1608004133
transform 1 0 5108 0 1 20
box -1 -28 4820 20841
use Sw-1  Sw-1_0
timestamp 1608004133
transform 1 0 8660 0 1 21115
box -70 45 891 509
<< end >>
