magic
tech sky130A
timestamp 1607400580
<< metal1 >>
rect 2192 15324 2211 15325
rect 2174 15302 2211 15324
rect 2192 10466 2211 15302
rect 1884 10455 2211 10466
rect 1884 10434 2208 10455
rect 7 10072 53 10120
rect 2199 9998 2218 10001
rect 2001 9976 2218 9998
rect 2199 5223 2218 9976
rect 2175 5202 2218 5223
rect 2175 5201 2212 5202
<< metal2 >>
rect 229 10411 256 10539
rect 229 10377 1465 10411
rect 229 9965 256 10377
<< metal3 >>
rect 1952 15284 1994 19847
rect 1219 15238 2008 15284
rect 102 10494 129 10495
rect 94 9977 129 10494
rect 94 9976 121 9977
rect 887 9952 929 11331
rect 1557 10516 1596 11696
rect 988 10506 1607 10516
rect 984 10481 1607 10506
rect 984 10078 1027 10481
rect 1759 10443 1801 12677
rect 1422 10441 1804 10443
rect 1067 10420 1804 10441
rect 1063 10412 1804 10420
rect 1063 10410 1449 10412
rect 984 9807 1031 10078
rect 1063 10037 1099 10410
rect 1950 10380 1985 15238
rect 1879 10379 1985 10380
rect 1160 10362 1985 10379
rect 1155 10350 1985 10362
rect 1155 10344 1984 10350
rect 1155 10340 1909 10344
rect 1155 10045 1188 10340
rect 1062 9873 1106 10037
rect 1155 10026 1192 10045
rect 1156 9944 1192 10026
rect 1155 9937 1999 9944
rect 1155 9908 2003 9937
rect 1062 9840 1832 9873
rect 1072 9837 1832 9840
rect 984 9767 1597 9807
rect 1553 9714 1593 9767
rect 1790 9726 1827 9837
rect 1966 5173 2003 9908
rect 1222 5131 2008 5173
<< metal4 >>
rect 425 10043 478 10157
rect 425 10001 1608 10043
rect 425 9954 515 10001
rect 465 9951 515 9954
use 5good  5good_0
timestamp 1607400580
transform 1 0 -48 0 1 -616
box 47 616 2227 10768
use 5good  5good_1
timestamp 1607400580
transform 1 0 -50 0 1 9485
box 47 616 2227 10768
use Sw-1  Sw-1_0
timestamp 1607400580
transform 1 0 1308 0 1 9932
box -70 45 891 509
<< end >>
