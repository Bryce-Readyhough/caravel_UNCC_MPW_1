magic
tech sky130A
magscale 1 2
timestamp 1608024904
<< locali >>
rect -280 8384 785 8444
rect -1000 8122 -482 8173
rect -280 7850 -220 8384
rect -1846 7720 -1232 7836
rect -964 7758 -505 7800
rect -425 7790 -220 7850
rect 17755 4791 18321 4831
rect 16470 4227 16759 4277
rect 17839 3025 18613 3065
rect -262 2561 780 2621
rect -1025 2408 -547 2465
rect -1828 2018 -1256 2134
rect -262 2125 -202 2561
rect 16436 2489 16759 2539
rect -980 2052 -582 2094
rect -502 2065 -202 2125
rect 17783 1195 19121 1235
rect 16530 663 16757 713
rect 17757 -619 19621 -579
rect 16392 -1155 16757 -1105
<< viali >>
rect -1962 7720 -1846 7836
rect 18321 4791 18361 4831
rect 16420 4227 16470 4277
rect 18613 3025 18653 3065
rect -1944 2018 -1828 2134
rect 16386 2489 16436 2539
rect 19121 1195 19161 1235
rect 16480 663 16530 713
rect 19621 -619 19661 -579
rect 16342 -1155 16392 -1105
<< metal1 >>
rect -10181 16574 -8107 16684
rect -7997 16574 255 16684
rect -9418 16080 -9412 16192
rect -9300 16080 358 16192
rect -10182 15836 -5132 15948
rect -5020 15836 -238 15948
rect -10182 15586 -5584 15698
rect -5472 15586 -134 15698
rect -10207 15336 -6049 15446
rect -5939 15336 -5 15446
rect -3293 14894 -3287 15136
rect -3045 14894 4787 15136
rect 11029 14474 11477 14616
rect 11619 14474 11625 14616
rect 10302 13198 12102 13310
rect 12214 13198 12220 13310
rect 10284 12986 12522 13098
rect 12634 12986 12640 13098
rect 10252 12773 12910 12885
rect 13022 12773 13028 12885
rect -2363 12404 -2357 12646
rect -2115 12404 4807 12646
rect 10806 12561 13280 12673
rect 13392 12561 13398 12673
rect -10077 12120 -6443 12230
rect -6333 12120 47 12230
rect -10130 11892 -6876 12004
rect -6764 11892 152 12004
rect -10156 11630 -7322 11742
rect -7210 11630 -4 11742
rect -10181 10754 -8108 10864
rect -7998 10754 489 10864
rect -5142 10128 -5132 10130
rect -10078 10018 -5132 10128
rect -5020 10128 -5010 10130
rect -5020 10018 -4 10128
rect -10078 10016 -4 10018
rect -10078 9766 -5586 9878
rect -5474 9766 22 9878
rect -6058 9626 -6048 9628
rect -10077 9516 -6048 9626
rect -5936 9626 -5926 9628
rect -5936 9516 47 9626
rect -26627 9148 -26621 9230
rect -26539 9148 -24229 9230
rect -3277 9074 -3271 9316
rect -3029 9074 4787 9316
rect -20810 8302 -19858 8354
rect -19806 8302 -19800 8354
rect -25242 8062 -25236 8114
rect -25184 8062 -24284 8114
rect -1140 8052 -1011 9074
rect 11073 8654 11477 8796
rect 11619 8654 11625 8796
rect -1968 7836 -1840 7848
rect -4208 7720 -4202 7836
rect -4086 7720 -1962 7836
rect -1846 7720 -1840 7836
rect -1968 7708 -1840 7720
rect -25936 7248 -25930 7300
rect -25878 7248 -24234 7300
rect -1112 6826 -983 7553
rect 10202 7378 12066 7490
rect 12178 7378 12184 7490
rect 10436 7166 12878 7278
rect 12990 7166 12996 7278
rect 10362 6953 13688 7065
rect 13800 6953 13806 7065
rect -2363 6584 -2357 6826
rect -2115 6584 4845 6826
rect 10774 6741 14424 6853
rect 14536 6741 14542 6853
rect -9843 6406 21 6410
rect -9843 6300 -6446 6406
rect -6456 6294 -6446 6300
rect -6334 6300 21 6406
rect -6334 6294 -6324 6300
rect -6886 6184 -6876 6186
rect -9896 6074 -6876 6184
rect -6764 6184 -6754 6186
rect -6764 6074 178 6184
rect -9896 6072 178 6074
rect -9870 5912 282 5922
rect -9870 5810 -7322 5912
rect -7332 5800 -7322 5810
rect -7210 5810 282 5912
rect -7210 5800 -7200 5810
rect -9819 5036 229 5038
rect -9819 4928 -8108 5036
rect -8118 4926 -8108 4928
rect -7998 4928 229 5036
rect 12357 5008 12363 5062
rect 12417 5008 16656 5062
rect -7998 4926 -7988 4928
rect 18315 4831 18367 4843
rect 18507 4831 18513 4837
rect 18315 4791 18321 4831
rect 18361 4791 18513 4831
rect 18315 4779 18367 4791
rect 18507 4785 18513 4791
rect 18565 4785 18571 4837
rect -5142 4302 -5132 4304
rect -9768 4192 -5132 4302
rect -5020 4302 -5010 4304
rect -5020 4192 -212 4302
rect 16123 4226 16129 4278
rect 16181 4277 16187 4278
rect 16414 4277 16476 4289
rect 16181 4227 16420 4277
rect 16470 4227 16476 4277
rect 16181 4226 16187 4227
rect 16414 4215 16476 4227
rect -9768 4190 -212 4192
rect -5594 4052 -5584 4054
rect -9716 3942 -5584 4052
rect -5472 4052 -5462 4054
rect -5472 3942 -82 4052
rect 12087 3948 12093 4002
rect 12147 3948 16618 4002
rect -9716 3940 -82 3942
rect -9637 3690 -6050 3800
rect -6060 3688 -6050 3690
rect -5938 3690 -213 3800
rect -5938 3688 -5928 3690
rect -3277 3250 -3271 3492
rect -3029 3250 4845 3492
rect -1131 2357 -1001 3250
rect 13191 3242 13197 3296
rect 13251 3242 16678 3296
rect 18607 3065 18659 3077
rect 18971 3065 18977 3071
rect 18607 3025 18613 3065
rect 18653 3025 18977 3065
rect 18607 3013 18659 3025
rect 18971 3019 18977 3025
rect 19029 3019 19035 3071
rect 11073 2828 11479 2970
rect 11621 2828 11627 2970
rect 16127 2488 16133 2540
rect 16185 2539 16191 2540
rect 16380 2539 16442 2551
rect 16185 2489 16386 2539
rect 16436 2489 16442 2539
rect 16185 2488 16191 2489
rect 16380 2477 16442 2489
rect 12883 2182 12889 2236
rect 12943 2182 16660 2236
rect -1950 2134 -1822 2146
rect -4666 2018 -4660 2134
rect -4544 2018 -1944 2134
rect -1828 2018 -1822 2134
rect -1950 2006 -1822 2018
rect -1123 1002 -993 1846
rect 10936 1552 12330 1664
rect 12442 1552 12448 1664
rect 10348 1340 13158 1452
rect 13270 1340 13276 1452
rect 14003 1412 14009 1466
rect 14063 1412 16736 1466
rect 10288 1127 13968 1239
rect 14080 1127 14086 1239
rect 19115 1235 19167 1247
rect 19397 1235 19403 1241
rect 19115 1195 19121 1235
rect 19161 1195 19403 1235
rect 19115 1183 19167 1195
rect 19397 1189 19403 1195
rect 19455 1189 19461 1241
rect -2379 760 -2373 1002
rect -2131 760 4845 1002
rect 10804 915 14688 1027
rect 14800 915 14806 1027
rect 16125 662 16131 714
rect 16183 713 16189 714
rect 16474 713 16536 725
rect 16183 663 16480 713
rect 16530 663 16536 713
rect 16183 662 16189 663
rect 16474 651 16536 663
rect -9429 474 -6440 584
rect -6450 472 -6440 474
rect -6328 474 47 584
rect -6328 472 -6318 474
rect -9404 352 152 358
rect 13717 352 13723 406
rect 13777 352 16656 406
rect -9404 246 -6876 352
rect -6886 240 -6876 246
rect -6764 246 152 352
rect -6764 240 -6754 246
rect -9378 94 204 96
rect -9378 -16 -7320 94
rect -7330 -18 -7320 -16
rect -7208 -16 204 94
rect -7208 -18 -7198 -16
rect 14717 -402 14723 -348
rect 14777 -402 16756 -348
rect 19615 -579 19667 -567
rect 19863 -579 19869 -573
rect 19615 -619 19621 -579
rect 19661 -619 19869 -579
rect 19615 -631 19667 -619
rect 19863 -625 19869 -619
rect 19921 -625 19927 -573
rect 16123 -1156 16129 -1104
rect 16181 -1105 16187 -1104
rect 16336 -1105 16398 -1093
rect 16181 -1155 16342 -1105
rect 16392 -1155 16398 -1105
rect 16181 -1156 16187 -1155
rect 16336 -1167 16398 -1155
rect 14455 -1462 14461 -1408
rect 14515 -1462 16658 -1408
rect 11469 -2001 11475 -1835
rect 11641 -2001 16536 -1835
rect 16370 -2175 16536 -2001
rect 16364 -2341 16370 -2175
rect 16536 -2341 16542 -2175
rect -19918 -2652 -19912 -2487
rect -19747 -2652 -2326 -2487
rect -2161 -2652 17180 -2487
rect 17345 -2652 17351 -2487
<< via1 >>
rect -8107 16574 -7997 16684
rect -9412 16080 -9300 16192
rect -5132 15836 -5020 15948
rect -5584 15586 -5472 15698
rect -6049 15336 -5939 15446
rect -3287 14894 -3045 15136
rect 11477 14474 11619 14616
rect 12102 13198 12214 13310
rect 12522 12986 12634 13098
rect 12910 12773 13022 12885
rect -2357 12404 -2115 12646
rect 13280 12561 13392 12673
rect -6443 12120 -6333 12230
rect -6876 11892 -6764 12004
rect -7322 11630 -7210 11742
rect -8108 10754 -7998 10864
rect -5132 10018 -5020 10130
rect -5586 9766 -5474 9878
rect -6048 9516 -5936 9628
rect -26621 9148 -26539 9230
rect -3271 9074 -3029 9316
rect -19858 8302 -19806 8354
rect -25236 8062 -25184 8114
rect 11477 8654 11619 8796
rect -4202 7720 -4086 7836
rect -25930 7248 -25878 7300
rect 12066 7378 12178 7490
rect 12878 7166 12990 7278
rect 13688 6953 13800 7065
rect -2357 6584 -2115 6826
rect 14424 6741 14536 6853
rect -6446 6294 -6334 6406
rect -6876 6074 -6764 6186
rect -7322 5800 -7210 5912
rect -8108 4926 -7998 5036
rect 12363 5008 12417 5062
rect 18513 4785 18565 4837
rect -5132 4192 -5020 4304
rect 16129 4226 16181 4278
rect -5584 3942 -5472 4054
rect 12093 3948 12147 4002
rect -6050 3688 -5938 3800
rect -3271 3250 -3029 3492
rect 13197 3242 13251 3296
rect 18977 3019 19029 3071
rect 11479 2828 11621 2970
rect 16133 2488 16185 2540
rect 12889 2182 12943 2236
rect -4660 2018 -4544 2134
rect 12330 1552 12442 1664
rect 13158 1340 13270 1452
rect 14009 1412 14063 1466
rect 13968 1127 14080 1239
rect 19403 1189 19455 1241
rect -2373 760 -2131 1002
rect 14688 915 14800 1027
rect 16131 662 16183 714
rect -6440 472 -6328 584
rect 13723 352 13777 406
rect -6876 240 -6764 352
rect -7320 -18 -7208 94
rect 14723 -402 14777 -348
rect 19869 -625 19921 -573
rect 16129 -1156 16181 -1104
rect 14461 -1462 14515 -1408
rect 11475 -2001 11641 -1835
rect 16370 -2341 16536 -2175
rect -19912 -2652 -19747 -2487
rect -2326 -2652 -2161 -2487
rect 17180 -2652 17345 -2487
<< metal2 >>
rect -26621 9230 -26539 24115
rect -26621 2029 -26539 9148
rect -25930 7300 -25878 24186
rect -25930 -8282 -25878 7248
rect -25236 8114 -25184 24356
rect -25236 -8014 -25184 8062
rect -23132 -8210 -23080 24382
rect -22740 -7916 -22688 24418
rect -22360 -8478 -22308 23824
rect -21968 -8570 -21916 24184
rect -19858 8354 -19806 24142
rect -19858 -2481 -19806 8302
rect -9412 16192 -9300 22956
rect -19912 -2487 -19747 -2481
rect -19912 -2658 -19747 -2652
rect -19858 -8002 -19806 -2658
rect -9412 -6638 -9300 16080
rect -8107 16684 -7997 23225
rect -8107 10874 -7997 16574
rect -8108 10864 -7997 10874
rect -7998 10754 -7997 10864
rect -8108 10744 -7997 10754
rect -8107 5046 -7997 10744
rect -8108 5036 -7997 5046
rect -7998 4926 -7997 5036
rect -8108 4916 -7997 4926
rect -8107 -6829 -7997 4916
rect -7322 11742 -7210 23352
rect -7322 5912 -7210 11630
rect -7322 104 -7210 5800
rect -6876 12004 -6764 23274
rect -6876 6186 -6764 11892
rect -6443 12230 -6333 23243
rect -6443 6416 -6333 12120
rect -6446 6406 -6333 6416
rect -6334 6294 -6333 6406
rect -6446 6284 -6333 6294
rect -6876 352 -6764 6074
rect -7322 94 -7208 104
rect -7322 -18 -7320 94
rect -7322 -28 -7208 -18
rect -7322 -6840 -7210 -28
rect -6876 -6826 -6764 240
rect -6443 594 -6333 6284
rect -6049 15446 -5939 23273
rect -6049 9638 -5939 15336
rect -5584 15698 -5472 23274
rect -5584 9888 -5472 15586
rect -5586 9878 -5472 9888
rect -5474 9766 -5472 9878
rect -5586 9756 -5472 9766
rect -6049 9628 -5936 9638
rect -6049 9516 -6048 9628
rect -6049 9506 -5936 9516
rect -6049 3810 -5939 9506
rect -5584 4054 -5472 9756
rect -6050 3800 -5938 3810
rect -6050 3678 -5938 3688
rect -6443 584 -6328 594
rect -6443 472 -6440 584
rect -6443 462 -6328 472
rect -6443 -6811 -6333 462
rect -6049 -6811 -5939 3678
rect -5584 -6744 -5472 3942
rect -5132 15948 -5020 23370
rect -5132 10130 -5020 15836
rect -5132 4304 -5020 10018
rect -5132 -6710 -5020 4192
rect -4660 2134 -4544 23340
rect -4660 -6690 -4544 2018
rect -4202 7836 -4086 23340
rect -3271 15142 -3029 23529
rect -3287 15136 -3029 15142
rect -3045 14894 -3029 15136
rect -3287 14888 -3029 14894
rect -4202 -6690 -4086 7720
rect -3271 9316 -3029 14888
rect -3271 3492 -3029 9074
rect -3271 -6803 -3029 3250
rect -2357 12646 -2115 23529
rect -2357 6826 -2115 12404
rect -2357 1008 -2115 6584
rect -2373 1002 -2115 1008
rect -2131 760 -2115 1002
rect -2373 754 -2115 760
rect -2357 -2487 -2115 754
rect 11477 14616 11619 23765
rect 11477 8796 11619 14474
rect 12102 13310 12214 23778
rect 12102 13192 12214 13198
rect 12522 13098 12634 23778
rect 12522 12980 12634 12986
rect 12910 12885 13022 23812
rect 12910 12767 13022 12773
rect 13280 12673 13392 23778
rect 13280 12555 13392 12561
rect 11477 2976 11619 8654
rect 12066 7490 12178 7996
rect 12066 4002 12178 7378
rect 12066 3948 12093 4002
rect 12147 3948 12178 4002
rect 11477 2970 11621 2976
rect 11477 2828 11479 2970
rect 11477 2822 11621 2828
rect 11477 -1829 11619 2822
rect 12066 -616 12178 3948
rect 12330 5062 12442 7982
rect 12330 5008 12363 5062
rect 12417 5008 12442 5062
rect 12330 1664 12442 5008
rect 12330 -644 12442 1552
rect 12878 7278 12990 8018
rect 12878 2236 12990 7166
rect 12878 2182 12889 2236
rect 12943 2182 12990 2236
rect 12878 -584 12990 2182
rect 13158 3296 13270 7990
rect 13158 3242 13197 3296
rect 13251 3242 13270 3296
rect 13158 1452 13270 3242
rect 13158 -556 13270 1340
rect 13688 7065 13800 8004
rect 13688 406 13800 6953
rect 13688 352 13723 406
rect 13777 352 13800 406
rect 13688 -556 13800 352
rect 13968 1466 14080 8048
rect 13968 1412 14009 1466
rect 14063 1412 14080 1466
rect 13968 1239 14080 1412
rect 13968 -644 14080 1127
rect 14424 6853 14536 8064
rect 14424 -1408 14536 6741
rect 14424 -1462 14461 -1408
rect 14515 -1462 14536 -1408
rect 11475 -1835 11641 -1829
rect 11475 -2007 11641 -2001
rect -2357 -2652 -2326 -2487
rect -2161 -2652 -2115 -2487
rect -2357 -6803 -2115 -2652
rect 11477 -6691 11619 -2007
rect 14424 -2706 14536 -1462
rect 14688 1027 14800 8048
rect 16130 4284 16180 23987
rect 16129 4278 16181 4284
rect 16129 4220 16181 4226
rect 14688 -348 14800 915
rect 14688 -402 14723 -348
rect 14777 -402 14800 -348
rect 14688 -2698 14800 -402
rect 16130 2546 16180 4220
rect 18014 3722 18064 5387
rect 18519 4843 18559 24188
rect 18513 4837 18565 4843
rect 18513 4779 18565 4785
rect 17761 3672 18064 3722
rect 16130 2540 16185 2546
rect 16130 2488 16133 2540
rect 16130 2482 16185 2488
rect 16130 720 16180 2482
rect 18014 1956 18064 3672
rect 17759 1906 18064 1956
rect 16130 714 16183 720
rect 16130 662 16131 714
rect 16130 656 16183 662
rect 16130 -1098 16180 656
rect 18014 126 18064 1906
rect 17755 76 18064 126
rect 16129 -1104 16181 -1098
rect 16129 -1162 16181 -1156
rect 16130 -7051 16180 -1162
rect 18014 -1688 18064 76
rect 17743 -1738 18064 -1688
rect 16370 -2175 16536 -2169
rect 16536 -2341 16910 -2175
rect 17076 -2341 17085 -2175
rect 16370 -2347 16536 -2341
rect 17180 -2487 17345 -2481
rect 18014 -2487 18064 -1738
rect 17345 -2652 18064 -2487
rect 17180 -2658 17345 -2652
rect 18014 -3723 18064 -2652
rect 18519 -7062 18559 4779
rect 18983 3077 19023 24108
rect 18977 3071 19029 3077
rect 18977 3013 19029 3019
rect 18983 -6966 19023 3013
rect 19409 1247 19449 24124
rect 19403 1241 19455 1247
rect 19403 1183 19455 1189
rect 19409 -7062 19449 1183
rect 19875 -567 19915 24188
rect 19869 -573 19921 -567
rect 19869 -631 19921 -625
rect 19875 -7158 19915 -631
<< via2 >>
rect 16910 -2341 17076 -2175
<< metal3 >>
rect 17871 4376 17943 5358
rect 17797 4306 17943 4376
rect 17871 2610 17943 4306
rect 17788 2540 17943 2610
rect 17871 780 17943 2540
rect 17786 710 17943 780
rect 17871 -1034 17943 710
rect 17786 -1104 17943 -1034
rect 16905 -2175 17081 -2170
rect 17871 -2175 17943 -1104
rect 16905 -2341 16910 -2175
rect 17076 -2341 17943 -2175
rect 16905 -2346 17081 -2341
rect 17871 -3734 17943 -2341
use neuron-labeled-extended-opamp  neuron-labeled-extended-opamp_2
timestamp 1606535953
transform 1 0 694 0 1 12268
box -1114 -638 10633 4416
use one-way  one-way_1
timestamp 1606105257
transform 1 0 -543 0 1 7572
box -37 0 183 688
use neuron-labeled-extended-opamp  neuron-labeled-extended-opamp_1
timestamp 1606535953
transform 1 0 694 0 1 6448
box -1114 -638 10633 4416
use inverter  inverter_1
timestamp 1606603647
transform 1 0 -1150 0 1 7804
box -126 -478 242 448
use 2x2-array  2x2-array_0
timestamp 1608024784
transform 1 0 -23516 0 1 6758
box -968 -870 3024 2996
use pass-gate-inv-2  pass-gate-inv-2_0
timestamp 1606604430
transform 1 0 17167 0 1 3624
box -669 -156 899 1683
use pass-gate-inv-2  pass-gate-inv-2_1
timestamp 1606604430
transform 1 0 17167 0 1 1858
box -669 -156 899 1683
use pass-gate-inv-2  pass-gate-inv-2_3
timestamp 1606604430
transform 1 0 17165 0 1 -1786
box -669 -156 899 1683
use pass-gate-inv-2  pass-gate-inv-2_2
timestamp 1606604430
transform 1 0 17165 0 1 28
box -669 -156 899 1683
use one-way  one-way_0
timestamp 1606105257
transform 1 0 -618 0 1 1859
box -37 0 183 688
use neuron-labeled-extended-opamp  neuron-labeled-extended-opamp_0
timestamp 1606535953
transform 1 0 694 0 1 622
box -1114 -638 10633 4416
use inverter  inverter_0
timestamp 1606603647
transform 1 0 -1166 0 1 2098
box -126 -478 242 448
<< labels >>
flabel metal2 -8082 23014 -8034 23104 0 FreeSans 1600 0 0 0 i_bias
port 0 nsew
flabel metal2 -7298 22968 -7250 23058 0 FreeSans 1600 0 0 0 vad
port 1 nsew
flabel metal2 -6850 22780 -6802 22870 0 FreeSans 1600 0 0 0 vr
port 2 nsew
flabel metal2 -6422 22634 -6374 22724 0 FreeSans 1600 0 0 0 vk
port 3 nsew
flabel metal2 -6026 23086 -5978 23176 0 FreeSans 1600 0 0 0 vth
port 4 nsew
flabel metal2 -5548 22932 -5500 23022 0 FreeSans 1600 0 0 0 vw
port 5 nsew
flabel metal2 -5104 22760 -5056 22850 0 FreeSans 1600 0 0 0 vau
port 6 nsew
flabel metal2 -4626 23074 -4578 23164 0 FreeSans 1600 0 0 0 vsyn0
port 7 nsew
flabel metal2 -4168 22878 -4120 22968 0 FreeSans 1600 0 0 0 vsyn1
port 8 nsew
flabel metal2 -3198 23286 -3150 23376 0 FreeSans 1600 0 0 0 vdd
port 9 nsew
flabel metal2 -2292 23270 -2244 23360 0 FreeSans 1600 0 0 0 vss
port 10 nsew
flabel metal2 11518 23554 11566 23644 0 FreeSans 1600 0 0 0 vdd_aux
port 11 nsew
flabel metal2 16144 23856 16164 23920 0 FreeSans 1600 0 0 0 sel
port 12 nsew
flabel metal2 18530 24070 18550 24134 0 FreeSans 1600 0 0 0 v_syn
port 13 nsew
flabel metal2 18990 23874 19010 23938 0 FreeSans 1600 0 0 0 u_syn
port 14 nsew
flabel metal2 19422 23636 19442 23700 0 FreeSans 1600 0 0 0 a_syn
port 15 nsew
flabel metal2 19884 23368 19904 23432 0 FreeSans 1600 0 0 0 axon_syn
port 16 nsew
flabel metal2 12134 23300 12186 23426 0 FreeSans 1600 0 0 0 v_buff
port 17 nsew
flabel metal2 12548 22954 12600 23080 0 FreeSans 1600 0 0 0 u_buff
port 18 nsew
flabel metal2 12936 22590 12988 22716 0 FreeSans 1600 0 0 0 a_buff
port 19 nsew
flabel metal2 13316 22094 13368 22220 0 FreeSans 1600 0 0 0 axon_buff
port 20 nsew
flabel metal2 -25226 24102 -25198 24160 0 FreeSans 1600 0 0 0 WL0
port 21 nsew
flabel metal2 -25914 23916 -25886 23974 0 FreeSans 1600 0 0 0 WL1
port 22 nsew
flabel metal2 -23120 23732 -23092 23790 0 FreeSans 1600 0 0 0 BL0
port 23 nsew
flabel metal2 -22728 23472 -22700 23530 0 FreeSans 1600 0 0 0 SL0
port 24 nsew
flabel metal2 -22352 23710 -22324 23768 0 FreeSans 1600 0 0 0 BL1
port 25 nsew
flabel metal2 -21954 23602 -21926 23660 0 FreeSans 1600 0 0 0 SL1
port 26 nsew
flabel metal2 -9378 22740 -9328 22830 0 FreeSans 800 0 0 0 i_in
port 27 nsew
flabel metal2 -26602 24006 -26556 24072 0 FreeSans 800 0 0 0 nwell
port 28 nsew
<< end >>
