magic
tech sky130A
magscale 1 2
timestamp 1606512719
<< error_p >>
rect -36 91 36 97
rect -36 57 -24 91
rect -36 51 36 57
<< nmos >>
rect -40 -81 40 19
<< ndiff >>
rect -98 7 -40 19
rect -98 -69 -86 7
rect -52 -69 -40 7
rect -98 -81 -40 -69
rect 40 7 98 19
rect 40 -69 52 7
rect 86 -69 98 7
rect 40 -81 98 -69
<< ndiffc >>
rect -86 -69 -52 7
rect 52 -69 86 7
<< poly >>
rect -40 91 40 107
rect -40 57 -24 91
rect 24 57 40 91
rect -40 19 40 57
rect -40 -107 40 -81
<< polycont >>
rect -24 57 24 91
<< locali >>
rect -40 57 -24 91
rect 24 57 40 91
rect -86 7 -52 23
rect -86 -85 -52 -69
rect 52 7 86 23
rect 52 -85 86 -69
<< viali >>
rect -24 57 24 91
rect -86 -69 -52 7
rect 52 -69 86 7
<< metal1 >>
rect -36 91 36 97
rect -36 57 -24 91
rect 24 57 36 91
rect -36 51 36 57
rect -92 7 -46 19
rect -92 -69 -86 7
rect -52 -69 -46 7
rect -92 -81 -46 -69
rect 46 7 92 19
rect 46 -69 52 7
rect 86 -69 92 7
rect 46 -81 92 -69
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 0.5 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
