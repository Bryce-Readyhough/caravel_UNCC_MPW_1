* NGSPICE file created from neuron-labeled-extended-opamp.ext - technology: sky130A

* Include SkyWater sky130 device models
* .include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical__lin.spice"
* .include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical.spice"
* .include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"

.lib "/home/mhasan13/pdk/pdk-prepared/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* DC source for current measure
Vdd vdd gnd DC 0.7V
Vgnd vss gnd DC 0.0V
Vth vth gnd DC 0.1V
Vk vk gnd DC 0.15V
Vw vw gnd DC 0.18V
Vr vr gnd DC 0.25V
Vau vau gnd DC 0.7V
Vad vad gnd DC 0.0V
Vdd_aux vdd_aux gnd DC 1.8V
Ibias i_bias gnd DC 1n

* Vdd VPWR gnd DC 0.7V
* Vgnd VGND gnd DC 0.0V
* Vth vth gnd DC 0.1V
* Vk vk gnd DC 0.15V
* Vw vw gnd DC 0.01V
* Vr vr gnd DC 0.37V
* Vau vau gnd DC 0.08V
* Vad vad gnd DC 0.25V

Idc vdd v DC 10p

.subckt sky130_fd_pr__nfet_01v8_r0atdz VSUBS a_n40_n107# a_n98_n81# a_40_n81#
X0 a_40_n81# a_n40_n107# a_n98_n81# VSUBS sky130_fd_pr__nfet_01v8 w=500000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4pknhj VSUBS a_n98_n86# w_n134_n148# a_40_n86# a_n40_n112#
X0 a_40_n86# a_n40_n112# a_n98_n86# w_n134_n148# sky130_fd_pr__pfet_01v8 w=500000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4ujh9u VSUBS w_n144_n198# a_n50_n162# a_n108_n136#
+ a_50_n136#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_01v8 w=1e+06u l=500000u
.ends

.subckt pmos-diff-amp in_1 in_2 out i_bias vdd vss
Xsky130_fd_pr__nfet_01v8_r0atdz_0 vss m1_91_n137# m1_91_n137# vss sky130_fd_pr__nfet_01v8_r0atdz
Xsky130_fd_pr__nfet_01v8_r0atdz_1 vss m1_91_n137# vss out sky130_fd_pr__nfet_01v8_r0atdz
Xsky130_fd_pr__pfet_01v8_4pknhj_0 vss m1_91_n137# vdd li_184_186# in_1 sky130_fd_pr__pfet_01v8_4pknhj
Xsky130_fd_pr__pfet_01v8_4ujh9u_0 vss vdd i_bias li_184_186# vdd sky130_fd_pr__pfet_01v8_4ujh9u
Xsky130_fd_pr__pfet_01v8_4pknhj_1 vss li_184_186# vdd out in_2 sky130_fd_pr__pfet_01v8_4pknhj
Xsky130_fd_pr__pfet_01v8_4ujh9u_1 vss vdd i_bias vdd i_bias sky130_fd_pr__pfet_01v8_4ujh9u
.ends

.subckt sky130_fd_pr__nfet_01v8_dlksd1 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_s3efqo VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lca7f7 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_u061qr VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_h2n75u VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_zt2j7p VSUBS a_n98_n120# a_n40_n146# a_40_n120# w_n134_n182#
X0 a_40_n120# a_n40_n146# a_n98_n120# w_n134_n182# sky130_fd_pr__pfet_01v8 w=1.2e+06u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ckptud VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_2vaynq VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_wpylm8 VSUBS a_n388_n400# a_n330_n426# a_330_n400#
X0 a_330_n400# a_n330_n426# a_n388_n400# VSUBS sky130_fd_pr__nfet_01v8 w=4e+06u l=3.3e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_9i6r5e VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_9hqhhq VSUBS a_n498_n500# a_n440_n526# a_440_n500#
X0 a_440_n500# a_n440_n526# a_n498_n500# VSUBS sky130_fd_pr__nfet_01v8 w=5e+06u l=4.4e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_h43ndc VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_6z4qh8 VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_tb02ql VSUBS a_n618_n800# a_n560_n826# a_560_n800#
X0 a_560_n800# a_n560_n826# a_n618_n800# VSUBS sky130_fd_pr__nfet_01v8 w=8e+06u l=5.6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_zgaw3c VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt neuron-labeled VPWR VGND vth vk vw vr vau vad v u# a# axon
XM10 VGND VGND vad a# sky130_fd_pr__nfet_01v8_dlksd1
XM11 VGND v a# VGND sky130_fd_pr__nfet_01v8_s3efqo
XM1 VGND a_35_1497# v vth sky130_fd_pr__nfet_01v8_lca7f7
XM2 VGND a_35_1497# VPWR VPWR a_35_1497# sky130_fd_pr__pfet_01v8_u061qr
XM3 VGND a_35_1497# VPWR VPWR v sky130_fd_pr__pfet_01v8_h2n75u
XM4 VGND VPWR a_35_1497# axon VPWR sky130_fd_pr__pfet_01v8_zt2j7p
XM5 VGND VGND a_35_1497# axon sky130_fd_pr__nfet_01v8_ckptud
XM6 VGND vw axon VPWR u# sky130_fd_pr__pfet_01v8_2vaynq
XCu VGND VGND u# VGND sky130_fd_pr__nfet_01v8_wpylm8
XM7 VGND VGND vr u# sky130_fd_pr__nfet_01v8_9i6r5e
XCv VGND VGND v VGND sky130_fd_pr__nfet_01v8_9hqhhq
XM8 VGND v u# VGND sky130_fd_pr__nfet_01v8_h43ndc
XM9 VGND vau axon VPWR a# sky130_fd_pr__pfet_01v8_6z4qh8
XCa VGND VGND a# VGND sky130_fd_pr__nfet_01v8_tb02ql
XMk VGND v vk VGND sky130_fd_pr__nfet_01v8_zgaw3c
.ends

.subckt neuron-labeled-extended-opamp v u a vau vw vth vk vr vad vdd vss axon i_bias
+ v_buff u_buff a_buff axon_buff vdd_aux
Xpmos-diff-amp_0 v v_buff v_buff i_bias vdd_aux vss pmos-diff-amp
Xpmos-diff-amp_1 u u_buff u_buff i_bias vdd_aux vss pmos-diff-amp
Xpmos-diff-amp_2 a a_buff a_buff i_bias vdd_aux vss pmos-diff-amp
Xneuron-labeled_0 vdd vss vth vk vw vr vau vad v u a axon neuron-labeled
Xpmos-diff-amp_3 axon axon_buff axon_buff i_bias vdd_aux vss pmos-diff-amp
.ends


* instantiate the neuron for sim
Xneuron v u a vau vw vth vk vr vad vdd vss axon i_bias
+ v_buff u_buff a_buff axon_buff vdd_aux neuron-labeled-extended-opamp

.IC V(v)=0 V(u)=0 V(a)=0

.control
* Sweep tran
tran 1u 20m uic
plot v(v)
plot v(v_buff)
.endc
.end

