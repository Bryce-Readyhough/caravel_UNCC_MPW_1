magic
tech sky130A
magscale 1 2
timestamp 1607400580
<< nwell >>
rect 10 760 664 822
rect 10 758 248 760
rect 10 706 244 758
rect 10 676 34 706
rect 10 602 30 676
rect 70 664 244 706
rect 250 664 664 760
rect 70 620 664 664
rect 70 616 574 620
rect 616 616 664 620
rect 70 602 664 616
rect 10 596 28 602
rect 216 594 664 602
rect 928 594 1178 976
rect 1442 768 1688 956
rect 1538 750 1688 768
rect 1442 592 1688 750
<< pwell >>
rect 480 524 1212 528
rect 6 458 30 524
rect 6 424 34 458
rect 70 424 1212 524
rect 6 374 1212 424
rect 6 312 1214 374
rect 36 274 1214 312
rect 36 272 492 274
rect 686 272 1214 274
<< psubdiff >>
rect 256 482 352 506
rect 256 436 280 482
rect 328 436 352 482
rect 256 412 352 436
<< nsubdiff >>
rect 966 910 1076 938
rect 966 866 998 910
rect 1046 866 1076 910
rect 966 836 1076 866
rect 1500 894 1606 920
rect 1500 850 1530 894
rect 1578 850 1606 894
rect 1500 830 1606 850
rect 254 734 356 762
rect 254 690 284 734
rect 328 690 356 734
rect 254 660 356 690
<< psubdiffcont >>
rect 280 436 328 482
<< nsubdiffcont >>
rect 998 866 1046 910
rect 1530 850 1578 894
rect 284 690 328 734
<< locali >>
rect 29 891 724 937
rect 29 719 75 891
rect 126 802 272 844
rect 326 802 570 844
rect 126 732 190 802
rect 274 752 338 802
rect 266 734 346 752
rect 506 734 570 802
rect 678 736 724 891
rect 978 910 1070 930
rect 978 866 998 910
rect 1046 866 1214 910
rect 978 848 1070 866
rect 1172 832 1214 866
rect 1510 894 1598 914
rect 1510 850 1530 894
rect 1578 850 1598 894
rect 1160 822 1254 832
rect 1160 764 1178 822
rect 1236 764 1254 822
rect 1510 802 1598 850
rect 1090 758 1254 764
rect 1370 798 1598 802
rect 1370 794 1754 798
rect 1370 768 1702 794
rect 266 690 284 734
rect 328 690 346 734
rect 266 672 346 690
rect 126 564 190 662
rect 414 626 448 724
rect 678 690 984 736
rect 1090 730 1214 758
rect 402 584 412 626
rect 450 584 460 626
rect 502 592 574 678
rect 678 592 712 690
rect 950 676 984 690
rect 1044 602 1104 676
rect 126 522 140 564
rect 178 522 190 564
rect 126 470 190 522
rect 264 482 346 500
rect 264 436 280 482
rect 328 436 346 482
rect 414 444 448 584
rect 502 546 712 592
rect 502 466 574 546
rect 264 420 346 436
rect 120 368 180 386
rect 120 332 196 368
rect 298 332 342 420
rect 424 414 448 444
rect 414 396 448 414
rect 678 404 712 546
rect 762 552 1104 602
rect 762 448 822 552
rect 498 370 558 386
rect 482 368 558 370
rect 482 332 574 368
rect 120 290 576 332
rect 298 220 342 290
rect 762 246 838 394
rect 904 334 950 552
rect 1178 514 1214 730
rect 1018 478 1214 514
rect 1044 448 1110 478
rect 1090 446 1110 448
rect 1146 422 1282 428
rect 1034 384 1094 392
rect 1018 372 1094 384
rect 1146 380 1230 422
rect 1268 380 1282 422
rect 1146 378 1282 380
rect 1018 334 1110 372
rect 904 332 1110 334
rect 1370 332 1406 768
rect 1538 752 1702 768
rect 1740 752 1754 794
rect 1538 750 1754 752
rect 1446 650 1504 734
rect 1538 728 1630 750
rect 1446 608 1456 650
rect 1494 608 1504 650
rect 904 298 1406 332
rect 1368 246 1378 252
rect 296 174 364 220
rect 412 174 422 220
rect 762 210 1378 246
rect 1416 246 1426 252
rect 1538 246 1614 672
rect 1416 210 1616 246
<< viali >>
rect 272 802 326 844
rect 1178 764 1236 822
rect 412 584 450 626
rect 140 522 178 564
rect 280 436 328 482
rect 1230 380 1268 422
rect 1702 752 1740 794
rect 1456 608 1494 650
rect 364 174 412 220
rect 1378 210 1416 252
<< metal1 >>
rect -24 966 1244 1018
rect 256 930 338 938
rect 256 878 264 930
rect 330 878 338 930
rect 256 850 338 878
rect 258 844 338 850
rect 258 802 272 844
rect 326 802 338 844
rect 258 774 338 802
rect 1168 822 1244 966
rect 1168 764 1178 822
rect 1236 764 1244 822
rect 1168 746 1244 764
rect 1686 796 1756 808
rect 1686 794 1782 796
rect 1686 752 1702 794
rect 1740 752 1782 794
rect 1686 734 1756 752
rect -64 666 32 676
rect -64 602 -56 666
rect 14 642 32 666
rect 1444 650 1508 664
rect 14 626 464 642
rect 14 610 412 626
rect 14 602 32 610
rect -64 594 32 602
rect 396 584 412 610
rect 450 584 464 626
rect 1444 608 1456 650
rect 1494 608 1508 650
rect 1444 596 1508 608
rect 126 564 200 578
rect 396 570 464 584
rect 126 558 140 564
rect -22 522 140 558
rect 178 522 200 564
rect -22 518 200 522
rect -22 338 18 518
rect 126 502 200 518
rect -24 302 18 338
rect 1214 422 1282 434
rect 1214 380 1230 422
rect 1268 418 1282 422
rect 1450 418 1502 596
rect 1268 384 1502 418
rect 1268 380 1282 384
rect 1214 368 1282 380
rect -24 276 822 302
rect -20 274 822 276
rect -20 262 492 274
rect 686 262 822 274
rect 420 232 512 234
rect 348 222 512 232
rect 764 224 806 262
rect 1214 224 1254 368
rect 348 220 454 222
rect 348 174 364 220
rect 412 174 454 220
rect 348 170 454 174
rect 506 170 512 222
rect 744 184 1254 224
rect 1358 252 1434 266
rect 1358 210 1378 252
rect 1416 210 1434 252
rect 348 162 512 170
rect 348 160 440 162
rect 1358 128 1434 210
rect -22 114 1434 128
rect -22 90 1418 114
<< via1 >>
rect 264 878 330 930
rect -56 602 14 666
rect 454 170 506 222
<< metal2 >>
rect 256 930 338 982
rect 256 878 264 930
rect 330 878 338 930
rect 256 868 338 878
rect -140 674 -56 680
rect -140 666 22 674
rect -140 658 -56 666
rect -140 600 -128 658
rect -72 602 -56 658
rect 14 602 22 666
rect -72 600 22 602
rect -140 594 22 600
rect -140 590 -56 594
rect 438 302 528 312
rect 438 246 448 302
rect 514 246 528 302
rect 438 234 528 246
rect 446 222 520 234
rect 446 170 454 222
rect 506 170 520 222
rect 446 162 520 170
<< via2 >>
rect -128 600 -72 658
rect 448 246 514 302
<< metal3 >>
rect -140 658 -56 712
rect -140 600 -128 658
rect -72 600 -56 658
rect -140 592 -56 600
rect 440 310 617 313
rect 438 304 617 310
rect 438 302 538 304
rect 438 246 448 302
rect 514 246 538 302
rect 438 236 538 246
rect 608 236 617 304
rect 438 227 617 236
rect 438 160 526 227
<< via3 >>
rect 538 236 608 304
<< metal4 >>
rect 528 304 620 316
rect 528 236 538 304
rect 608 236 620 304
rect 528 166 620 236
use sky130_fd_pr__nfet_01v8_dma3uj  sky130_fd_pr__nfet_01v8_dma3uj_0
timestamp 1606234862
transform 1 0 77 0 1 277
box -57 69 141 457
use sky130_fd_pr__pfet_01v8_hf7xew  sky130_fd_pr__pfet_01v8_hf7xew_0
timestamp 1606234862
transform 1 0 125 0 1 719
box -109 -123 137 95
use sky130_fd_pr__nfet_01v8_raze6j  sky130_fd_pr__nfet_01v8_raze6j_0
timestamp 1606234862
transform 1 0 121 0 1 120
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_p8bhg1  sky130_fd_pr__nfet_01v8_p8bhg1_0
timestamp 1606234862
transform 1 0 73 0 1 99
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_j74adr  sky130_fd_pr__nfet_01v8_j74adr_0
timestamp 1606234862
transform 1 0 377 0 1 97
box 21 249 219 395
use sky130_fd_pr__pfet_01v8_b4l3oq  sky130_fd_pr__pfet_01v8_b4l3oq_0
timestamp 1606237748
transform 1 0 505 0 1 725
box -111 -127 135 91
use sky130_fd_pr__nfet_01v8_5uk7v6  sky130_fd_pr__nfet_01v8_5uk7v6_0
timestamp 1606234862
transform 1 0 277 0 1 748
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_h5gdbm  sky130_fd_pr__nfet_01v8_h5gdbm_0
timestamp 1606237748
transform 1 0 763 0 1 93
box -101 255 97 401
use sky130_fd_pr__nfet_01v8_lz0viw  sky130_fd_pr__nfet_01v8_lz0viw_0
timestamp 1606237748
transform 1 0 1047 0 1 91
box -55 255 149 401
use sky130_fd_pr__pfet_01v8_htftno  sky130_fd_pr__pfet_01v8_htftno_0
timestamp 1606240701
transform 1 0 1119 0 1 727
box -187 -133 59 85
use sky130_fd_pr__pfet_01v8_k0ujpa  sky130_fd_pr__pfet_01v8_k0ujpa_0
timestamp 1606237748
transform 1 0 1693 0 1 733
box -251 -141 -5 77
<< end >>
