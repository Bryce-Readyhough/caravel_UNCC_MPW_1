magic
tech sky130A
magscale 1 2
timestamp 1607536219
<< error_p >>
rect -7836 710700 -6596 710702
rect 11284 710700 12524 710702
rect 47284 710700 48524 710702
rect 83284 710700 84524 710702
rect 119284 710700 120524 710702
rect 155284 710700 156524 710702
rect 191284 710700 192524 710702
rect 227284 710700 228524 710702
rect 263284 710700 264524 710702
rect 299284 710700 300524 710702
rect 335284 710700 336524 710702
rect 371284 710700 372524 710702
rect 407284 710700 408524 710702
rect 443520 710700 444524 710702
rect 479284 710700 480524 710702
rect 515284 710700 516524 710702
rect 551284 710700 552524 710702
rect 590520 710700 591760 710702
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect 29284 710378 30524 710380
rect 65284 710378 66524 710380
rect 101284 710378 102524 710380
rect 137284 710378 138524 710380
rect 173284 710378 174524 710380
rect 209284 710378 210524 710380
rect 245284 710378 246524 710380
rect 281284 710378 282240 710380
rect 317284 710378 318524 710380
rect 353284 710378 354524 710380
rect 389284 710378 390524 710380
rect 425284 710378 426524 710380
rect 461284 710378 462524 710380
rect 497284 710378 498524 710380
rect 533284 710378 534524 710380
rect 569284 710378 570524 710380
rect -6916 709780 -5676 709782
rect 25684 709780 26924 709782
rect 61684 709780 62924 709782
rect 97684 709780 98924 709782
rect 133684 709780 134924 709782
rect 169684 709780 170924 709782
rect 205684 709780 206924 709782
rect 241920 709780 242924 709782
rect 277684 709780 278924 709782
rect 313684 709780 314924 709782
rect 349684 709780 350924 709782
rect 385684 709780 386924 709782
rect 421684 709780 422924 709782
rect 457684 709780 458924 709782
rect 493684 709780 494924 709782
rect 529684 709780 530924 709782
rect 565684 709780 566924 709782
rect 589600 709780 590840 709782
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect 11284 709458 12524 709460
rect 47284 709458 48524 709460
rect 83284 709458 84524 709460
rect 119284 709458 120524 709460
rect 155284 709458 156524 709460
rect 191284 709458 192524 709460
rect 227284 709458 228524 709460
rect 263284 709458 264524 709460
rect 299284 709458 300524 709460
rect 335284 709458 336524 709460
rect 371284 709458 372524 709460
rect 407284 709458 408524 709460
rect 443520 709458 444524 709460
rect 479284 709458 480524 709460
rect 515284 709458 516524 709460
rect 551284 709458 552524 709460
rect -5996 708860 -4756 708862
rect 7684 708860 8924 708862
rect 43684 708860 44924 708862
rect 79684 708860 80640 708862
rect 115684 708860 116924 708862
rect 151684 708860 152924 708862
rect 187684 708860 188924 708862
rect 223684 708860 224924 708862
rect 259684 708860 260924 708862
rect 295684 708860 296924 708862
rect 331684 708860 332924 708862
rect 367684 708860 368924 708862
rect 403684 708860 404924 708862
rect 439684 708860 440924 708862
rect 475684 708860 476924 708862
rect 511684 708860 512924 708862
rect 547684 708860 548924 708862
rect 588680 708860 589920 708862
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect 25684 708538 26924 708540
rect 61684 708538 62924 708540
rect 97684 708538 98924 708540
rect 133684 708538 134924 708540
rect 169684 708538 170924 708540
rect 205684 708538 206924 708540
rect 241920 708538 242924 708540
rect 277684 708538 278924 708540
rect 313684 708538 314924 708540
rect 349684 708538 350924 708540
rect 385684 708538 386924 708540
rect 421684 708538 422924 708540
rect 457684 708538 458924 708540
rect 493684 708538 494924 708540
rect 529684 708538 530924 708540
rect 565684 708538 566924 708540
rect -5076 707940 -3836 707942
rect 22084 707940 23324 707942
rect 58084 707940 59324 707942
rect 94084 707940 95324 707942
rect 130084 707940 131324 707942
rect 166084 707940 167324 707942
rect 202084 707940 203324 707942
rect 238084 707940 239324 707942
rect 274084 707940 275324 707942
rect 310084 707940 311324 707942
rect 346084 707940 347324 707942
rect 382084 707940 383040 707942
rect 418084 707940 419324 707942
rect 454084 707940 455324 707942
rect 490084 707940 491324 707942
rect 526084 707940 527324 707942
rect 562084 707940 563324 707942
rect 587760 707940 589000 707942
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect 7684 707618 8924 707620
rect 43684 707618 44924 707620
rect 79684 707618 80640 707620
rect 115684 707618 116924 707620
rect 151684 707618 152924 707620
rect 187684 707618 188924 707620
rect 223684 707618 224924 707620
rect 259684 707618 260924 707620
rect 295684 707618 296924 707620
rect 331684 707618 332924 707620
rect 367684 707618 368924 707620
rect 403684 707618 404924 707620
rect 439684 707618 440924 707620
rect 475684 707618 476924 707620
rect 511684 707618 512924 707620
rect 547684 707618 548924 707620
rect -4156 707020 -2916 707022
rect 4084 707020 5324 707022
rect 40320 707020 41324 707022
rect 76084 707020 77324 707022
rect 112084 707020 113324 707022
rect 148084 707020 149324 707022
rect 184084 707020 185324 707022
rect 220084 707020 221324 707022
rect 256084 707020 257324 707022
rect 292084 707020 293324 707022
rect 328084 707020 329324 707022
rect 364084 707020 365324 707022
rect 400084 707020 401324 707022
rect 436084 707020 437324 707022
rect 472084 707020 473324 707022
rect 508084 707020 509324 707022
rect 544320 707020 545324 707022
rect 580084 707020 581324 707022
rect 586840 707020 588080 707022
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect 22084 706698 23324 706700
rect 58084 706698 59324 706700
rect 94084 706698 95324 706700
rect 130084 706698 131324 706700
rect 166084 706698 167324 706700
rect 202084 706698 203324 706700
rect 238084 706698 239324 706700
rect 274084 706698 275324 706700
rect 310084 706698 311324 706700
rect 346084 706698 347324 706700
rect 382084 706698 383040 706700
rect 418084 706698 419324 706700
rect 454084 706698 455324 706700
rect 490084 706698 491324 706700
rect 526084 706698 527324 706700
rect 562084 706698 563324 706700
rect -3236 706100 -1996 706102
rect 18484 706100 19724 706102
rect 54484 706100 55724 706102
rect 90484 706100 91724 706102
rect 126484 706100 127724 706102
rect 162484 706100 163724 706102
rect 198484 706100 199724 706102
rect 234484 706100 235724 706102
rect 270484 706100 271724 706102
rect 306484 706100 307724 706102
rect 342720 706100 343724 706102
rect 378484 706100 379724 706102
rect 414484 706100 415724 706102
rect 450484 706100 451724 706102
rect 486484 706100 487724 706102
rect 522484 706100 523724 706102
rect 558484 706100 559724 706102
rect 585920 706100 587160 706102
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect 4084 705778 5324 705780
rect 40320 705778 41324 705780
rect 76084 705778 77324 705780
rect 112084 705778 113324 705780
rect 148084 705778 149324 705780
rect 184084 705778 185324 705780
rect 220084 705778 221324 705780
rect 256084 705778 257324 705780
rect 292084 705778 293324 705780
rect 328084 705778 329324 705780
rect 364084 705778 365324 705780
rect 400084 705778 401324 705780
rect 436084 705778 437324 705780
rect 472084 705778 473324 705780
rect 508084 705778 509324 705780
rect 544320 705778 545324 705780
rect 580084 705778 581324 705780
rect -2316 705180 -1076 705182
rect 484 705180 1724 705182
rect 36484 705180 37724 705182
rect 72484 705180 73724 705182
rect 108484 705180 109724 705182
rect 144484 705180 145724 705182
rect 180484 705180 181440 705182
rect 216484 705180 217724 705182
rect 252484 705180 253724 705182
rect 288484 705180 289724 705182
rect 324484 705180 325724 705182
rect 360484 705180 361724 705182
rect 396484 705180 397724 705182
rect 432484 705180 433724 705182
rect 468484 705180 469724 705182
rect 504484 705180 505724 705182
rect 540484 705180 541724 705182
rect 576484 705180 577724 705182
rect 585000 705180 586240 705182
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect 18484 704858 19724 704860
rect 54484 704858 55724 704860
rect 90484 704858 91724 704860
rect 126484 704858 127724 704860
rect 162484 704858 163724 704860
rect 198484 704858 199724 704860
rect 234484 704858 235724 704860
rect 270484 704858 271724 704860
rect 306484 704858 307724 704860
rect 342720 704858 343724 704860
rect 378484 704858 379724 704860
rect 414484 704858 415724 704860
rect 450484 704858 451724 704860
rect 486484 704858 487724 704860
rect 522484 704858 523724 704860
rect 558484 704858 559724 704860
rect 18484 -924 19724 -922
rect 54484 -924 55724 -922
rect 90484 -924 91724 -922
rect 126484 -924 127724 -922
rect 162484 -924 163724 -922
rect 198484 -924 199724 -922
rect 234484 -924 235724 -922
rect 270484 -924 271724 -922
rect 306484 -924 307724 -922
rect 342720 -924 343724 -922
rect 378484 -924 379724 -922
rect 414484 -924 415724 -922
rect 450484 -924 451724 -922
rect 486484 -924 487724 -922
rect 522484 -924 523724 -922
rect 558484 -924 559724 -922
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect -2316 -1246 -1260 -1244
rect 484 -1246 1724 -1244
rect 36484 -1246 37724 -1244
rect 72484 -1246 73724 -1244
rect 108484 -1246 109724 -1244
rect 144484 -1246 145724 -1244
rect 180484 -1246 181440 -1244
rect 216484 -1246 217724 -1244
rect 252484 -1246 253724 -1244
rect 288484 -1246 289724 -1244
rect 324484 -1246 325724 -1244
rect 360484 -1246 361724 -1244
rect 396484 -1246 397724 -1244
rect 432484 -1246 433724 -1244
rect 468484 -1246 469724 -1244
rect 504484 -1246 505724 -1244
rect 540484 -1246 541724 -1244
rect 576484 -1246 577724 -1244
rect 585000 -1246 586240 -1244
rect 4084 -1844 5324 -1842
rect 40320 -1844 41324 -1842
rect 76084 -1844 77324 -1842
rect 112084 -1844 113324 -1842
rect 148084 -1844 149324 -1842
rect 184084 -1844 185324 -1842
rect 220084 -1844 221324 -1842
rect 256084 -1844 257324 -1842
rect 292084 -1844 293324 -1842
rect 328084 -1844 329324 -1842
rect 364084 -1844 365324 -1842
rect 400084 -1844 401324 -1842
rect 436084 -1844 437324 -1842
rect 472084 -1844 473324 -1842
rect 508084 -1844 509324 -1842
rect 544320 -1844 545324 -1842
rect 580084 -1844 581324 -1842
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect -3236 -2166 -1996 -2164
rect 18484 -2166 19724 -2164
rect 54484 -2166 55724 -2164
rect 90484 -2166 91724 -2164
rect 126484 -2166 127724 -2164
rect 162484 -2166 163724 -2164
rect 198484 -2166 199724 -2164
rect 234484 -2166 235724 -2164
rect 270484 -2166 271724 -2164
rect 306484 -2166 307724 -2164
rect 342720 -2166 343724 -2164
rect 378484 -2166 379724 -2164
rect 414484 -2166 415724 -2164
rect 450484 -2166 451724 -2164
rect 486484 -2166 487724 -2164
rect 522484 -2166 523724 -2164
rect 558484 -2166 559724 -2164
rect 585920 -2166 587160 -2164
rect 22084 -2764 23324 -2762
rect 58084 -2764 59324 -2762
rect 94084 -2764 95324 -2762
rect 130084 -2764 131324 -2762
rect 166084 -2764 167324 -2762
rect 202084 -2764 203324 -2762
rect 238084 -2764 239324 -2762
rect 274084 -2764 275324 -2762
rect 310084 -2764 311324 -2762
rect 346084 -2764 347324 -2762
rect 382084 -2764 383040 -2762
rect 418084 -2764 419324 -2762
rect 454084 -2764 455324 -2762
rect 490084 -2764 491324 -2762
rect 526084 -2764 527324 -2762
rect 562084 -2764 563324 -2762
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect -4156 -3086 -2916 -3084
rect 4084 -3086 5324 -3084
rect 40320 -3086 41324 -3084
rect 76084 -3086 77324 -3084
rect 112084 -3086 113324 -3084
rect 148084 -3086 149324 -3084
rect 184084 -3086 185324 -3084
rect 220084 -3086 221324 -3084
rect 256084 -3086 257324 -3084
rect 292084 -3086 293324 -3084
rect 328084 -3086 329324 -3084
rect 364084 -3086 365324 -3084
rect 400084 -3086 401324 -3084
rect 436084 -3086 437324 -3084
rect 472084 -3086 473324 -3084
rect 508084 -3086 509324 -3084
rect 544320 -3086 545324 -3084
rect 580084 -3086 581324 -3084
rect 586840 -3086 588080 -3084
rect 7684 -3684 8924 -3682
rect 43684 -3684 44924 -3682
rect 79684 -3684 80640 -3682
rect 115684 -3684 116924 -3682
rect 151684 -3684 152924 -3682
rect 187684 -3684 188924 -3682
rect 223684 -3684 224924 -3682
rect 259684 -3684 260924 -3682
rect 295684 -3684 296924 -3682
rect 331684 -3684 332924 -3682
rect 367684 -3684 368924 -3682
rect 403684 -3684 404924 -3682
rect 439684 -3684 440924 -3682
rect 475684 -3684 476924 -3682
rect 511684 -3684 512924 -3682
rect 547684 -3684 548924 -3682
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect -5076 -4006 -3836 -4004
rect 22084 -4006 23324 -4004
rect 58084 -4006 59324 -4004
rect 94084 -4006 95324 -4004
rect 130084 -4006 131324 -4004
rect 166084 -4006 167324 -4004
rect 202084 -4006 203324 -4004
rect 238084 -4006 239324 -4004
rect 274084 -4006 275324 -4004
rect 310084 -4006 311324 -4004
rect 346084 -4006 347324 -4004
rect 382084 -4006 383040 -4004
rect 418084 -4006 419324 -4004
rect 454084 -4006 455324 -4004
rect 490084 -4006 491324 -4004
rect 526084 -4006 527324 -4004
rect 562084 -4006 563324 -4004
rect 587760 -4006 589000 -4004
rect 25684 -4604 26924 -4602
rect 61684 -4604 62924 -4602
rect 97684 -4604 98924 -4602
rect 133684 -4604 134924 -4602
rect 169684 -4604 170924 -4602
rect 205684 -4604 206924 -4602
rect 241920 -4604 242924 -4602
rect 277684 -4604 278924 -4602
rect 313684 -4604 314924 -4602
rect 349684 -4604 350924 -4602
rect 385684 -4604 386924 -4602
rect 421684 -4604 422924 -4602
rect 457684 -4604 458924 -4602
rect 493684 -4604 494924 -4602
rect 529684 -4604 530924 -4602
rect 565684 -4604 566924 -4602
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect -5996 -4926 -4756 -4924
rect 7684 -4926 8924 -4924
rect 43684 -4926 44924 -4924
rect 79684 -4926 80640 -4924
rect 115684 -4926 116924 -4924
rect 151684 -4926 152924 -4924
rect 187684 -4926 188924 -4924
rect 223684 -4926 224924 -4924
rect 259684 -4926 260924 -4924
rect 295684 -4926 296924 -4924
rect 331684 -4926 332924 -4924
rect 367684 -4926 368924 -4924
rect 403684 -4926 404924 -4924
rect 439684 -4926 440924 -4924
rect 475684 -4926 476924 -4924
rect 511684 -4926 512924 -4924
rect 547684 -4926 548924 -4924
rect 588680 -4926 589920 -4924
rect 11284 -5524 12524 -5522
rect 47284 -5524 48524 -5522
rect 83284 -5524 84524 -5522
rect 119284 -5524 120524 -5522
rect 155284 -5524 156524 -5522
rect 191284 -5524 192524 -5522
rect 227284 -5524 228524 -5522
rect 263284 -5524 264524 -5522
rect 299284 -5524 300524 -5522
rect 335284 -5524 336524 -5522
rect 371284 -5524 372524 -5522
rect 407284 -5524 408524 -5522
rect 443520 -5524 444524 -5522
rect 479284 -5524 480524 -5522
rect 515284 -5524 516524 -5522
rect 551284 -5524 552524 -5522
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect -6916 -5846 -5676 -5844
rect 25684 -5846 26924 -5844
rect 61684 -5846 62924 -5844
rect 97684 -5846 98924 -5844
rect 133684 -5846 134924 -5844
rect 169684 -5846 170924 -5844
rect 205684 -5846 206924 -5844
rect 241920 -5846 242924 -5844
rect 277684 -5846 278924 -5844
rect 313684 -5846 314924 -5844
rect 349684 -5846 350924 -5844
rect 385684 -5846 386924 -5844
rect 421684 -5846 422924 -5844
rect 457684 -5846 458924 -5844
rect 493684 -5846 494924 -5844
rect 529684 -5846 530924 -5844
rect 565684 -5846 566924 -5844
rect 589600 -5846 590840 -5844
rect 29284 -6444 30524 -6442
rect 65284 -6444 66524 -6442
rect 101284 -6444 102524 -6442
rect 137284 -6444 138524 -6442
rect 173284 -6444 174524 -6442
rect 209284 -6444 210524 -6442
rect 245284 -6444 246524 -6442
rect 281284 -6444 282240 -6442
rect 317284 -6444 318524 -6442
rect 353284 -6444 354524 -6442
rect 389284 -6444 390524 -6442
rect 425284 -6444 426524 -6442
rect 461284 -6444 462524 -6442
rect 497284 -6444 498524 -6442
rect 533284 -6444 534524 -6442
rect 569284 -6444 570524 -6442
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect -7836 -6766 -6596 -6764
rect 11284 -6766 12524 -6764
rect 47284 -6766 48524 -6764
rect 83284 -6766 84524 -6764
rect 119284 -6766 120524 -6764
rect 155284 -6766 156524 -6764
rect 191284 -6766 192524 -6764
rect 227284 -6766 228524 -6764
rect 263284 -6766 264524 -6764
rect 299284 -6766 300524 -6764
rect 335284 -6766 336524 -6764
rect 371284 -6766 372524 -6764
rect 407284 -6766 408524 -6764
rect 443520 -6766 444524 -6764
rect 479284 -6766 480524 -6764
rect 515284 -6766 516524 -6764
rect 551284 -6766 552524 -6764
rect 590520 -6766 591760 -6764
<< metal1 >>
rect 142378 275806 142532 277754
rect 142314 275784 142532 275806
rect 142314 275662 142484 275784
rect 142314 275558 142340 275662
rect 142448 275558 142484 275662
rect 142314 275530 142484 275558
rect 63662 274224 63776 274248
rect 63566 274206 63776 274224
rect 63566 274150 63576 274206
rect 63640 274152 63776 274206
rect 63640 274150 63666 274152
rect 63566 274142 63666 274150
<< via1 >>
rect 142340 275558 142448 275662
rect 63576 274150 63640 274206
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 603336 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 56754 603276 56938 603336
rect 56998 603276 57007 603336
rect 56754 602274 56866 603276
rect 121614 595400 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 121614 595340 121800 595400
rect 121860 595340 121869 595400
rect 121614 594646 121726 595340
rect 186474 589686 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 186474 589626 186660 589686
rect 186720 589626 186729 589686
rect 186474 589192 186586 589626
rect 251426 583194 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 251426 583134 251614 583194
rect 251674 583134 251683 583194
rect 251426 581996 251538 583134
rect 316286 575592 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 332056 696698 332168 696707
rect 316286 575532 316464 575592
rect 316524 575532 316533 575592
rect 316286 574432 316398 575532
rect 142076 275692 142176 278820
rect 142076 275662 142518 275692
rect 142076 275558 142340 275662
rect 142448 275558 142518 275662
rect 142076 275474 142512 275558
rect 142326 275470 142512 275474
rect 142326 275338 142350 275470
rect 142482 275338 142512 275470
rect 142326 275314 142512 275338
rect 63570 274206 63648 274214
rect 63570 274150 63576 274206
rect 63640 274150 63648 274206
rect 63570 272772 63648 274150
rect 63562 272550 63764 272772
rect 63562 272370 63592 272550
rect 63726 272370 63764 272550
rect 63562 272344 63764 272370
rect 315538 5927 315590 474312
rect 316232 52869 316284 474312
rect 318336 99769 318388 474312
rect 318728 146676 318780 474312
rect 319108 193613 319160 474312
rect 319500 240545 319552 474312
rect 332056 470694 332168 696586
rect 337266 662844 337382 662853
rect 336808 615942 336924 615951
rect 336336 568994 336448 569003
rect 335884 522082 335996 522091
rect 335419 475161 335529 475170
rect 333361 287497 333471 474312
rect 334146 334416 334258 474312
rect 334592 381348 334704 474312
rect 335025 428257 335135 474312
rect 335419 471069 335529 475051
rect 335884 470678 335996 521970
rect 336336 470944 336448 568882
rect 336808 471044 336924 615826
rect 337266 470960 337382 662728
rect 353570 653602 353682 653611
rect 335025 428138 335135 428147
rect 334592 381227 334704 381236
rect 334146 334295 334258 334304
rect 338197 318925 338439 472873
rect 338197 318674 338439 318683
rect 333361 287378 333471 287387
rect 339111 286369 339353 472273
rect 352945 355401 353087 473973
rect 353570 471344 353682 653490
rect 353990 647282 354102 647291
rect 353990 470918 354102 647170
rect 354378 640380 354490 640389
rect 354378 470022 354490 640268
rect 354748 634930 354860 634939
rect 381146 634934 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 640382 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 647280 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 653614 575930 704960
rect 575515 653470 575524 653614
rect 575668 653470 575930 653614
rect 575818 653310 575930 653470
rect 510777 647168 510786 647280
rect 510898 647168 511070 647280
rect 510958 646946 511070 647168
rect 445895 640270 445904 640382
rect 446016 640270 446210 640382
rect 446098 640102 446210 640270
rect 380941 634822 380950 634934
rect 381062 634822 381258 634934
rect 354748 470146 354860 634818
rect 381146 634578 381258 634822
rect 361324 603276 361333 603336
rect 361393 603276 361402 603336
rect 360867 595400 360927 595409
rect 360867 595331 360927 595340
rect 360441 589686 360501 589695
rect 360441 589617 360501 589626
rect 359977 583194 360037 583203
rect 359977 583125 360037 583134
rect 357584 575532 357593 575592
rect 357653 575532 357662 575592
rect 357598 471249 357648 575532
rect 359987 471714 360027 583125
rect 360451 472136 360491 589617
rect 360877 471864 360917 595331
rect 361343 471536 361383 603276
rect 352945 355250 353087 355259
rect 339111 286118 339353 286127
rect 319496 240536 319556 240545
rect 319496 240467 319556 240476
rect 319104 193604 319164 193613
rect 319104 193535 319164 193544
rect 318715 146616 318724 146676
rect 318784 146616 318793 146676
rect 318332 99760 318392 99769
rect 318332 99691 318392 99700
rect 316228 52860 316288 52869
rect 316228 52791 316288 52800
rect 315534 5918 315594 5927
rect 315534 5849 315594 5858
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 56938 603276 56998 603336
rect 121800 595340 121860 595400
rect 186660 589626 186720 589686
rect 251614 583134 251674 583194
rect 332056 696586 332168 696698
rect 316464 575532 316524 575592
rect 142350 275338 142482 275470
rect 63592 272370 63726 272550
rect 337266 662728 337382 662844
rect 336808 615826 336924 615942
rect 336336 568882 336448 568994
rect 335884 521970 335996 522082
rect 335419 475051 335529 475161
rect 353570 653490 353682 653602
rect 335025 428147 335135 428257
rect 334592 381236 334704 381348
rect 334146 334304 334258 334416
rect 338197 318683 338439 318925
rect 333361 287387 333471 287497
rect 353990 647170 354102 647282
rect 354378 640268 354490 640380
rect 575524 653470 575668 653614
rect 510786 647168 510898 647280
rect 445904 640270 446016 640382
rect 354748 634818 354860 634930
rect 380950 634822 381062 634934
rect 361333 603276 361393 603336
rect 360867 595340 360927 595400
rect 360441 589626 360501 589686
rect 359977 583134 360037 583194
rect 357593 575532 357653 575592
rect 352945 355259 353087 355401
rect 339111 286127 339353 286369
rect 319496 240476 319556 240536
rect 319104 193544 319164 193604
rect 318724 146616 318784 146676
rect 318332 99700 318392 99760
rect 316228 52800 316288 52860
rect 315534 5858 315594 5918
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696698 332428 696780
rect -960 696586 332056 696698
rect 332168 696586 332428 696698
rect -960 696540 332428 696586
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 583520 674508 584960 674748
rect -960 667844 480 668084
rect 337074 662844 584960 662916
rect 337074 662728 337266 662844
rect 337382 662728 584960 662844
rect 337074 662676 584960 662728
rect -960 653428 480 653668
rect 575519 653614 575673 653619
rect 575519 653613 575524 653614
rect 353392 653602 575524 653613
rect 353392 653490 353570 653602
rect 353682 653490 575524 653602
rect 353392 653471 575524 653490
rect 575519 653470 575524 653471
rect 575668 653613 575673 653614
rect 575668 653471 575746 653613
rect 575668 653470 575673 653471
rect 575519 653465 575673 653470
rect 583520 650980 584960 651220
rect 353985 647282 354107 647287
rect 353985 647280 353990 647282
rect 353968 647170 353990 647280
rect 354102 647280 354107 647282
rect 510781 647280 510903 647285
rect 354102 647170 510786 647280
rect 353968 647168 510786 647170
rect 510898 647168 510908 647280
rect 353985 647165 354107 647168
rect 510781 647163 510903 647168
rect 354373 640382 354495 640385
rect 445899 640382 446021 640387
rect 354324 640380 445904 640382
rect 354324 640270 354378 640380
rect 354373 640268 354378 640270
rect 354490 640270 445904 640380
rect 446016 640270 446080 640382
rect 354490 640268 354495 640270
rect 354373 640263 354495 640268
rect 445899 640265 446021 640270
rect 583520 639284 584960 639524
rect -960 639012 39992 639252
rect -960 624732 480 624972
rect -960 610316 480 610556
rect -960 595900 480 596140
rect -960 581620 480 581860
rect -960 567204 480 567444
rect -960 552924 480 553164
rect -960 538508 480 538748
rect -960 524092 480 524332
rect -960 509812 480 510052
rect -960 495396 480 495636
rect -960 480980 480 481220
rect -960 466700 480 466940
rect -960 452284 480 452524
rect -960 437868 480 438108
rect -960 423588 480 423828
rect -960 409172 480 409412
rect -960 394892 480 395132
rect -960 380476 480 380716
rect -960 366060 480 366300
rect -960 351780 480 352020
rect -960 337364 480 337604
rect -960 322948 480 323188
rect -960 308668 480 308908
rect -960 294252 480 294492
rect -960 279972 480 280212
rect 39752 272582 39992 639012
rect 354743 634934 354865 634935
rect 380945 634934 381067 634939
rect 354688 634930 380950 634934
rect 354688 634822 354748 634930
rect 354743 634818 354748 634822
rect 354860 634822 380950 634930
rect 381062 634822 381112 634934
rect 354860 634818 354865 634822
rect 354743 634813 354865 634818
rect 380945 634817 381067 634822
rect 583520 627588 584960 627828
rect 336614 615942 584960 615996
rect 336614 615826 336808 615942
rect 336924 615826 584960 615942
rect 336614 615756 584960 615826
rect 583520 604060 584960 604300
rect 56933 603336 57003 603341
rect 361328 603336 361398 603341
rect 56894 603276 56938 603336
rect 56998 603276 361333 603336
rect 361393 603276 361398 603336
rect 56933 603271 57003 603276
rect 361328 603271 361398 603276
rect 121795 595400 121865 595405
rect 360862 595400 360932 595405
rect 121774 595340 121800 595400
rect 121860 595340 360867 595400
rect 360927 595340 360932 595400
rect 121795 595335 121865 595340
rect 360862 595335 360932 595340
rect 583520 592364 584960 592604
rect 186655 589686 186725 589691
rect 360436 589686 360506 589691
rect 186618 589626 186660 589686
rect 186720 589626 360441 589686
rect 360501 589626 360506 589686
rect 186655 589621 186725 589626
rect 360436 589621 360506 589626
rect 251609 583194 251679 583199
rect 359972 583194 360042 583199
rect 251574 583134 251614 583194
rect 251674 583134 359977 583194
rect 360037 583134 360042 583194
rect 251609 583129 251679 583134
rect 359972 583129 360042 583134
rect 583520 580668 584960 580908
rect 316459 575592 316529 575597
rect 357588 575592 357658 575597
rect 316420 575532 316464 575592
rect 316524 575532 357593 575592
rect 357653 575532 357658 575592
rect 316459 575527 316529 575532
rect 357588 575527 357658 575532
rect 336118 568994 584960 569076
rect 336118 568882 336336 568994
rect 336448 568882 584960 568994
rect 336118 568836 584960 568882
rect 583520 557140 584960 557380
rect 583520 545444 584960 545684
rect 583520 533748 584960 533988
rect 335720 522082 584960 522156
rect 335720 521970 335884 522082
rect 335996 521970 584960 522082
rect 335720 521916 584960 521970
rect 583520 510220 584960 510460
rect 583520 498524 584960 498764
rect 583520 486692 584960 486932
rect 335322 475161 584960 475236
rect 335322 475051 335419 475161
rect 335529 475051 584960 475161
rect 335322 474996 584960 475051
rect 583520 463300 584960 463540
rect 583520 451604 584960 451844
rect 291924 439772 584960 440012
rect 142326 275470 142520 275502
rect 142326 275338 142350 275470
rect 142482 275338 142520 275470
rect 142326 275236 142520 275338
rect 142326 275062 142344 275236
rect 142490 275062 142520 275236
rect 142326 275044 142520 275062
rect 39752 272550 63786 272582
rect 39752 272370 63592 272550
rect 63726 272370 63786 272550
rect 39752 272342 63786 272370
rect 65590 271641 65720 273361
rect 57253 271511 65720 271641
rect -960 265556 480 265796
rect 57253 255578 57383 271511
rect 66054 270831 66220 273228
rect 60039 270665 66220 270831
rect 57253 255063 57612 255578
rect -960 251140 480 251380
rect -960 236860 480 237100
rect -960 222444 480 222684
rect -960 208028 480 208268
rect -960 193748 480 193988
rect -960 179332 480 179572
rect -960 164916 480 165156
rect -960 150636 480 150876
rect -960 136220 480 136460
rect -960 121940 480 122180
rect -960 107524 480 107764
rect -960 93108 480 93348
rect -960 78828 480 79068
rect -960 64412 480 64652
rect -960 49996 480 50236
rect -960 35716 480 35956
rect -960 21300 480 21540
rect 57372 17732 57612 255063
rect 60039 255051 60205 270665
rect 66856 270246 67000 272942
rect 63154 270102 67000 270246
rect 67756 272560 68072 272704
rect 60384 255051 60624 255070
rect 60039 254345 60624 255051
rect 60384 64652 60624 254345
rect 63154 254866 63298 270102
rect 67756 269714 67900 272560
rect 66978 269570 67900 269714
rect 68130 272330 68494 272474
rect 63154 254206 63476 254866
rect 63236 111572 63476 254206
rect 66978 254140 67122 269570
rect 68130 268124 68274 272330
rect 68556 272086 68966 272230
rect 68556 268562 68700 272086
rect 68932 271824 69432 271968
rect 68932 269018 69076 271824
rect 69376 271562 69790 271706
rect 69376 269358 69520 271562
rect 69772 271314 70222 271458
rect 69772 269702 69916 271314
rect 70222 271052 70758 271196
rect 70222 270084 70366 271052
rect 70222 269940 86682 270084
rect 69772 269558 83444 269702
rect 69376 269214 80316 269358
rect 68932 268874 77792 269018
rect 68556 268418 74446 268562
rect 68130 267980 70786 268124
rect 66978 253478 67234 254140
rect 66994 158492 67234 253478
rect 70642 253714 70786 267980
rect 70642 252794 70888 253714
rect 70648 205412 70888 252794
rect 74302 252332 74446 268418
rect 77648 253148 77792 268874
rect 80172 254108 80316 269214
rect 83300 255360 83444 269558
rect 86538 256508 86682 269940
rect 291924 256508 292164 439772
rect 334910 428257 584960 428316
rect 334910 428147 335025 428257
rect 335135 428147 584960 428257
rect 334910 428076 584960 428147
rect 583520 416380 584960 416620
rect 583520 404684 584960 404924
rect 86538 256268 292164 256508
rect 300952 392852 584960 393092
rect 86538 256222 86682 256268
rect 300952 255360 301192 392852
rect 334468 381348 584960 381396
rect 334468 381236 334592 381348
rect 334704 381236 584960 381348
rect 334468 381156 584960 381236
rect 583520 369460 584960 369700
rect 583520 357764 584960 358004
rect 352940 355401 353092 355406
rect 352940 355259 352945 355401
rect 353087 355259 353092 355401
rect 352940 355254 353092 355259
rect 352945 351927 353087 355254
rect 352945 351779 353087 351785
rect 83300 255120 301192 255360
rect 303884 345932 584960 346172
rect 83300 255092 83444 255120
rect 303884 254108 304124 345932
rect 334014 334416 584960 334476
rect 334014 334304 334146 334416
rect 334258 334304 584960 334416
rect 334014 334236 584960 334304
rect 583520 322540 584960 322780
rect 338192 318925 338444 318930
rect 338192 318683 338197 318925
rect 338439 318683 338444 318925
rect 338192 318678 338444 318683
rect 338197 316681 338439 318678
rect 338197 316433 338439 316439
rect 583520 310708 584960 310948
rect 80172 253870 304124 254108
rect 80244 253868 304124 253870
rect 306042 299012 584960 299252
rect 306042 253148 306282 299012
rect 333064 287497 584960 287556
rect 333064 287387 333361 287497
rect 333471 287387 584960 287497
rect 333064 287316 584960 287387
rect 339106 286369 339358 286374
rect 339106 286127 339111 286369
rect 339353 286127 339358 286369
rect 339106 286122 339358 286127
rect 339111 284223 339353 286122
rect 339111 283975 339353 283981
rect 583520 275620 584960 275860
rect 583520 263788 584960 264028
rect 77648 252920 306282 253148
rect 77724 252908 306282 252920
rect 74302 252092 584960 252332
rect 74302 252068 74446 252092
rect 319410 240536 584960 240636
rect 319410 240476 319496 240536
rect 319556 240476 584960 240536
rect 319410 240396 584960 240476
rect 583520 228700 584960 228940
rect 583520 216868 584960 217108
rect 70648 205172 584960 205412
rect 319026 193604 584960 193716
rect 319026 193544 319104 193604
rect 319164 193544 584960 193604
rect 319026 193476 584960 193544
rect 583520 181780 584960 182020
rect 583520 169948 584960 170188
rect 66994 158252 584960 158492
rect 318698 146676 584960 146796
rect 318698 146616 318724 146676
rect 318784 146616 584960 146676
rect 318698 146556 584960 146616
rect 583520 134724 584960 134964
rect 583520 123028 584960 123268
rect 63236 111332 584960 111572
rect 317720 99760 584960 99876
rect 317720 99700 318332 99760
rect 318392 99700 584960 99760
rect 317720 99636 584960 99700
rect 583520 87804 584960 88044
rect 583520 76108 584960 76348
rect 60384 64412 584960 64652
rect 316182 52860 584960 52956
rect 316182 52800 316228 52860
rect 316288 52800 584960 52860
rect 316182 52716 584960 52800
rect 583520 40884 584960 41124
rect 583520 29188 584960 29428
rect 57372 17492 584960 17732
rect -960 7020 480 7260
rect 314984 5918 584960 6036
rect 314984 5858 315534 5918
rect 315594 5858 584960 5918
rect 314984 5796 584960 5858
<< via3 >>
rect 142344 275062 142490 275236
rect 352945 351785 353087 351927
rect 338197 316439 338439 316681
rect 339111 283981 339353 284223
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 703520 1404 704282
rect 4404 703520 5004 706122
rect 8004 703520 8604 707962
rect 11604 703520 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 703520 19404 705202
rect 22404 703520 23004 707042
rect 26004 703520 26604 708882
rect 29604 703520 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 703520 37404 704282
rect 40404 703520 41004 706122
rect 44004 703520 44604 707962
rect 47604 703520 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 703520 55404 705202
rect 58404 703520 59004 707042
rect 62004 703520 62604 708882
rect 65604 703520 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 703520 73404 704282
rect 76404 703520 77004 706122
rect 80004 703520 80604 707962
rect 83604 703520 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 703520 91404 705202
rect 94404 703520 95004 707042
rect 98004 703520 98604 708882
rect 101604 703520 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 703520 109404 704282
rect 112404 703520 113004 706122
rect 116004 703520 116604 707962
rect 119604 703520 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 703520 127404 705202
rect 130404 703520 131004 707042
rect 134004 703520 134604 708882
rect 137604 703520 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 703520 145404 704282
rect 148404 703520 149004 706122
rect 152004 703520 152604 707962
rect 155604 703520 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 703520 163404 705202
rect 166404 703520 167004 707042
rect 170004 703520 170604 708882
rect 173604 703520 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 703520 181404 704282
rect 184404 703520 185004 706122
rect 188004 703520 188604 707962
rect 191604 703520 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 703520 199404 705202
rect 202404 703520 203004 707042
rect 206004 703520 206604 708882
rect 209604 703520 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 703520 217404 704282
rect 220404 703520 221004 706122
rect 224004 703520 224604 707962
rect 227604 703520 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 703520 235404 705202
rect 238404 703520 239004 707042
rect 242004 703520 242604 708882
rect 245604 703520 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 703520 253404 704282
rect 256404 703520 257004 706122
rect 260004 703520 260604 707962
rect 263604 703520 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 703520 271404 705202
rect 274404 703520 275004 707042
rect 278004 703520 278604 708882
rect 281604 703520 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 703520 289404 704282
rect 292404 703520 293004 706122
rect 296004 703520 296604 707962
rect 299604 703520 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 703520 307404 705202
rect 310404 703520 311004 707042
rect 314004 703520 314604 708882
rect 317604 703520 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 703520 325404 704282
rect 328404 703520 329004 706122
rect 332004 703520 332604 707962
rect 335604 703520 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 703520 343404 705202
rect 346404 703520 347004 707042
rect 350004 703520 350604 708882
rect 353604 703520 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 703520 361404 704282
rect 364404 703520 365004 706122
rect 368004 703520 368604 707962
rect 371604 703520 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 703520 379404 705202
rect 382404 703520 383004 707042
rect 386004 703520 386604 708882
rect 389604 703520 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 703520 397404 704282
rect 400404 703520 401004 706122
rect 404004 703520 404604 707962
rect 407604 703520 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 703520 415404 705202
rect 418404 703520 419004 707042
rect 422004 703520 422604 708882
rect 425604 703520 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 703520 433404 704282
rect 436404 703520 437004 706122
rect 440004 703520 440604 707962
rect 443604 703520 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 703520 451404 705202
rect 454404 703520 455004 707042
rect 458004 703520 458604 708882
rect 461604 703520 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 703520 469404 704282
rect 472404 703520 473004 706122
rect 476004 703520 476604 707962
rect 479604 703520 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 703520 487404 705202
rect 490404 703520 491004 707042
rect 494004 703520 494604 708882
rect 497604 703520 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 703520 505404 704282
rect 508404 703520 509004 706122
rect 512004 703520 512604 707962
rect 515604 703520 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 703520 523404 705202
rect 526404 703520 527004 707042
rect 530004 703520 530604 708882
rect 533604 703520 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 703520 541404 704282
rect 544404 703520 545004 706122
rect 548004 703520 548604 707962
rect 551604 703520 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 703520 559404 705202
rect 562404 703520 563004 707042
rect 566004 703520 566604 708882
rect 569604 703520 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 703520 577404 704282
rect 580404 703520 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 352944 351927 353088 351928
rect 352944 351785 352945 351927
rect 353087 351785 353088 351927
rect 352944 351784 353088 351785
rect 352945 343742 353087 351784
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 338196 316681 338440 316682
rect 338196 316439 338197 316681
rect 338439 316439 338440 316681
rect 338196 316438 338440 316439
rect 338197 312212 338439 316438
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 339110 284223 339354 284224
rect 339110 283981 339111 284223
rect 339353 283981 339354 284223
rect 339110 283980 339354 283981
rect 339111 281750 339353 283980
rect 140822 278664 141080 278678
rect 140822 278180 141670 278664
rect 140822 276188 141080 278180
rect 140696 275776 141198 276188
rect 132054 275532 141198 275776
rect 132054 275304 141168 275532
rect 132160 264340 132618 275304
rect 142130 275236 142730 275278
rect 142130 275062 142344 275236
rect 142490 275062 142730 275236
rect 132160 264072 132772 264340
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect 132172 229856 132772 264072
rect 142130 249324 142730 275062
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 142130 248724 296604 249324
rect 132172 229256 278604 229856
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 -346 1404 480
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 480
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 480
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 480
rect 18804 -1266 19404 480
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 -3106 23004 480
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 -4946 26604 480
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 480
rect 36804 -346 37404 480
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 -2186 41004 480
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 -4026 44604 480
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 480
rect 54804 -1266 55404 480
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 -3106 59004 480
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 -4946 62604 480
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 480
rect 72804 -346 73404 480
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 -2186 77004 480
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 -4026 80604 480
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 480
rect 90804 -1266 91404 480
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 -3106 95004 480
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 -4946 98604 480
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 480
rect 108804 -346 109404 480
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 -2186 113004 480
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 -4026 116604 480
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 480
rect 126804 -1266 127404 480
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 -3106 131004 480
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 -4946 134604 480
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 480
rect 144804 -346 145404 480
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 -2186 149004 480
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 -4026 152604 480
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 480
rect 162804 -1266 163404 480
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 -3106 167004 480
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 -4946 170604 480
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 480
rect 180804 -346 181404 480
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 -2186 185004 480
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 -4026 188604 480
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 480
rect 198804 -1266 199404 480
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 -3106 203004 480
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 -4946 206604 480
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 480
rect 216804 -346 217404 480
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 -2186 221004 480
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 -4026 224604 480
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 480
rect 234804 -1266 235404 480
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 -3106 239004 480
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 -4946 242604 480
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 480
rect 252804 -346 253404 480
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 -2186 257004 480
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 -4026 260604 480
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 480
rect 270804 -1266 271404 480
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 -3106 275004 480
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 -4946 278604 229256
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 480
rect 288804 -346 289404 480
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 -2186 293004 480
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 -4026 296604 248724
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 480
rect 306804 -1266 307404 480
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 -3106 311004 480
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 -4946 314604 480
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 480
rect 324804 -346 325404 480
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 -2186 329004 480
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 -4026 332604 480
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 480
rect 342804 -1266 343404 480
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 -3106 347004 480
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 -4946 350604 480
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 480
rect 360804 -346 361404 480
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 -2186 365004 480
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 -4026 368604 480
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 480
rect 378804 -1266 379404 480
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 -3106 383004 480
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 -4946 386604 480
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 480
rect 396804 -346 397404 480
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 -2186 401004 480
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 -4026 404604 480
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 480
rect 414804 -1266 415404 480
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 -3106 419004 480
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 -4946 422604 480
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 480
rect 432804 -346 433404 480
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 -2186 437004 480
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 -4026 440604 480
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 480
rect 450804 -1266 451404 480
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 -3106 455004 480
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 -4946 458604 480
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 480
rect 468804 -346 469404 480
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 -2186 473004 480
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 -4026 476604 480
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 480
rect 486804 -1266 487404 480
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 -3106 491004 480
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 -4946 494604 480
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 480
rect 504804 -346 505404 480
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 -2186 509004 480
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 -4026 512604 480
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 480
rect 522804 -1266 523404 480
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 -3106 527004 480
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 -4946 530604 480
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 480
rect 540804 -346 541404 480
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 -2186 545004 480
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 -4026 548604 480
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 480
rect 558804 -1266 559404 480
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 -3106 563004 480
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 -4946 566604 480
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 480
rect 576804 -346 577404 480
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 -2186 581004 480
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 352856 343422 353176 343742
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 338158 311892 338478 312212
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 339072 281430 339392 281750
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 590840 697276 591440 697278
rect -8436 697254 480 697276
rect -8436 697018 -7334 697254
rect -7098 697018 480 697254
rect -8436 696934 480 697018
rect -8436 696698 -7334 696934
rect -7098 696698 480 696934
rect -8436 696676 480 696698
rect 583520 697254 592360 697276
rect 583520 697018 591022 697254
rect 591258 697018 592360 697254
rect 583520 696934 592360 697018
rect 583520 696698 591022 696934
rect 591258 696698 592360 696934
rect 583520 696676 592360 696698
rect -7516 696674 -6916 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 589000 693676 589600 693678
rect -6596 693654 480 693676
rect -6596 693418 -5494 693654
rect -5258 693418 480 693654
rect -6596 693334 480 693418
rect -6596 693098 -5494 693334
rect -5258 693098 480 693334
rect -6596 693076 480 693098
rect 583520 693654 590520 693676
rect 583520 693418 589182 693654
rect 589418 693418 590520 693654
rect 583520 693334 590520 693418
rect 583520 693098 589182 693334
rect 589418 693098 590520 693334
rect 583520 693076 590520 693098
rect -5676 693074 -5076 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 587160 690076 587760 690078
rect -4756 690054 480 690076
rect -4756 689818 -3654 690054
rect -3418 689818 480 690054
rect -4756 689734 480 689818
rect -4756 689498 -3654 689734
rect -3418 689498 480 689734
rect -4756 689476 480 689498
rect 583520 690054 588680 690076
rect 583520 689818 587342 690054
rect 587578 689818 588680 690054
rect 583520 689734 588680 689818
rect 583520 689498 587342 689734
rect 587578 689498 588680 689734
rect 583520 689476 588680 689498
rect -3836 689474 -3236 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 585320 686476 585920 686478
rect -2916 686454 480 686476
rect -2916 686218 -1814 686454
rect -1578 686218 480 686454
rect -2916 686134 480 686218
rect -2916 685898 -1814 686134
rect -1578 685898 480 686134
rect -2916 685876 480 685898
rect 583520 686454 586840 686476
rect 583520 686218 585502 686454
rect 585738 686218 586840 686454
rect 583520 686134 586840 686218
rect 583520 685898 585502 686134
rect 585738 685898 586840 686134
rect 583520 685876 586840 685898
rect -1996 685874 -1396 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 591760 679276 592360 679278
rect -8436 679254 480 679276
rect -8436 679018 -8254 679254
rect -8018 679018 480 679254
rect -8436 678934 480 679018
rect -8436 678698 -8254 678934
rect -8018 678698 480 678934
rect -8436 678676 480 678698
rect 583520 679254 592360 679276
rect 583520 679018 591942 679254
rect 592178 679018 592360 679254
rect 583520 678934 592360 679018
rect 583520 678698 591942 678934
rect 592178 678698 592360 678934
rect 583520 678676 592360 678698
rect -8436 678674 -7836 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 589920 675676 590520 675678
rect -6596 675654 480 675676
rect -6596 675418 -6414 675654
rect -6178 675418 480 675654
rect -6596 675334 480 675418
rect -6596 675098 -6414 675334
rect -6178 675098 480 675334
rect -6596 675076 480 675098
rect 583520 675654 590520 675676
rect 583520 675418 590102 675654
rect 590338 675418 590520 675654
rect 583520 675334 590520 675418
rect 583520 675098 590102 675334
rect 590338 675098 590520 675334
rect 583520 675076 590520 675098
rect -6596 675074 -5996 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 588080 672076 588680 672078
rect -4756 672054 480 672076
rect -4756 671818 -4574 672054
rect -4338 671818 480 672054
rect -4756 671734 480 671818
rect -4756 671498 -4574 671734
rect -4338 671498 480 671734
rect -4756 671476 480 671498
rect 583520 672054 588680 672076
rect 583520 671818 588262 672054
rect 588498 671818 588680 672054
rect 583520 671734 588680 671818
rect 583520 671498 588262 671734
rect 588498 671498 588680 671734
rect 583520 671476 588680 671498
rect -4756 671474 -4156 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 586240 668476 586840 668478
rect -2916 668454 480 668476
rect -2916 668218 -2734 668454
rect -2498 668218 480 668454
rect -2916 668134 480 668218
rect -2916 667898 -2734 668134
rect -2498 667898 480 668134
rect -2916 667876 480 667898
rect 583520 668454 586840 668476
rect 583520 668218 586422 668454
rect 586658 668218 586840 668454
rect 583520 668134 586840 668218
rect 583520 667898 586422 668134
rect 586658 667898 586840 668134
rect 583520 667876 586840 667898
rect -2916 667874 -2316 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 590840 661276 591440 661278
rect -8436 661254 480 661276
rect -8436 661018 -7334 661254
rect -7098 661018 480 661254
rect -8436 660934 480 661018
rect -8436 660698 -7334 660934
rect -7098 660698 480 660934
rect -8436 660676 480 660698
rect 583520 661254 592360 661276
rect 583520 661018 591022 661254
rect 591258 661018 592360 661254
rect 583520 660934 592360 661018
rect 583520 660698 591022 660934
rect 591258 660698 592360 660934
rect 583520 660676 592360 660698
rect -7516 660674 -6916 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 589000 657676 589600 657678
rect -6596 657654 480 657676
rect -6596 657418 -5494 657654
rect -5258 657418 480 657654
rect -6596 657334 480 657418
rect -6596 657098 -5494 657334
rect -5258 657098 480 657334
rect -6596 657076 480 657098
rect 583520 657654 590520 657676
rect 583520 657418 589182 657654
rect 589418 657418 590520 657654
rect 583520 657334 590520 657418
rect 583520 657098 589182 657334
rect 589418 657098 590520 657334
rect 583520 657076 590520 657098
rect -5676 657074 -5076 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 587160 654076 587760 654078
rect -4756 654054 480 654076
rect -4756 653818 -3654 654054
rect -3418 653818 480 654054
rect -4756 653734 480 653818
rect -4756 653498 -3654 653734
rect -3418 653498 480 653734
rect -4756 653476 480 653498
rect 583520 654054 588680 654076
rect 583520 653818 587342 654054
rect 587578 653818 588680 654054
rect 583520 653734 588680 653818
rect 583520 653498 587342 653734
rect 587578 653498 588680 653734
rect 583520 653476 588680 653498
rect -3836 653474 -3236 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 585320 650476 585920 650478
rect -2916 650454 480 650476
rect -2916 650218 -1814 650454
rect -1578 650218 480 650454
rect -2916 650134 480 650218
rect -2916 649898 -1814 650134
rect -1578 649898 480 650134
rect -2916 649876 480 649898
rect 583520 650454 586840 650476
rect 583520 650218 585502 650454
rect 585738 650218 586840 650454
rect 583520 650134 586840 650218
rect 583520 649898 585502 650134
rect 585738 649898 586840 650134
rect 583520 649876 586840 649898
rect -1996 649874 -1396 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 591760 643276 592360 643278
rect -8436 643254 480 643276
rect -8436 643018 -8254 643254
rect -8018 643018 480 643254
rect -8436 642934 480 643018
rect -8436 642698 -8254 642934
rect -8018 642698 480 642934
rect -8436 642676 480 642698
rect 583520 643254 592360 643276
rect 583520 643018 591942 643254
rect 592178 643018 592360 643254
rect 583520 642934 592360 643018
rect 583520 642698 591942 642934
rect 592178 642698 592360 642934
rect 583520 642676 592360 642698
rect -8436 642674 -7836 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 589920 639676 590520 639678
rect -6596 639654 480 639676
rect -6596 639418 -6414 639654
rect -6178 639418 480 639654
rect -6596 639334 480 639418
rect -6596 639098 -6414 639334
rect -6178 639098 480 639334
rect -6596 639076 480 639098
rect 583520 639654 590520 639676
rect 583520 639418 590102 639654
rect 590338 639418 590520 639654
rect 583520 639334 590520 639418
rect 583520 639098 590102 639334
rect 590338 639098 590520 639334
rect 583520 639076 590520 639098
rect -6596 639074 -5996 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 588080 636076 588680 636078
rect -4756 636054 480 636076
rect -4756 635818 -4574 636054
rect -4338 635818 480 636054
rect -4756 635734 480 635818
rect -4756 635498 -4574 635734
rect -4338 635498 480 635734
rect -4756 635476 480 635498
rect 583520 636054 588680 636076
rect 583520 635818 588262 636054
rect 588498 635818 588680 636054
rect 583520 635734 588680 635818
rect 583520 635498 588262 635734
rect 588498 635498 588680 635734
rect 583520 635476 588680 635498
rect -4756 635474 -4156 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 586240 632476 586840 632478
rect -2916 632454 480 632476
rect -2916 632218 -2734 632454
rect -2498 632218 480 632454
rect -2916 632134 480 632218
rect -2916 631898 -2734 632134
rect -2498 631898 480 632134
rect -2916 631876 480 631898
rect 583520 632454 586840 632476
rect 583520 632218 586422 632454
rect 586658 632218 586840 632454
rect 583520 632134 586840 632218
rect 583520 631898 586422 632134
rect 586658 631898 586840 632134
rect 583520 631876 586840 631898
rect -2916 631874 -2316 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 590840 625276 591440 625278
rect -8436 625254 480 625276
rect -8436 625018 -7334 625254
rect -7098 625018 480 625254
rect -8436 624934 480 625018
rect -8436 624698 -7334 624934
rect -7098 624698 480 624934
rect -8436 624676 480 624698
rect 583520 625254 592360 625276
rect 583520 625018 591022 625254
rect 591258 625018 592360 625254
rect 583520 624934 592360 625018
rect 583520 624698 591022 624934
rect 591258 624698 592360 624934
rect 583520 624676 592360 624698
rect -7516 624674 -6916 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 589000 621676 589600 621678
rect -6596 621654 480 621676
rect -6596 621418 -5494 621654
rect -5258 621418 480 621654
rect -6596 621334 480 621418
rect -6596 621098 -5494 621334
rect -5258 621098 480 621334
rect -6596 621076 480 621098
rect 583520 621654 590520 621676
rect 583520 621418 589182 621654
rect 589418 621418 590520 621654
rect 583520 621334 590520 621418
rect 583520 621098 589182 621334
rect 589418 621098 590520 621334
rect 583520 621076 590520 621098
rect -5676 621074 -5076 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 587160 618076 587760 618078
rect -4756 618054 480 618076
rect -4756 617818 -3654 618054
rect -3418 617818 480 618054
rect -4756 617734 480 617818
rect -4756 617498 -3654 617734
rect -3418 617498 480 617734
rect -4756 617476 480 617498
rect 583520 618054 588680 618076
rect 583520 617818 587342 618054
rect 587578 617818 588680 618054
rect 583520 617734 588680 617818
rect 583520 617498 587342 617734
rect 587578 617498 588680 617734
rect 583520 617476 588680 617498
rect -3836 617474 -3236 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 585320 614476 585920 614478
rect -2916 614454 480 614476
rect -2916 614218 -1814 614454
rect -1578 614218 480 614454
rect -2916 614134 480 614218
rect -2916 613898 -1814 614134
rect -1578 613898 480 614134
rect -2916 613876 480 613898
rect 583520 614454 586840 614476
rect 583520 614218 585502 614454
rect 585738 614218 586840 614454
rect 583520 614134 586840 614218
rect 583520 613898 585502 614134
rect 585738 613898 586840 614134
rect 583520 613876 586840 613898
rect -1996 613874 -1396 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 591760 607276 592360 607278
rect -8436 607254 480 607276
rect -8436 607018 -8254 607254
rect -8018 607018 480 607254
rect -8436 606934 480 607018
rect -8436 606698 -8254 606934
rect -8018 606698 480 606934
rect -8436 606676 480 606698
rect 583520 607254 592360 607276
rect 583520 607018 591942 607254
rect 592178 607018 592360 607254
rect 583520 606934 592360 607018
rect 583520 606698 591942 606934
rect 592178 606698 592360 606934
rect 583520 606676 592360 606698
rect -8436 606674 -7836 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 589920 603676 590520 603678
rect -6596 603654 480 603676
rect -6596 603418 -6414 603654
rect -6178 603418 480 603654
rect -6596 603334 480 603418
rect -6596 603098 -6414 603334
rect -6178 603098 480 603334
rect -6596 603076 480 603098
rect 583520 603654 590520 603676
rect 583520 603418 590102 603654
rect 590338 603418 590520 603654
rect 583520 603334 590520 603418
rect 583520 603098 590102 603334
rect 590338 603098 590520 603334
rect 583520 603076 590520 603098
rect -6596 603074 -5996 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 588080 600076 588680 600078
rect -4756 600054 480 600076
rect -4756 599818 -4574 600054
rect -4338 599818 480 600054
rect -4756 599734 480 599818
rect -4756 599498 -4574 599734
rect -4338 599498 480 599734
rect -4756 599476 480 599498
rect 583520 600054 588680 600076
rect 583520 599818 588262 600054
rect 588498 599818 588680 600054
rect 583520 599734 588680 599818
rect 583520 599498 588262 599734
rect 588498 599498 588680 599734
rect 583520 599476 588680 599498
rect -4756 599474 -4156 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 586240 596476 586840 596478
rect -2916 596454 480 596476
rect -2916 596218 -2734 596454
rect -2498 596218 480 596454
rect -2916 596134 480 596218
rect -2916 595898 -2734 596134
rect -2498 595898 480 596134
rect -2916 595876 480 595898
rect 583520 596454 586840 596476
rect 583520 596218 586422 596454
rect 586658 596218 586840 596454
rect 583520 596134 586840 596218
rect 583520 595898 586422 596134
rect 586658 595898 586840 596134
rect 583520 595876 586840 595898
rect -2916 595874 -2316 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 590840 589276 591440 589278
rect -8436 589254 480 589276
rect -8436 589018 -7334 589254
rect -7098 589018 480 589254
rect -8436 588934 480 589018
rect -8436 588698 -7334 588934
rect -7098 588698 480 588934
rect -8436 588676 480 588698
rect 583520 589254 592360 589276
rect 583520 589018 591022 589254
rect 591258 589018 592360 589254
rect 583520 588934 592360 589018
rect 583520 588698 591022 588934
rect 591258 588698 592360 588934
rect 583520 588676 592360 588698
rect -7516 588674 -6916 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 589000 585676 589600 585678
rect -6596 585654 480 585676
rect -6596 585418 -5494 585654
rect -5258 585418 480 585654
rect -6596 585334 480 585418
rect -6596 585098 -5494 585334
rect -5258 585098 480 585334
rect -6596 585076 480 585098
rect 583520 585654 590520 585676
rect 583520 585418 589182 585654
rect 589418 585418 590520 585654
rect 583520 585334 590520 585418
rect 583520 585098 589182 585334
rect 589418 585098 590520 585334
rect 583520 585076 590520 585098
rect -5676 585074 -5076 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 587160 582076 587760 582078
rect -4756 582054 480 582076
rect -4756 581818 -3654 582054
rect -3418 581818 480 582054
rect -4756 581734 480 581818
rect -4756 581498 -3654 581734
rect -3418 581498 480 581734
rect -4756 581476 480 581498
rect 583520 582054 588680 582076
rect 583520 581818 587342 582054
rect 587578 581818 588680 582054
rect 583520 581734 588680 581818
rect 583520 581498 587342 581734
rect 587578 581498 588680 581734
rect 583520 581476 588680 581498
rect -3836 581474 -3236 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 585320 578476 585920 578478
rect -2916 578454 480 578476
rect -2916 578218 -1814 578454
rect -1578 578218 480 578454
rect -2916 578134 480 578218
rect -2916 577898 -1814 578134
rect -1578 577898 480 578134
rect -2916 577876 480 577898
rect 583520 578454 586840 578476
rect 583520 578218 585502 578454
rect 585738 578218 586840 578454
rect 583520 578134 586840 578218
rect 583520 577898 585502 578134
rect 585738 577898 586840 578134
rect 583520 577876 586840 577898
rect -1996 577874 -1396 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 591760 571276 592360 571278
rect -8436 571254 480 571276
rect -8436 571018 -8254 571254
rect -8018 571018 480 571254
rect -8436 570934 480 571018
rect -8436 570698 -8254 570934
rect -8018 570698 480 570934
rect -8436 570676 480 570698
rect 583520 571254 592360 571276
rect 583520 571018 591942 571254
rect 592178 571018 592360 571254
rect 583520 570934 592360 571018
rect 583520 570698 591942 570934
rect 592178 570698 592360 570934
rect 583520 570676 592360 570698
rect -8436 570674 -7836 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 589920 567676 590520 567678
rect -6596 567654 480 567676
rect -6596 567418 -6414 567654
rect -6178 567418 480 567654
rect -6596 567334 480 567418
rect -6596 567098 -6414 567334
rect -6178 567098 480 567334
rect -6596 567076 480 567098
rect 583520 567654 590520 567676
rect 583520 567418 590102 567654
rect 590338 567418 590520 567654
rect 583520 567334 590520 567418
rect 583520 567098 590102 567334
rect 590338 567098 590520 567334
rect 583520 567076 590520 567098
rect -6596 567074 -5996 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 588080 564076 588680 564078
rect -4756 564054 480 564076
rect -4756 563818 -4574 564054
rect -4338 563818 480 564054
rect -4756 563734 480 563818
rect -4756 563498 -4574 563734
rect -4338 563498 480 563734
rect -4756 563476 480 563498
rect 583520 564054 588680 564076
rect 583520 563818 588262 564054
rect 588498 563818 588680 564054
rect 583520 563734 588680 563818
rect 583520 563498 588262 563734
rect 588498 563498 588680 563734
rect 583520 563476 588680 563498
rect -4756 563474 -4156 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 586240 560476 586840 560478
rect -2916 560454 480 560476
rect -2916 560218 -2734 560454
rect -2498 560218 480 560454
rect -2916 560134 480 560218
rect -2916 559898 -2734 560134
rect -2498 559898 480 560134
rect -2916 559876 480 559898
rect 583520 560454 586840 560476
rect 583520 560218 586422 560454
rect 586658 560218 586840 560454
rect 583520 560134 586840 560218
rect 583520 559898 586422 560134
rect 586658 559898 586840 560134
rect 583520 559876 586840 559898
rect -2916 559874 -2316 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 590840 553276 591440 553278
rect -8436 553254 480 553276
rect -8436 553018 -7334 553254
rect -7098 553018 480 553254
rect -8436 552934 480 553018
rect -8436 552698 -7334 552934
rect -7098 552698 480 552934
rect -8436 552676 480 552698
rect 583520 553254 592360 553276
rect 583520 553018 591022 553254
rect 591258 553018 592360 553254
rect 583520 552934 592360 553018
rect 583520 552698 591022 552934
rect 591258 552698 592360 552934
rect 583520 552676 592360 552698
rect -7516 552674 -6916 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 589000 549676 589600 549678
rect -6596 549654 480 549676
rect -6596 549418 -5494 549654
rect -5258 549418 480 549654
rect -6596 549334 480 549418
rect -6596 549098 -5494 549334
rect -5258 549098 480 549334
rect -6596 549076 480 549098
rect 583520 549654 590520 549676
rect 583520 549418 589182 549654
rect 589418 549418 590520 549654
rect 583520 549334 590520 549418
rect 583520 549098 589182 549334
rect 589418 549098 590520 549334
rect 583520 549076 590520 549098
rect -5676 549074 -5076 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 587160 546076 587760 546078
rect -4756 546054 480 546076
rect -4756 545818 -3654 546054
rect -3418 545818 480 546054
rect -4756 545734 480 545818
rect -4756 545498 -3654 545734
rect -3418 545498 480 545734
rect -4756 545476 480 545498
rect 583520 546054 588680 546076
rect 583520 545818 587342 546054
rect 587578 545818 588680 546054
rect 583520 545734 588680 545818
rect 583520 545498 587342 545734
rect 587578 545498 588680 545734
rect 583520 545476 588680 545498
rect -3836 545474 -3236 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 585320 542476 585920 542478
rect -2916 542454 480 542476
rect -2916 542218 -1814 542454
rect -1578 542218 480 542454
rect -2916 542134 480 542218
rect -2916 541898 -1814 542134
rect -1578 541898 480 542134
rect -2916 541876 480 541898
rect 583520 542454 586840 542476
rect 583520 542218 585502 542454
rect 585738 542218 586840 542454
rect 583520 542134 586840 542218
rect 583520 541898 585502 542134
rect 585738 541898 586840 542134
rect 583520 541876 586840 541898
rect -1996 541874 -1396 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 591760 535276 592360 535278
rect -8436 535254 480 535276
rect -8436 535018 -8254 535254
rect -8018 535018 480 535254
rect -8436 534934 480 535018
rect -8436 534698 -8254 534934
rect -8018 534698 480 534934
rect -8436 534676 480 534698
rect 583520 535254 592360 535276
rect 583520 535018 591942 535254
rect 592178 535018 592360 535254
rect 583520 534934 592360 535018
rect 583520 534698 591942 534934
rect 592178 534698 592360 534934
rect 583520 534676 592360 534698
rect -8436 534674 -7836 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 589920 531676 590520 531678
rect -6596 531654 480 531676
rect -6596 531418 -6414 531654
rect -6178 531418 480 531654
rect -6596 531334 480 531418
rect -6596 531098 -6414 531334
rect -6178 531098 480 531334
rect -6596 531076 480 531098
rect 583520 531654 590520 531676
rect 583520 531418 590102 531654
rect 590338 531418 590520 531654
rect 583520 531334 590520 531418
rect 583520 531098 590102 531334
rect 590338 531098 590520 531334
rect 583520 531076 590520 531098
rect -6596 531074 -5996 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 588080 528076 588680 528078
rect -4756 528054 480 528076
rect -4756 527818 -4574 528054
rect -4338 527818 480 528054
rect -4756 527734 480 527818
rect -4756 527498 -4574 527734
rect -4338 527498 480 527734
rect -4756 527476 480 527498
rect 583520 528054 588680 528076
rect 583520 527818 588262 528054
rect 588498 527818 588680 528054
rect 583520 527734 588680 527818
rect 583520 527498 588262 527734
rect 588498 527498 588680 527734
rect 583520 527476 588680 527498
rect -4756 527474 -4156 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 586240 524476 586840 524478
rect -2916 524454 480 524476
rect -2916 524218 -2734 524454
rect -2498 524218 480 524454
rect -2916 524134 480 524218
rect -2916 523898 -2734 524134
rect -2498 523898 480 524134
rect -2916 523876 480 523898
rect 583520 524454 586840 524476
rect 583520 524218 586422 524454
rect 586658 524218 586840 524454
rect 583520 524134 586840 524218
rect 583520 523898 586422 524134
rect 586658 523898 586840 524134
rect 583520 523876 586840 523898
rect -2916 523874 -2316 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 590840 517276 591440 517278
rect -8436 517254 480 517276
rect -8436 517018 -7334 517254
rect -7098 517018 480 517254
rect -8436 516934 480 517018
rect -8436 516698 -7334 516934
rect -7098 516698 480 516934
rect -8436 516676 480 516698
rect 583520 517254 592360 517276
rect 583520 517018 591022 517254
rect 591258 517018 592360 517254
rect 583520 516934 592360 517018
rect 583520 516698 591022 516934
rect 591258 516698 592360 516934
rect 583520 516676 592360 516698
rect -7516 516674 -6916 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 589000 513676 589600 513678
rect -6596 513654 480 513676
rect -6596 513418 -5494 513654
rect -5258 513418 480 513654
rect -6596 513334 480 513418
rect -6596 513098 -5494 513334
rect -5258 513098 480 513334
rect -6596 513076 480 513098
rect 583520 513654 590520 513676
rect 583520 513418 589182 513654
rect 589418 513418 590520 513654
rect 583520 513334 590520 513418
rect 583520 513098 589182 513334
rect 589418 513098 590520 513334
rect 583520 513076 590520 513098
rect -5676 513074 -5076 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 587160 510076 587760 510078
rect -4756 510054 480 510076
rect -4756 509818 -3654 510054
rect -3418 509818 480 510054
rect -4756 509734 480 509818
rect -4756 509498 -3654 509734
rect -3418 509498 480 509734
rect -4756 509476 480 509498
rect 583520 510054 588680 510076
rect 583520 509818 587342 510054
rect 587578 509818 588680 510054
rect 583520 509734 588680 509818
rect 583520 509498 587342 509734
rect 587578 509498 588680 509734
rect 583520 509476 588680 509498
rect -3836 509474 -3236 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 585320 506476 585920 506478
rect -2916 506454 480 506476
rect -2916 506218 -1814 506454
rect -1578 506218 480 506454
rect -2916 506134 480 506218
rect -2916 505898 -1814 506134
rect -1578 505898 480 506134
rect -2916 505876 480 505898
rect 583520 506454 586840 506476
rect 583520 506218 585502 506454
rect 585738 506218 586840 506454
rect 583520 506134 586840 506218
rect 583520 505898 585502 506134
rect 585738 505898 586840 506134
rect 583520 505876 586840 505898
rect -1996 505874 -1396 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 591760 499276 592360 499278
rect -8436 499254 480 499276
rect -8436 499018 -8254 499254
rect -8018 499018 480 499254
rect -8436 498934 480 499018
rect -8436 498698 -8254 498934
rect -8018 498698 480 498934
rect -8436 498676 480 498698
rect 583520 499254 592360 499276
rect 583520 499018 591942 499254
rect 592178 499018 592360 499254
rect 583520 498934 592360 499018
rect 583520 498698 591942 498934
rect 592178 498698 592360 498934
rect 583520 498676 592360 498698
rect -8436 498674 -7836 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 589920 495676 590520 495678
rect -6596 495654 480 495676
rect -6596 495418 -6414 495654
rect -6178 495418 480 495654
rect -6596 495334 480 495418
rect -6596 495098 -6414 495334
rect -6178 495098 480 495334
rect -6596 495076 480 495098
rect 583520 495654 590520 495676
rect 583520 495418 590102 495654
rect 590338 495418 590520 495654
rect 583520 495334 590520 495418
rect 583520 495098 590102 495334
rect 590338 495098 590520 495334
rect 583520 495076 590520 495098
rect -6596 495074 -5996 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 588080 492076 588680 492078
rect -4756 492054 480 492076
rect -4756 491818 -4574 492054
rect -4338 491818 480 492054
rect -4756 491734 480 491818
rect -4756 491498 -4574 491734
rect -4338 491498 480 491734
rect -4756 491476 480 491498
rect 583520 492054 588680 492076
rect 583520 491818 588262 492054
rect 588498 491818 588680 492054
rect 583520 491734 588680 491818
rect 583520 491498 588262 491734
rect 588498 491498 588680 491734
rect 583520 491476 588680 491498
rect -4756 491474 -4156 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 586240 488476 586840 488478
rect -2916 488454 480 488476
rect -2916 488218 -2734 488454
rect -2498 488218 480 488454
rect -2916 488134 480 488218
rect -2916 487898 -2734 488134
rect -2498 487898 480 488134
rect -2916 487876 480 487898
rect 583520 488454 586840 488476
rect 583520 488218 586422 488454
rect 586658 488218 586840 488454
rect 583520 488134 586840 488218
rect 583520 487898 586422 488134
rect 586658 487898 586840 488134
rect 583520 487876 586840 487898
rect -2916 487874 -2316 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 590840 481276 591440 481278
rect -8436 481254 480 481276
rect -8436 481018 -7334 481254
rect -7098 481018 480 481254
rect -8436 480934 480 481018
rect -8436 480698 -7334 480934
rect -7098 480698 480 480934
rect -8436 480676 480 480698
rect 583520 481254 592360 481276
rect 583520 481018 591022 481254
rect 591258 481018 592360 481254
rect 583520 480934 592360 481018
rect 583520 480698 591022 480934
rect 591258 480698 592360 480934
rect 583520 480676 592360 480698
rect -7516 480674 -6916 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 589000 477676 589600 477678
rect -6596 477654 480 477676
rect -6596 477418 -5494 477654
rect -5258 477418 480 477654
rect -6596 477334 480 477418
rect -6596 477098 -5494 477334
rect -5258 477098 480 477334
rect -6596 477076 480 477098
rect 583520 477654 590520 477676
rect 583520 477418 589182 477654
rect 589418 477418 590520 477654
rect 583520 477334 590520 477418
rect 583520 477098 589182 477334
rect 589418 477098 590520 477334
rect 583520 477076 590520 477098
rect -5676 477074 -5076 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 587160 474076 587760 474078
rect -4756 474054 480 474076
rect -4756 473818 -3654 474054
rect -3418 473818 480 474054
rect -4756 473734 480 473818
rect -4756 473498 -3654 473734
rect -3418 473498 480 473734
rect -4756 473476 480 473498
rect 583520 474054 588680 474076
rect 583520 473818 587342 474054
rect 587578 473818 588680 474054
rect 583520 473734 588680 473818
rect 583520 473498 587342 473734
rect 587578 473498 588680 473734
rect 583520 473476 588680 473498
rect -3836 473474 -3236 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 585320 470476 585920 470478
rect -2916 470454 480 470476
rect -2916 470218 -1814 470454
rect -1578 470218 480 470454
rect -2916 470134 480 470218
rect -2916 469898 -1814 470134
rect -1578 469898 480 470134
rect -2916 469876 480 469898
rect 583520 470454 586840 470476
rect 583520 470218 585502 470454
rect 585738 470218 586840 470454
rect 583520 470134 586840 470218
rect 583520 469898 585502 470134
rect 585738 469898 586840 470134
rect 583520 469876 586840 469898
rect -1996 469874 -1396 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 591760 463276 592360 463278
rect -8436 463254 480 463276
rect -8436 463018 -8254 463254
rect -8018 463018 480 463254
rect -8436 462934 480 463018
rect -8436 462698 -8254 462934
rect -8018 462698 480 462934
rect -8436 462676 480 462698
rect 583520 463254 592360 463276
rect 583520 463018 591942 463254
rect 592178 463018 592360 463254
rect 583520 462934 592360 463018
rect 583520 462698 591942 462934
rect 592178 462698 592360 462934
rect 583520 462676 592360 462698
rect -8436 462674 -7836 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 589920 459676 590520 459678
rect -6596 459654 480 459676
rect -6596 459418 -6414 459654
rect -6178 459418 480 459654
rect -6596 459334 480 459418
rect -6596 459098 -6414 459334
rect -6178 459098 480 459334
rect -6596 459076 480 459098
rect 583520 459654 590520 459676
rect 583520 459418 590102 459654
rect 590338 459418 590520 459654
rect 583520 459334 590520 459418
rect 583520 459098 590102 459334
rect 590338 459098 590520 459334
rect 583520 459076 590520 459098
rect -6596 459074 -5996 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 588080 456076 588680 456078
rect -4756 456054 480 456076
rect -4756 455818 -4574 456054
rect -4338 455818 480 456054
rect -4756 455734 480 455818
rect -4756 455498 -4574 455734
rect -4338 455498 480 455734
rect -4756 455476 480 455498
rect 583520 456054 588680 456076
rect 583520 455818 588262 456054
rect 588498 455818 588680 456054
rect 583520 455734 588680 455818
rect 583520 455498 588262 455734
rect 588498 455498 588680 455734
rect 583520 455476 588680 455498
rect -4756 455474 -4156 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 586240 452476 586840 452478
rect -2916 452454 480 452476
rect -2916 452218 -2734 452454
rect -2498 452218 480 452454
rect -2916 452134 480 452218
rect -2916 451898 -2734 452134
rect -2498 451898 480 452134
rect -2916 451876 480 451898
rect 583520 452454 586840 452476
rect 583520 452218 586422 452454
rect 586658 452218 586840 452454
rect 583520 452134 586840 452218
rect 583520 451898 586422 452134
rect 586658 451898 586840 452134
rect 583520 451876 586840 451898
rect -2916 451874 -2316 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 590840 445276 591440 445278
rect -8436 445254 480 445276
rect -8436 445018 -7334 445254
rect -7098 445018 480 445254
rect -8436 444934 480 445018
rect -8436 444698 -7334 444934
rect -7098 444698 480 444934
rect -8436 444676 480 444698
rect 583520 445254 592360 445276
rect 583520 445018 591022 445254
rect 591258 445018 592360 445254
rect 583520 444934 592360 445018
rect 583520 444698 591022 444934
rect 591258 444698 592360 444934
rect 583520 444676 592360 444698
rect -7516 444674 -6916 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 589000 441676 589600 441678
rect -6596 441654 480 441676
rect -6596 441418 -5494 441654
rect -5258 441418 480 441654
rect -6596 441334 480 441418
rect -6596 441098 -5494 441334
rect -5258 441098 480 441334
rect -6596 441076 480 441098
rect 583520 441654 590520 441676
rect 583520 441418 589182 441654
rect 589418 441418 590520 441654
rect 583520 441334 590520 441418
rect 583520 441098 589182 441334
rect 589418 441098 590520 441334
rect 583520 441076 590520 441098
rect -5676 441074 -5076 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 587160 438076 587760 438078
rect -4756 438054 480 438076
rect -4756 437818 -3654 438054
rect -3418 437818 480 438054
rect -4756 437734 480 437818
rect -4756 437498 -3654 437734
rect -3418 437498 480 437734
rect -4756 437476 480 437498
rect 583520 438054 588680 438076
rect 583520 437818 587342 438054
rect 587578 437818 588680 438054
rect 583520 437734 588680 437818
rect 583520 437498 587342 437734
rect 587578 437498 588680 437734
rect 583520 437476 588680 437498
rect -3836 437474 -3236 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 585320 434476 585920 434478
rect -2916 434454 480 434476
rect -2916 434218 -1814 434454
rect -1578 434218 480 434454
rect -2916 434134 480 434218
rect -2916 433898 -1814 434134
rect -1578 433898 480 434134
rect -2916 433876 480 433898
rect 583520 434454 586840 434476
rect 583520 434218 585502 434454
rect 585738 434218 586840 434454
rect 583520 434134 586840 434218
rect 583520 433898 585502 434134
rect 585738 433898 586840 434134
rect 583520 433876 586840 433898
rect -1996 433874 -1396 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 591760 427276 592360 427278
rect -8436 427254 480 427276
rect -8436 427018 -8254 427254
rect -8018 427018 480 427254
rect -8436 426934 480 427018
rect -8436 426698 -8254 426934
rect -8018 426698 480 426934
rect -8436 426676 480 426698
rect 583520 427254 592360 427276
rect 583520 427018 591942 427254
rect 592178 427018 592360 427254
rect 583520 426934 592360 427018
rect 583520 426698 591942 426934
rect 592178 426698 592360 426934
rect 583520 426676 592360 426698
rect -8436 426674 -7836 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 589920 423676 590520 423678
rect -6596 423654 480 423676
rect -6596 423418 -6414 423654
rect -6178 423418 480 423654
rect -6596 423334 480 423418
rect -6596 423098 -6414 423334
rect -6178 423098 480 423334
rect -6596 423076 480 423098
rect 583520 423654 590520 423676
rect 583520 423418 590102 423654
rect 590338 423418 590520 423654
rect 583520 423334 590520 423418
rect 583520 423098 590102 423334
rect 590338 423098 590520 423334
rect 583520 423076 590520 423098
rect -6596 423074 -5996 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 588080 420076 588680 420078
rect -4756 420054 480 420076
rect -4756 419818 -4574 420054
rect -4338 419818 480 420054
rect -4756 419734 480 419818
rect -4756 419498 -4574 419734
rect -4338 419498 480 419734
rect -4756 419476 480 419498
rect 583520 420054 588680 420076
rect 583520 419818 588262 420054
rect 588498 419818 588680 420054
rect 583520 419734 588680 419818
rect 583520 419498 588262 419734
rect 588498 419498 588680 419734
rect 583520 419476 588680 419498
rect -4756 419474 -4156 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 586240 416476 586840 416478
rect -2916 416454 480 416476
rect -2916 416218 -2734 416454
rect -2498 416218 480 416454
rect -2916 416134 480 416218
rect -2916 415898 -2734 416134
rect -2498 415898 480 416134
rect -2916 415876 480 415898
rect 582212 416454 586840 416476
rect 582212 416218 586422 416454
rect 586658 416218 586840 416454
rect 582212 416134 586840 416218
rect 582212 415898 586422 416134
rect 586658 415898 586840 416134
rect 582212 415876 586840 415898
rect -2916 415874 -2316 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 590840 409276 591440 409278
rect -8436 409254 480 409276
rect -8436 409018 -7334 409254
rect -7098 409018 480 409254
rect -8436 408934 480 409018
rect -8436 408698 -7334 408934
rect -7098 408698 480 408934
rect -8436 408676 480 408698
rect 583520 409254 592360 409276
rect 583520 409018 591022 409254
rect 591258 409018 592360 409254
rect 583520 408934 592360 409018
rect 583520 408698 591022 408934
rect 591258 408698 592360 408934
rect 583520 408676 592360 408698
rect -7516 408674 -6916 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 589000 405676 589600 405678
rect -6596 405654 480 405676
rect -6596 405418 -5494 405654
rect -5258 405418 480 405654
rect -6596 405334 480 405418
rect -6596 405098 -5494 405334
rect -5258 405098 480 405334
rect -6596 405076 480 405098
rect 583520 405654 590520 405676
rect 583520 405418 589182 405654
rect 589418 405418 590520 405654
rect 583520 405334 590520 405418
rect 583520 405098 589182 405334
rect 589418 405098 590520 405334
rect 583520 405076 590520 405098
rect -5676 405074 -5076 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 587160 402076 587760 402078
rect -4756 402054 480 402076
rect -4756 401818 -3654 402054
rect -3418 401818 480 402054
rect -4756 401734 480 401818
rect -4756 401498 -3654 401734
rect -3418 401498 480 401734
rect -4756 401476 480 401498
rect 582598 402054 588680 402076
rect 582598 401818 587342 402054
rect 587578 401818 588680 402054
rect 582598 401734 588680 401818
rect 582598 401498 587342 401734
rect 587578 401498 588680 401734
rect 582598 401476 588680 401498
rect -3836 401474 -3236 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 585320 398476 585920 398478
rect -2916 398454 480 398476
rect -2916 398218 -1814 398454
rect -1578 398218 480 398454
rect -2916 398134 480 398218
rect -2916 397898 -1814 398134
rect -1578 397898 480 398134
rect -2916 397876 480 397898
rect 583520 398454 586840 398476
rect 583520 398218 585502 398454
rect 585738 398218 586840 398454
rect 583520 398134 586840 398218
rect 583520 397898 585502 398134
rect 585738 397898 586840 398134
rect 583520 397876 586840 397898
rect -1996 397874 -1396 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 591760 391276 592360 391278
rect -8436 391254 480 391276
rect -8436 391018 -8254 391254
rect -8018 391018 480 391254
rect -8436 390934 480 391018
rect -8436 390698 -8254 390934
rect -8018 390698 480 390934
rect -8436 390676 480 390698
rect 583520 391254 592360 391276
rect 583520 391018 591942 391254
rect 592178 391018 592360 391254
rect 583520 390934 592360 391018
rect 583520 390698 591942 390934
rect 592178 390698 592360 390934
rect 583520 390676 592360 390698
rect -8436 390674 -7836 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 589920 387676 590520 387678
rect -6596 387654 480 387676
rect -6596 387418 -6414 387654
rect -6178 387418 480 387654
rect -6596 387334 480 387418
rect -6596 387098 -6414 387334
rect -6178 387098 480 387334
rect -6596 387076 480 387098
rect 583520 387654 590520 387676
rect 583520 387418 590102 387654
rect 590338 387418 590520 387654
rect 583520 387334 590520 387418
rect 583520 387098 590102 387334
rect 590338 387098 590520 387334
rect 583520 387076 590520 387098
rect -6596 387074 -5996 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 588080 384076 588680 384078
rect -4756 384054 480 384076
rect -4756 383818 -4574 384054
rect -4338 383818 480 384054
rect -4756 383734 480 383818
rect -4756 383498 -4574 383734
rect -4338 383498 480 383734
rect -4756 383476 480 383498
rect 583036 384054 588680 384076
rect 583036 383818 588262 384054
rect 588498 383818 588680 384054
rect 583036 383734 588680 383818
rect 583036 383498 588262 383734
rect 588498 383498 588680 383734
rect 583036 383476 588680 383498
rect -4756 383474 -4156 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 586240 380476 586840 380478
rect -2916 380454 480 380476
rect -2916 380218 -2734 380454
rect -2498 380218 480 380454
rect -2916 380134 480 380218
rect -2916 379898 -2734 380134
rect -2498 379898 480 380134
rect -2916 379876 480 379898
rect 582542 380454 586840 380476
rect 582542 380218 586422 380454
rect 586658 380218 586840 380454
rect 582542 380134 586840 380218
rect 582542 379898 586422 380134
rect 586658 379898 586840 380134
rect 582542 379876 586840 379898
rect -2916 379874 -2316 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 590840 373276 591440 373278
rect -8436 373254 480 373276
rect -8436 373018 -7334 373254
rect -7098 373018 480 373254
rect -8436 372934 480 373018
rect -8436 372698 -7334 372934
rect -7098 372698 480 372934
rect -8436 372676 480 372698
rect 583520 373254 592360 373276
rect 583520 373018 591022 373254
rect 591258 373018 592360 373254
rect 583520 372934 592360 373018
rect 583520 372698 591022 372934
rect 591258 372698 592360 372934
rect 583520 372676 592360 372698
rect -7516 372674 -6916 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 589000 369676 589600 369678
rect -6596 369654 480 369676
rect -6596 369418 -5494 369654
rect -5258 369418 480 369654
rect -6596 369334 480 369418
rect -6596 369098 -5494 369334
rect -5258 369098 480 369334
rect -6596 369076 480 369098
rect 583520 369654 590520 369676
rect 583520 369418 589182 369654
rect 589418 369418 590520 369654
rect 583520 369334 590520 369418
rect 583520 369098 589182 369334
rect 589418 369098 590520 369334
rect 583520 369076 590520 369098
rect -5676 369074 -5076 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 587160 366076 587760 366078
rect -4756 366054 480 366076
rect -4756 365818 -3654 366054
rect -3418 365818 480 366054
rect -4756 365734 480 365818
rect -4756 365498 -3654 365734
rect -3418 365498 480 365734
rect -4756 365476 480 365498
rect 583520 366054 588680 366076
rect 583520 365818 587342 366054
rect 587578 365818 588680 366054
rect 583520 365734 588680 365818
rect 583520 365498 587342 365734
rect 587578 365498 588680 365734
rect 583520 365476 588680 365498
rect -3836 365474 -3236 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 585320 362476 585920 362478
rect -2916 362454 480 362476
rect -2916 362218 -1814 362454
rect -1578 362218 480 362454
rect -2916 362134 480 362218
rect -2916 361898 -1814 362134
rect -1578 361898 480 362134
rect -2916 361876 480 361898
rect 583520 362454 586840 362476
rect 583520 362218 585502 362454
rect 585738 362218 586840 362454
rect 583520 362134 586840 362218
rect 583520 361898 585502 362134
rect 585738 361898 586840 362134
rect 583520 361876 586840 361898
rect -1996 361874 -1396 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 591760 355276 592360 355278
rect -8436 355254 480 355276
rect -8436 355018 -8254 355254
rect -8018 355018 480 355254
rect -8436 354934 480 355018
rect -8436 354698 -8254 354934
rect -8018 354698 480 354934
rect -8436 354676 480 354698
rect 583520 355254 592360 355276
rect 583520 355018 591942 355254
rect 592178 355018 592360 355254
rect 583520 354934 592360 355018
rect 583520 354698 591942 354934
rect 592178 354698 592360 354934
rect 583520 354676 592360 354698
rect -8436 354674 -7836 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 589920 351676 590520 351678
rect -6596 351654 480 351676
rect -6596 351418 -6414 351654
rect -6178 351418 480 351654
rect -6596 351334 480 351418
rect -6596 351098 -6414 351334
rect -6178 351098 480 351334
rect -6596 351076 480 351098
rect 583520 351654 590520 351676
rect 583520 351418 590102 351654
rect 590338 351418 590520 351654
rect 583520 351334 590520 351418
rect 583520 351098 590102 351334
rect 590338 351098 590520 351334
rect 583520 351076 590520 351098
rect -6596 351074 -5996 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 588080 348076 588680 348078
rect -4756 348054 480 348076
rect -4756 347818 -4574 348054
rect -4338 347818 480 348054
rect -4756 347734 480 347818
rect -4756 347498 -4574 347734
rect -4338 347498 480 347734
rect -4756 347476 480 347498
rect 583520 348054 588680 348076
rect 583520 347818 588262 348054
rect 588498 347818 588680 348054
rect 583520 347734 588680 347818
rect 583520 347498 588262 347734
rect 588498 347498 588680 347734
rect 583520 347476 588680 347498
rect -4756 347474 -4156 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 586240 344476 586840 344478
rect -2916 344454 480 344476
rect -2916 344218 -2734 344454
rect -2498 344218 480 344454
rect -2916 344134 480 344218
rect -2916 343898 -2734 344134
rect -2498 343898 480 344134
rect -2916 343876 480 343898
rect 583520 344454 586840 344476
rect 583520 344218 586422 344454
rect 586658 344218 586840 344454
rect 583520 344134 586840 344218
rect 583520 343898 586422 344134
rect 586658 343898 586840 344134
rect 583520 343876 586840 343898
rect -2916 343874 -2316 343876
rect 586240 343874 586840 343876
rect 352832 343742 353200 343766
rect 352832 343422 352856 343742
rect 353176 343422 353200 343742
rect 352832 343398 353200 343422
rect -7516 337276 -6916 337278
rect 352856 337276 353176 343398
rect 590840 337276 591440 337278
rect -8436 337254 480 337276
rect -8436 337018 -7334 337254
rect -7098 337018 480 337254
rect -8436 336934 480 337018
rect -8436 336698 -7334 336934
rect -7098 336698 480 336934
rect -8436 336676 480 336698
rect 351420 337254 592360 337276
rect 351420 337018 591022 337254
rect 591258 337018 592360 337254
rect 351420 336934 592360 337018
rect 351420 336698 591022 336934
rect 591258 336698 592360 336934
rect 351420 336676 592360 336698
rect -7516 336674 -6916 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 589000 333676 589600 333678
rect -6596 333654 480 333676
rect -6596 333418 -5494 333654
rect -5258 333418 480 333654
rect -6596 333334 480 333418
rect -6596 333098 -5494 333334
rect -5258 333098 480 333334
rect -6596 333076 480 333098
rect 583520 333654 590520 333676
rect 583520 333418 589182 333654
rect 589418 333418 590520 333654
rect 583520 333334 590520 333418
rect 583520 333098 589182 333334
rect 589418 333098 590520 333334
rect 583520 333076 590520 333098
rect -5676 333074 -5076 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 587160 330076 587760 330078
rect -4756 330054 480 330076
rect -4756 329818 -3654 330054
rect -3418 329818 480 330054
rect -4756 329734 480 329818
rect -4756 329498 -3654 329734
rect -3418 329498 480 329734
rect -4756 329476 480 329498
rect 583520 330054 588680 330076
rect 583520 329818 587342 330054
rect 587578 329818 588680 330054
rect 583520 329734 588680 329818
rect 583520 329498 587342 329734
rect 587578 329498 588680 329734
rect 583520 329476 588680 329498
rect -3836 329474 -3236 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 585320 326476 585920 326478
rect -2916 326454 480 326476
rect -2916 326218 -1814 326454
rect -1578 326218 480 326454
rect -2916 326134 480 326218
rect -2916 325898 -1814 326134
rect -1578 325898 480 326134
rect -2916 325876 480 325898
rect 583520 326454 586840 326476
rect 583520 326218 585502 326454
rect 585738 326218 586840 326454
rect 583520 326134 586840 326218
rect 583520 325898 585502 326134
rect 585738 325898 586840 326134
rect 583520 325876 586840 325898
rect -1996 325874 -1396 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 591760 319276 592360 319278
rect -8436 319254 480 319276
rect -8436 319018 -8254 319254
rect -8018 319018 480 319254
rect -8436 318934 480 319018
rect -8436 318698 -8254 318934
rect -8018 318698 480 318934
rect -8436 318676 480 318698
rect 583520 319254 592360 319276
rect 583520 319018 591942 319254
rect 592178 319018 592360 319254
rect 583520 318934 592360 319018
rect 583520 318698 591942 318934
rect 592178 318698 592360 318934
rect 583520 318676 592360 318698
rect -8436 318674 -7836 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 589920 315676 590520 315678
rect -6596 315654 480 315676
rect -6596 315418 -6414 315654
rect -6178 315418 480 315654
rect -6596 315334 480 315418
rect -6596 315098 -6414 315334
rect -6178 315098 480 315334
rect -6596 315076 480 315098
rect 583520 315654 590520 315676
rect 583520 315418 590102 315654
rect 590338 315418 590520 315654
rect 583520 315334 590520 315418
rect 583520 315098 590102 315334
rect 590338 315098 590520 315334
rect 583520 315076 590520 315098
rect -6596 315074 -5996 315076
rect 589920 315074 590520 315076
rect 338134 312212 338502 312236
rect -4756 312076 -4156 312078
rect -4756 312054 480 312076
rect -4756 311818 -4574 312054
rect -4338 311818 480 312054
rect 338134 311892 338158 312212
rect 338478 311892 338502 312212
rect 588080 312076 588680 312078
rect 338134 311868 338502 311892
rect 583520 312054 588680 312076
rect -4756 311734 480 311818
rect -4756 311498 -4574 311734
rect -4338 311498 480 311734
rect -4756 311476 480 311498
rect -4756 311474 -4156 311476
rect -2916 308476 -2316 308478
rect -2916 308454 480 308476
rect -2916 308218 -2734 308454
rect -2498 308218 480 308454
rect -2916 308134 480 308218
rect -2916 307898 -2734 308134
rect -2498 307898 480 308134
rect -2916 307876 480 307898
rect -2916 307874 -2316 307876
rect -7516 301276 -6916 301278
rect -8436 301254 480 301276
rect -8436 301018 -7334 301254
rect -7098 301018 480 301254
rect -8436 300934 480 301018
rect -8436 300698 -7334 300934
rect -7098 300698 480 300934
rect -8436 300676 480 300698
rect -7516 300674 -6916 300676
rect -5676 297676 -5076 297678
rect 338158 297676 338478 311868
rect 583520 311818 588262 312054
rect 588498 311818 588680 312054
rect 583520 311734 588680 311818
rect 583520 311498 588262 311734
rect 588498 311498 588680 311734
rect 583520 311476 588680 311498
rect 588080 311474 588680 311476
rect 586240 308476 586840 308478
rect 583520 308454 586840 308476
rect 583520 308218 586422 308454
rect 586658 308218 586840 308454
rect 583520 308134 586840 308218
rect 583520 307898 586422 308134
rect 586658 307898 586840 308134
rect 583520 307876 586840 307898
rect 586240 307874 586840 307876
rect 590840 301276 591440 301278
rect 583290 301254 592360 301276
rect 583290 301018 591022 301254
rect 591258 301018 592360 301254
rect 583290 300934 592360 301018
rect 583290 300698 591022 300934
rect 591258 300698 592360 300934
rect 583290 300676 592360 300698
rect 590840 300674 591440 300676
rect 589000 297676 589600 297678
rect -6596 297654 480 297676
rect -6596 297418 -5494 297654
rect -5258 297418 480 297654
rect -6596 297334 480 297418
rect -6596 297098 -5494 297334
rect -5258 297098 480 297334
rect -6596 297076 480 297098
rect 336214 297654 590520 297676
rect 336214 297418 589182 297654
rect 589418 297418 590520 297654
rect 336214 297334 590520 297418
rect 336214 297098 589182 297334
rect 589418 297098 590520 297334
rect 336214 297076 590520 297098
rect -5676 297074 -5076 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 587160 294076 587760 294078
rect -4756 294054 480 294076
rect -4756 293818 -3654 294054
rect -3418 293818 480 294054
rect -4756 293734 480 293818
rect -4756 293498 -3654 293734
rect -3418 293498 480 293734
rect -4756 293476 480 293498
rect 583520 294054 588680 294076
rect 583520 293818 587342 294054
rect 587578 293818 588680 294054
rect 583520 293734 588680 293818
rect 583520 293498 587342 293734
rect 587578 293498 588680 293734
rect 583520 293476 588680 293498
rect -3836 293474 -3236 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 585320 290476 585920 290478
rect -2916 290454 480 290476
rect -2916 290218 -1814 290454
rect -1578 290218 480 290454
rect -2916 290134 480 290218
rect -2916 289898 -1814 290134
rect -1578 289898 480 290134
rect -2916 289876 480 289898
rect 583520 290454 586840 290476
rect 583520 290218 585502 290454
rect 585738 290218 586840 290454
rect 583520 290134 586840 290218
rect 583520 289898 585502 290134
rect 585738 289898 586840 290134
rect 583520 289876 586840 289898
rect -1996 289874 -1396 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 591760 283276 592360 283278
rect -8436 283254 480 283276
rect -8436 283018 -8254 283254
rect -8018 283018 480 283254
rect -8436 282934 480 283018
rect -8436 282698 -8254 282934
rect -8018 282698 480 282934
rect -8436 282676 480 282698
rect 583520 283254 592360 283276
rect 583520 283018 591942 283254
rect 592178 283018 592360 283254
rect 583520 282934 592360 283018
rect 583520 282698 591942 282934
rect 592178 282698 592360 282934
rect 583520 282676 592360 282698
rect -8436 282674 -7836 282676
rect 591760 282674 592360 282676
rect 339048 281750 339416 281774
rect 339048 281430 339072 281750
rect 339392 281430 339416 281750
rect 339048 281406 339416 281430
rect -6596 279676 -5996 279678
rect 339072 279676 339392 281406
rect 589920 279676 590520 279678
rect -6596 279654 480 279676
rect -6596 279418 -6414 279654
rect -6178 279418 480 279654
rect -6596 279334 480 279418
rect -6596 279098 -6414 279334
rect -6178 279098 480 279334
rect -6596 279076 480 279098
rect 337710 279654 590520 279676
rect 337710 279418 590102 279654
rect 590338 279418 590520 279654
rect 337710 279334 590520 279418
rect 337710 279098 590102 279334
rect 590338 279098 590520 279334
rect 337710 279076 590520 279098
rect -6596 279074 -5996 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 588080 276076 588680 276078
rect -4756 276054 480 276076
rect -4756 275818 -4574 276054
rect -4338 275818 480 276054
rect -4756 275734 480 275818
rect -4756 275498 -4574 275734
rect -4338 275498 480 275734
rect -4756 275476 480 275498
rect 583520 276054 588680 276076
rect 583520 275818 588262 276054
rect 588498 275818 588680 276054
rect 583520 275734 588680 275818
rect 583520 275498 588262 275734
rect 588498 275498 588680 275734
rect 583520 275476 588680 275498
rect -4756 275474 -4156 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 586240 272476 586840 272478
rect -2916 272454 480 272476
rect -2916 272218 -2734 272454
rect -2498 272218 480 272454
rect -2916 272134 480 272218
rect -2916 271898 -2734 272134
rect -2498 271898 480 272134
rect -2916 271876 480 271898
rect 583520 272454 586840 272476
rect 583520 272218 586422 272454
rect 586658 272218 586840 272454
rect 583520 272134 586840 272218
rect 583520 271898 586422 272134
rect 586658 271898 586840 272134
rect 583520 271876 586840 271898
rect -2916 271874 -2316 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 590840 265276 591440 265278
rect -8436 265254 480 265276
rect -8436 265018 -7334 265254
rect -7098 265018 480 265254
rect -8436 264934 480 265018
rect -8436 264698 -7334 264934
rect -7098 264698 480 264934
rect -8436 264676 480 264698
rect 583520 265254 592360 265276
rect 583520 265018 591022 265254
rect 591258 265018 592360 265254
rect 583520 264934 592360 265018
rect 583520 264698 591022 264934
rect 591258 264698 592360 264934
rect 583520 264676 592360 264698
rect -7516 264674 -6916 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 589000 261676 589600 261678
rect -6596 261654 480 261676
rect -6596 261418 -5494 261654
rect -5258 261418 480 261654
rect -6596 261334 480 261418
rect -6596 261098 -5494 261334
rect -5258 261098 480 261334
rect -6596 261076 480 261098
rect 583520 261654 590520 261676
rect 583520 261418 589182 261654
rect 589418 261418 590520 261654
rect 583520 261334 590520 261418
rect 583520 261098 589182 261334
rect 589418 261098 590520 261334
rect 583520 261076 590520 261098
rect -5676 261074 -5076 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 587160 258076 587760 258078
rect -4756 258054 480 258076
rect -4756 257818 -3654 258054
rect -3418 257818 480 258054
rect -4756 257734 480 257818
rect -4756 257498 -3654 257734
rect -3418 257498 480 257734
rect -4756 257476 480 257498
rect 583520 258054 588680 258076
rect 583520 257818 587342 258054
rect 587578 257818 588680 258054
rect 583520 257734 588680 257818
rect 583520 257498 587342 257734
rect 587578 257498 588680 257734
rect 583520 257476 588680 257498
rect -3836 257474 -3236 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 585320 254476 585920 254478
rect -2916 254454 480 254476
rect -2916 254218 -1814 254454
rect -1578 254218 480 254454
rect -2916 254134 480 254218
rect -2916 253898 -1814 254134
rect -1578 253898 480 254134
rect -2916 253876 480 253898
rect 583520 254454 586840 254476
rect 583520 254218 585502 254454
rect 585738 254218 586840 254454
rect 583520 254134 586840 254218
rect 583520 253898 585502 254134
rect 585738 253898 586840 254134
rect 583520 253876 586840 253898
rect -1996 253874 -1396 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 591760 247276 592360 247278
rect -8436 247254 480 247276
rect -8436 247018 -8254 247254
rect -8018 247018 480 247254
rect -8436 246934 480 247018
rect -8436 246698 -8254 246934
rect -8018 246698 480 246934
rect -8436 246676 480 246698
rect 583520 247254 592360 247276
rect 583520 247018 591942 247254
rect 592178 247018 592360 247254
rect 583520 246934 592360 247018
rect 583520 246698 591942 246934
rect 592178 246698 592360 246934
rect 583520 246676 592360 246698
rect -8436 246674 -7836 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 589920 243676 590520 243678
rect -6596 243654 480 243676
rect -6596 243418 -6414 243654
rect -6178 243418 480 243654
rect -6596 243334 480 243418
rect -6596 243098 -6414 243334
rect -6178 243098 480 243334
rect -6596 243076 480 243098
rect 583520 243654 590520 243676
rect 583520 243418 590102 243654
rect 590338 243418 590520 243654
rect 583520 243334 590520 243418
rect 583520 243098 590102 243334
rect 590338 243098 590520 243334
rect 583520 243076 590520 243098
rect -6596 243074 -5996 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 588080 240076 588680 240078
rect -4756 240054 480 240076
rect -4756 239818 -4574 240054
rect -4338 239818 480 240054
rect -4756 239734 480 239818
rect -4756 239498 -4574 239734
rect -4338 239498 480 239734
rect -4756 239476 480 239498
rect 583520 240054 588680 240076
rect 583520 239818 588262 240054
rect 588498 239818 588680 240054
rect 583520 239734 588680 239818
rect 583520 239498 588262 239734
rect 588498 239498 588680 239734
rect 583520 239476 588680 239498
rect -4756 239474 -4156 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 586240 236476 586840 236478
rect -2916 236454 480 236476
rect -2916 236218 -2734 236454
rect -2498 236218 480 236454
rect -2916 236134 480 236218
rect -2916 235898 -2734 236134
rect -2498 235898 480 236134
rect -2916 235876 480 235898
rect 583520 236454 586840 236476
rect 583520 236218 586422 236454
rect 586658 236218 586840 236454
rect 583520 236134 586840 236218
rect 583520 235898 586422 236134
rect 586658 235898 586840 236134
rect 583520 235876 586840 235898
rect -2916 235874 -2316 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 590840 229276 591440 229278
rect -8436 229254 480 229276
rect -8436 229018 -7334 229254
rect -7098 229018 480 229254
rect -8436 228934 480 229018
rect -8436 228698 -7334 228934
rect -7098 228698 480 228934
rect -8436 228676 480 228698
rect 583520 229254 592360 229276
rect 583520 229018 591022 229254
rect 591258 229018 592360 229254
rect 583520 228934 592360 229018
rect 583520 228698 591022 228934
rect 591258 228698 592360 228934
rect 583520 228676 592360 228698
rect -7516 228674 -6916 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 589000 225676 589600 225678
rect -6596 225654 480 225676
rect -6596 225418 -5494 225654
rect -5258 225418 480 225654
rect -6596 225334 480 225418
rect -6596 225098 -5494 225334
rect -5258 225098 480 225334
rect -6596 225076 480 225098
rect 583520 225654 590520 225676
rect 583520 225418 589182 225654
rect 589418 225418 590520 225654
rect 583520 225334 590520 225418
rect 583520 225098 589182 225334
rect 589418 225098 590520 225334
rect 583520 225076 590520 225098
rect -5676 225074 -5076 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 587160 222076 587760 222078
rect -4756 222054 480 222076
rect -4756 221818 -3654 222054
rect -3418 221818 480 222054
rect -4756 221734 480 221818
rect -4756 221498 -3654 221734
rect -3418 221498 480 221734
rect -4756 221476 480 221498
rect 583520 222054 588680 222076
rect 583520 221818 587342 222054
rect 587578 221818 588680 222054
rect 583520 221734 588680 221818
rect 583520 221498 587342 221734
rect 587578 221498 588680 221734
rect 583520 221476 588680 221498
rect -3836 221474 -3236 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 585320 218476 585920 218478
rect -2916 218454 480 218476
rect -2916 218218 -1814 218454
rect -1578 218218 480 218454
rect -2916 218134 480 218218
rect -2916 217898 -1814 218134
rect -1578 217898 480 218134
rect -2916 217876 480 217898
rect 583520 218454 586840 218476
rect 583520 218218 585502 218454
rect 585738 218218 586840 218454
rect 583520 218134 586840 218218
rect 583520 217898 585502 218134
rect 585738 217898 586840 218134
rect 583520 217876 586840 217898
rect -1996 217874 -1396 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 591760 211276 592360 211278
rect -8436 211254 480 211276
rect -8436 211018 -8254 211254
rect -8018 211018 480 211254
rect -8436 210934 480 211018
rect -8436 210698 -8254 210934
rect -8018 210698 480 210934
rect -8436 210676 480 210698
rect 583520 211254 592360 211276
rect 583520 211018 591942 211254
rect 592178 211018 592360 211254
rect 583520 210934 592360 211018
rect 583520 210698 591942 210934
rect 592178 210698 592360 210934
rect 583520 210676 592360 210698
rect -8436 210674 -7836 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 589920 207676 590520 207678
rect -6596 207654 480 207676
rect -6596 207418 -6414 207654
rect -6178 207418 480 207654
rect -6596 207334 480 207418
rect -6596 207098 -6414 207334
rect -6178 207098 480 207334
rect -6596 207076 480 207098
rect 583520 207654 590520 207676
rect 583520 207418 590102 207654
rect 590338 207418 590520 207654
rect 583520 207334 590520 207418
rect 583520 207098 590102 207334
rect 590338 207098 590520 207334
rect 583520 207076 590520 207098
rect -6596 207074 -5996 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 588080 204076 588680 204078
rect -4756 204054 480 204076
rect -4756 203818 -4574 204054
rect -4338 203818 480 204054
rect -4756 203734 480 203818
rect -4756 203498 -4574 203734
rect -4338 203498 480 203734
rect -4756 203476 480 203498
rect 583520 204054 588680 204076
rect 583520 203818 588262 204054
rect 588498 203818 588680 204054
rect 583520 203734 588680 203818
rect 583520 203498 588262 203734
rect 588498 203498 588680 203734
rect 583520 203476 588680 203498
rect -4756 203474 -4156 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 586240 200476 586840 200478
rect -2916 200454 480 200476
rect -2916 200218 -2734 200454
rect -2498 200218 480 200454
rect -2916 200134 480 200218
rect -2916 199898 -2734 200134
rect -2498 199898 480 200134
rect -2916 199876 480 199898
rect 583520 200454 586840 200476
rect 583520 200218 586422 200454
rect 586658 200218 586840 200454
rect 583520 200134 586840 200218
rect 583520 199898 586422 200134
rect 586658 199898 586840 200134
rect 583520 199876 586840 199898
rect -2916 199874 -2316 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 590840 193276 591440 193278
rect -8436 193254 480 193276
rect -8436 193018 -7334 193254
rect -7098 193018 480 193254
rect -8436 192934 480 193018
rect -8436 192698 -7334 192934
rect -7098 192698 480 192934
rect -8436 192676 480 192698
rect 583520 193254 592360 193276
rect 583520 193018 591022 193254
rect 591258 193018 592360 193254
rect 583520 192934 592360 193018
rect 583520 192698 591022 192934
rect 591258 192698 592360 192934
rect 583520 192676 592360 192698
rect -7516 192674 -6916 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 589000 189676 589600 189678
rect -6596 189654 480 189676
rect -6596 189418 -5494 189654
rect -5258 189418 480 189654
rect -6596 189334 480 189418
rect -6596 189098 -5494 189334
rect -5258 189098 480 189334
rect -6596 189076 480 189098
rect 583520 189654 590520 189676
rect 583520 189418 589182 189654
rect 589418 189418 590520 189654
rect 583520 189334 590520 189418
rect 583520 189098 589182 189334
rect 589418 189098 590520 189334
rect 583520 189076 590520 189098
rect -5676 189074 -5076 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 587160 186076 587760 186078
rect -4756 186054 480 186076
rect -4756 185818 -3654 186054
rect -3418 185818 480 186054
rect -4756 185734 480 185818
rect -4756 185498 -3654 185734
rect -3418 185498 480 185734
rect -4756 185476 480 185498
rect 583520 186054 588680 186076
rect 583520 185818 587342 186054
rect 587578 185818 588680 186054
rect 583520 185734 588680 185818
rect 583520 185498 587342 185734
rect 587578 185498 588680 185734
rect 583520 185476 588680 185498
rect -3836 185474 -3236 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 585320 182476 585920 182478
rect -2916 182454 480 182476
rect -2916 182218 -1814 182454
rect -1578 182218 480 182454
rect -2916 182134 480 182218
rect -2916 181898 -1814 182134
rect -1578 181898 480 182134
rect -2916 181876 480 181898
rect 583520 182454 586840 182476
rect 583520 182218 585502 182454
rect 585738 182218 586840 182454
rect 583520 182134 586840 182218
rect 583520 181898 585502 182134
rect 585738 181898 586840 182134
rect 583520 181876 586840 181898
rect -1996 181874 -1396 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 591760 175276 592360 175278
rect -8436 175254 480 175276
rect -8436 175018 -8254 175254
rect -8018 175018 480 175254
rect -8436 174934 480 175018
rect -8436 174698 -8254 174934
rect -8018 174698 480 174934
rect -8436 174676 480 174698
rect 583520 175254 592360 175276
rect 583520 175018 591942 175254
rect 592178 175018 592360 175254
rect 583520 174934 592360 175018
rect 583520 174698 591942 174934
rect 592178 174698 592360 174934
rect 583520 174676 592360 174698
rect -8436 174674 -7836 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 589920 171676 590520 171678
rect -6596 171654 480 171676
rect -6596 171418 -6414 171654
rect -6178 171418 480 171654
rect -6596 171334 480 171418
rect -6596 171098 -6414 171334
rect -6178 171098 480 171334
rect -6596 171076 480 171098
rect 583520 171654 590520 171676
rect 583520 171418 590102 171654
rect 590338 171418 590520 171654
rect 583520 171334 590520 171418
rect 583520 171098 590102 171334
rect 590338 171098 590520 171334
rect 583520 171076 590520 171098
rect -6596 171074 -5996 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 588080 168076 588680 168078
rect -4756 168054 480 168076
rect -4756 167818 -4574 168054
rect -4338 167818 480 168054
rect -4756 167734 480 167818
rect -4756 167498 -4574 167734
rect -4338 167498 480 167734
rect -4756 167476 480 167498
rect 583520 168054 588680 168076
rect 583520 167818 588262 168054
rect 588498 167818 588680 168054
rect 583520 167734 588680 167818
rect 583520 167498 588262 167734
rect 588498 167498 588680 167734
rect 583520 167476 588680 167498
rect -4756 167474 -4156 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 586240 164476 586840 164478
rect -2916 164454 480 164476
rect -2916 164218 -2734 164454
rect -2498 164218 480 164454
rect -2916 164134 480 164218
rect -2916 163898 -2734 164134
rect -2498 163898 480 164134
rect -2916 163876 480 163898
rect 583520 164454 586840 164476
rect 583520 164218 586422 164454
rect 586658 164218 586840 164454
rect 583520 164134 586840 164218
rect 583520 163898 586422 164134
rect 586658 163898 586840 164134
rect 583520 163876 586840 163898
rect -2916 163874 -2316 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 590840 157276 591440 157278
rect -8436 157254 480 157276
rect -8436 157018 -7334 157254
rect -7098 157018 480 157254
rect -8436 156934 480 157018
rect -8436 156698 -7334 156934
rect -7098 156698 480 156934
rect -8436 156676 480 156698
rect 583520 157254 592360 157276
rect 583520 157018 591022 157254
rect 591258 157018 592360 157254
rect 583520 156934 592360 157018
rect 583520 156698 591022 156934
rect 591258 156698 592360 156934
rect 583520 156676 592360 156698
rect -7516 156674 -6916 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 589000 153676 589600 153678
rect -6596 153654 480 153676
rect -6596 153418 -5494 153654
rect -5258 153418 480 153654
rect -6596 153334 480 153418
rect -6596 153098 -5494 153334
rect -5258 153098 480 153334
rect -6596 153076 480 153098
rect 583520 153654 590520 153676
rect 583520 153418 589182 153654
rect 589418 153418 590520 153654
rect 583520 153334 590520 153418
rect 583520 153098 589182 153334
rect 589418 153098 590520 153334
rect 583520 153076 590520 153098
rect -5676 153074 -5076 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 587160 150076 587760 150078
rect -4756 150054 480 150076
rect -4756 149818 -3654 150054
rect -3418 149818 480 150054
rect -4756 149734 480 149818
rect -4756 149498 -3654 149734
rect -3418 149498 480 149734
rect -4756 149476 480 149498
rect 583520 150054 588680 150076
rect 583520 149818 587342 150054
rect 587578 149818 588680 150054
rect 583520 149734 588680 149818
rect 583520 149498 587342 149734
rect 587578 149498 588680 149734
rect 583520 149476 588680 149498
rect -3836 149474 -3236 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 585320 146476 585920 146478
rect -2916 146454 480 146476
rect -2916 146218 -1814 146454
rect -1578 146218 480 146454
rect -2916 146134 480 146218
rect -2916 145898 -1814 146134
rect -1578 145898 480 146134
rect -2916 145876 480 145898
rect 583520 146454 586840 146476
rect 583520 146218 585502 146454
rect 585738 146218 586840 146454
rect 583520 146134 586840 146218
rect 583520 145898 585502 146134
rect 585738 145898 586840 146134
rect 583520 145876 586840 145898
rect -1996 145874 -1396 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 591760 139276 592360 139278
rect -8436 139254 480 139276
rect -8436 139018 -8254 139254
rect -8018 139018 480 139254
rect -8436 138934 480 139018
rect -8436 138698 -8254 138934
rect -8018 138698 480 138934
rect -8436 138676 480 138698
rect 583520 139254 592360 139276
rect 583520 139018 591942 139254
rect 592178 139018 592360 139254
rect 583520 138934 592360 139018
rect 583520 138698 591942 138934
rect 592178 138698 592360 138934
rect 583520 138676 592360 138698
rect -8436 138674 -7836 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 589920 135676 590520 135678
rect -6596 135654 480 135676
rect -6596 135418 -6414 135654
rect -6178 135418 480 135654
rect -6596 135334 480 135418
rect -6596 135098 -6414 135334
rect -6178 135098 480 135334
rect -6596 135076 480 135098
rect 583520 135654 590520 135676
rect 583520 135418 590102 135654
rect 590338 135418 590520 135654
rect 583520 135334 590520 135418
rect 583520 135098 590102 135334
rect 590338 135098 590520 135334
rect 583520 135076 590520 135098
rect -6596 135074 -5996 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 588080 132076 588680 132078
rect -4756 132054 480 132076
rect -4756 131818 -4574 132054
rect -4338 131818 480 132054
rect -4756 131734 480 131818
rect -4756 131498 -4574 131734
rect -4338 131498 480 131734
rect -4756 131476 480 131498
rect 583520 132054 588680 132076
rect 583520 131818 588262 132054
rect 588498 131818 588680 132054
rect 583520 131734 588680 131818
rect 583520 131498 588262 131734
rect 588498 131498 588680 131734
rect 583520 131476 588680 131498
rect -4756 131474 -4156 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 586240 128476 586840 128478
rect -2916 128454 480 128476
rect -2916 128218 -2734 128454
rect -2498 128218 480 128454
rect -2916 128134 480 128218
rect -2916 127898 -2734 128134
rect -2498 127898 480 128134
rect -2916 127876 480 127898
rect 583520 128454 586840 128476
rect 583520 128218 586422 128454
rect 586658 128218 586840 128454
rect 583520 128134 586840 128218
rect 583520 127898 586422 128134
rect 586658 127898 586840 128134
rect 583520 127876 586840 127898
rect -2916 127874 -2316 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 590840 121276 591440 121278
rect -8436 121254 480 121276
rect -8436 121018 -7334 121254
rect -7098 121018 480 121254
rect -8436 120934 480 121018
rect -8436 120698 -7334 120934
rect -7098 120698 480 120934
rect -8436 120676 480 120698
rect 583520 121254 592360 121276
rect 583520 121018 591022 121254
rect 591258 121018 592360 121254
rect 583520 120934 592360 121018
rect 583520 120698 591022 120934
rect 591258 120698 592360 120934
rect 583520 120676 592360 120698
rect -7516 120674 -6916 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 589000 117676 589600 117678
rect -6596 117654 480 117676
rect -6596 117418 -5494 117654
rect -5258 117418 480 117654
rect -6596 117334 480 117418
rect -6596 117098 -5494 117334
rect -5258 117098 480 117334
rect -6596 117076 480 117098
rect 583520 117654 590520 117676
rect 583520 117418 589182 117654
rect 589418 117418 590520 117654
rect 583520 117334 590520 117418
rect 583520 117098 589182 117334
rect 589418 117098 590520 117334
rect 583520 117076 590520 117098
rect -5676 117074 -5076 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 587160 114076 587760 114078
rect -4756 114054 480 114076
rect -4756 113818 -3654 114054
rect -3418 113818 480 114054
rect -4756 113734 480 113818
rect -4756 113498 -3654 113734
rect -3418 113498 480 113734
rect -4756 113476 480 113498
rect 583520 114054 588680 114076
rect 583520 113818 587342 114054
rect 587578 113818 588680 114054
rect 583520 113734 588680 113818
rect 583520 113498 587342 113734
rect 587578 113498 588680 113734
rect 583520 113476 588680 113498
rect -3836 113474 -3236 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 585320 110476 585920 110478
rect -2916 110454 480 110476
rect -2916 110218 -1814 110454
rect -1578 110218 480 110454
rect -2916 110134 480 110218
rect -2916 109898 -1814 110134
rect -1578 109898 480 110134
rect -2916 109876 480 109898
rect 583520 110454 586840 110476
rect 583520 110218 585502 110454
rect 585738 110218 586840 110454
rect 583520 110134 586840 110218
rect 583520 109898 585502 110134
rect 585738 109898 586840 110134
rect 583520 109876 586840 109898
rect -1996 109874 -1396 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 591760 103276 592360 103278
rect -8436 103254 480 103276
rect -8436 103018 -8254 103254
rect -8018 103018 480 103254
rect -8436 102934 480 103018
rect -8436 102698 -8254 102934
rect -8018 102698 480 102934
rect -8436 102676 480 102698
rect 583520 103254 592360 103276
rect 583520 103018 591942 103254
rect 592178 103018 592360 103254
rect 583520 102934 592360 103018
rect 583520 102698 591942 102934
rect 592178 102698 592360 102934
rect 583520 102676 592360 102698
rect -8436 102674 -7836 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 589920 99676 590520 99678
rect -6596 99654 480 99676
rect -6596 99418 -6414 99654
rect -6178 99418 480 99654
rect -6596 99334 480 99418
rect -6596 99098 -6414 99334
rect -6178 99098 480 99334
rect -6596 99076 480 99098
rect 583520 99654 590520 99676
rect 583520 99418 590102 99654
rect 590338 99418 590520 99654
rect 583520 99334 590520 99418
rect 583520 99098 590102 99334
rect 590338 99098 590520 99334
rect 583520 99076 590520 99098
rect -6596 99074 -5996 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 588080 96076 588680 96078
rect -4756 96054 480 96076
rect -4756 95818 -4574 96054
rect -4338 95818 480 96054
rect -4756 95734 480 95818
rect -4756 95498 -4574 95734
rect -4338 95498 480 95734
rect -4756 95476 480 95498
rect 583520 96054 588680 96076
rect 583520 95818 588262 96054
rect 588498 95818 588680 96054
rect 583520 95734 588680 95818
rect 583520 95498 588262 95734
rect 588498 95498 588680 95734
rect 583520 95476 588680 95498
rect -4756 95474 -4156 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 586240 92476 586840 92478
rect -2916 92454 480 92476
rect -2916 92218 -2734 92454
rect -2498 92218 480 92454
rect -2916 92134 480 92218
rect -2916 91898 -2734 92134
rect -2498 91898 480 92134
rect -2916 91876 480 91898
rect 583520 92454 586840 92476
rect 583520 92218 586422 92454
rect 586658 92218 586840 92454
rect 583520 92134 586840 92218
rect 583520 91898 586422 92134
rect 586658 91898 586840 92134
rect 583520 91876 586840 91898
rect -2916 91874 -2316 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 590840 85276 591440 85278
rect -8436 85254 480 85276
rect -8436 85018 -7334 85254
rect -7098 85018 480 85254
rect -8436 84934 480 85018
rect -8436 84698 -7334 84934
rect -7098 84698 480 84934
rect -8436 84676 480 84698
rect 583520 85254 592360 85276
rect 583520 85018 591022 85254
rect 591258 85018 592360 85254
rect 583520 84934 592360 85018
rect 583520 84698 591022 84934
rect 591258 84698 592360 84934
rect 583520 84676 592360 84698
rect -7516 84674 -6916 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 589000 81676 589600 81678
rect -6596 81654 480 81676
rect -6596 81418 -5494 81654
rect -5258 81418 480 81654
rect -6596 81334 480 81418
rect -6596 81098 -5494 81334
rect -5258 81098 480 81334
rect -6596 81076 480 81098
rect 583520 81654 590520 81676
rect 583520 81418 589182 81654
rect 589418 81418 590520 81654
rect 583520 81334 590520 81418
rect 583520 81098 589182 81334
rect 589418 81098 590520 81334
rect 583520 81076 590520 81098
rect -5676 81074 -5076 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 587160 78076 587760 78078
rect -4756 78054 480 78076
rect -4756 77818 -3654 78054
rect -3418 77818 480 78054
rect -4756 77734 480 77818
rect -4756 77498 -3654 77734
rect -3418 77498 480 77734
rect -4756 77476 480 77498
rect 583520 78054 588680 78076
rect 583520 77818 587342 78054
rect 587578 77818 588680 78054
rect 583520 77734 588680 77818
rect 583520 77498 587342 77734
rect 587578 77498 588680 77734
rect 583520 77476 588680 77498
rect -3836 77474 -3236 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 585320 74476 585920 74478
rect -2916 74454 480 74476
rect -2916 74218 -1814 74454
rect -1578 74218 480 74454
rect -2916 74134 480 74218
rect -2916 73898 -1814 74134
rect -1578 73898 480 74134
rect -2916 73876 480 73898
rect 583520 74454 586840 74476
rect 583520 74218 585502 74454
rect 585738 74218 586840 74454
rect 583520 74134 586840 74218
rect 583520 73898 585502 74134
rect 585738 73898 586840 74134
rect 583520 73876 586840 73898
rect -1996 73874 -1396 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 591760 67276 592360 67278
rect -8436 67254 480 67276
rect -8436 67018 -8254 67254
rect -8018 67018 480 67254
rect -8436 66934 480 67018
rect -8436 66698 -8254 66934
rect -8018 66698 480 66934
rect -8436 66676 480 66698
rect 583520 67254 592360 67276
rect 583520 67018 591942 67254
rect 592178 67018 592360 67254
rect 583520 66934 592360 67018
rect 583520 66698 591942 66934
rect 592178 66698 592360 66934
rect 583520 66676 592360 66698
rect -8436 66674 -7836 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 589920 63676 590520 63678
rect -6596 63654 480 63676
rect -6596 63418 -6414 63654
rect -6178 63418 480 63654
rect -6596 63334 480 63418
rect -6596 63098 -6414 63334
rect -6178 63098 480 63334
rect -6596 63076 480 63098
rect 583520 63654 590520 63676
rect 583520 63418 590102 63654
rect 590338 63418 590520 63654
rect 583520 63334 590520 63418
rect 583520 63098 590102 63334
rect 590338 63098 590520 63334
rect 583520 63076 590520 63098
rect -6596 63074 -5996 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 588080 60076 588680 60078
rect -4756 60054 480 60076
rect -4756 59818 -4574 60054
rect -4338 59818 480 60054
rect -4756 59734 480 59818
rect -4756 59498 -4574 59734
rect -4338 59498 480 59734
rect -4756 59476 480 59498
rect 583520 60054 588680 60076
rect 583520 59818 588262 60054
rect 588498 59818 588680 60054
rect 583520 59734 588680 59818
rect 583520 59498 588262 59734
rect 588498 59498 588680 59734
rect 583520 59476 588680 59498
rect -4756 59474 -4156 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 586240 56476 586840 56478
rect -2916 56454 480 56476
rect -2916 56218 -2734 56454
rect -2498 56218 480 56454
rect -2916 56134 480 56218
rect -2916 55898 -2734 56134
rect -2498 55898 480 56134
rect -2916 55876 480 55898
rect 583520 56454 586840 56476
rect 583520 56218 586422 56454
rect 586658 56218 586840 56454
rect 583520 56134 586840 56218
rect 583520 55898 586422 56134
rect 586658 55898 586840 56134
rect 583520 55876 586840 55898
rect -2916 55874 -2316 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 590840 49276 591440 49278
rect -8436 49254 480 49276
rect -8436 49018 -7334 49254
rect -7098 49018 480 49254
rect -8436 48934 480 49018
rect -8436 48698 -7334 48934
rect -7098 48698 480 48934
rect -8436 48676 480 48698
rect 583520 49254 592360 49276
rect 583520 49018 591022 49254
rect 591258 49018 592360 49254
rect 583520 48934 592360 49018
rect 583520 48698 591022 48934
rect 591258 48698 592360 48934
rect 583520 48676 592360 48698
rect -7516 48674 -6916 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 589000 45676 589600 45678
rect -6596 45654 480 45676
rect -6596 45418 -5494 45654
rect -5258 45418 480 45654
rect -6596 45334 480 45418
rect -6596 45098 -5494 45334
rect -5258 45098 480 45334
rect -6596 45076 480 45098
rect 583520 45654 590520 45676
rect 583520 45418 589182 45654
rect 589418 45418 590520 45654
rect 583520 45334 590520 45418
rect 583520 45098 589182 45334
rect 589418 45098 590520 45334
rect 583520 45076 590520 45098
rect -5676 45074 -5076 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 587160 42076 587760 42078
rect -4756 42054 480 42076
rect -4756 41818 -3654 42054
rect -3418 41818 480 42054
rect -4756 41734 480 41818
rect -4756 41498 -3654 41734
rect -3418 41498 480 41734
rect -4756 41476 480 41498
rect 583520 42054 588680 42076
rect 583520 41818 587342 42054
rect 587578 41818 588680 42054
rect 583520 41734 588680 41818
rect 583520 41498 587342 41734
rect 587578 41498 588680 41734
rect 583520 41476 588680 41498
rect -3836 41474 -3236 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 585320 38476 585920 38478
rect -2916 38454 480 38476
rect -2916 38218 -1814 38454
rect -1578 38218 480 38454
rect -2916 38134 480 38218
rect -2916 37898 -1814 38134
rect -1578 37898 480 38134
rect -2916 37876 480 37898
rect 583520 38454 586840 38476
rect 583520 38218 585502 38454
rect 585738 38218 586840 38454
rect 583520 38134 586840 38218
rect 583520 37898 585502 38134
rect 585738 37898 586840 38134
rect 583520 37876 586840 37898
rect -1996 37874 -1396 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 591760 31276 592360 31278
rect -8436 31254 480 31276
rect -8436 31018 -8254 31254
rect -8018 31018 480 31254
rect -8436 30934 480 31018
rect -8436 30698 -8254 30934
rect -8018 30698 480 30934
rect -8436 30676 480 30698
rect 583520 31254 592360 31276
rect 583520 31018 591942 31254
rect 592178 31018 592360 31254
rect 583520 30934 592360 31018
rect 583520 30698 591942 30934
rect 592178 30698 592360 30934
rect 583520 30676 592360 30698
rect -8436 30674 -7836 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 589920 27676 590520 27678
rect -6596 27654 480 27676
rect -6596 27418 -6414 27654
rect -6178 27418 480 27654
rect -6596 27334 480 27418
rect -6596 27098 -6414 27334
rect -6178 27098 480 27334
rect -6596 27076 480 27098
rect 583520 27654 590520 27676
rect 583520 27418 590102 27654
rect 590338 27418 590520 27654
rect 583520 27334 590520 27418
rect 583520 27098 590102 27334
rect 590338 27098 590520 27334
rect 583520 27076 590520 27098
rect -6596 27074 -5996 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 588080 24076 588680 24078
rect -4756 24054 480 24076
rect -4756 23818 -4574 24054
rect -4338 23818 480 24054
rect -4756 23734 480 23818
rect -4756 23498 -4574 23734
rect -4338 23498 480 23734
rect -4756 23476 480 23498
rect 583520 24054 588680 24076
rect 583520 23818 588262 24054
rect 588498 23818 588680 24054
rect 583520 23734 588680 23818
rect 583520 23498 588262 23734
rect 588498 23498 588680 23734
rect 583520 23476 588680 23498
rect -4756 23474 -4156 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 586240 20476 586840 20478
rect -2916 20454 480 20476
rect -2916 20218 -2734 20454
rect -2498 20218 480 20454
rect -2916 20134 480 20218
rect -2916 19898 -2734 20134
rect -2498 19898 480 20134
rect -2916 19876 480 19898
rect 583520 20454 586840 20476
rect 583520 20218 586422 20454
rect 586658 20218 586840 20454
rect 583520 20134 586840 20218
rect 583520 19898 586422 20134
rect 586658 19898 586840 20134
rect 583520 19876 586840 19898
rect -2916 19874 -2316 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 590840 13276 591440 13278
rect -8436 13254 480 13276
rect -8436 13018 -7334 13254
rect -7098 13018 480 13254
rect -8436 12934 480 13018
rect -8436 12698 -7334 12934
rect -7098 12698 480 12934
rect -8436 12676 480 12698
rect 583520 13254 592360 13276
rect 583520 13018 591022 13254
rect 591258 13018 592360 13254
rect 583520 12934 592360 13018
rect 583520 12698 591022 12934
rect 591258 12698 592360 12934
rect 583520 12676 592360 12698
rect -7516 12674 -6916 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 589000 9676 589600 9678
rect -6596 9654 480 9676
rect -6596 9418 -5494 9654
rect -5258 9418 480 9654
rect -6596 9334 480 9418
rect -6596 9098 -5494 9334
rect -5258 9098 480 9334
rect -6596 9076 480 9098
rect 583520 9654 590520 9676
rect 583520 9418 589182 9654
rect 589418 9418 590520 9654
rect 583520 9334 590520 9418
rect 583520 9098 589182 9334
rect 589418 9098 590520 9334
rect 583520 9076 590520 9098
rect -5676 9074 -5076 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 587160 6076 587760 6078
rect -4756 6054 480 6076
rect -4756 5818 -3654 6054
rect -3418 5818 480 6054
rect -4756 5734 480 5818
rect -4756 5498 -3654 5734
rect -3418 5498 480 5734
rect -4756 5476 480 5498
rect 583520 6054 588680 6076
rect 583520 5818 587342 6054
rect 587578 5818 588680 6054
rect 583520 5734 588680 5818
rect 583520 5498 587342 5734
rect 587578 5498 588680 5734
rect 583520 5476 588680 5498
rect -3836 5474 -3236 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 585320 2476 585920 2478
rect -2916 2454 480 2476
rect -2916 2218 -1814 2454
rect -1578 2218 480 2454
rect -2916 2134 480 2218
rect -2916 1898 -1814 2134
rect -1578 1898 480 2134
rect -2916 1876 480 1898
rect 583520 2454 586840 2476
rect 583520 2218 585502 2454
rect 585738 2218 586840 2454
rect 583520 2134 586840 2218
rect 583520 1898 585502 2134
rect 585738 1898 586840 2134
rect 583520 1876 586840 1898
rect -1996 1874 -1396 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use chip-w-opamp  chip-w-opamp_0
timestamp 1606718978
transform 1 0 341468 0 1 448419
box -25936 -8570 19927 24418
use 10good  10good_0
timestamp 1607536219
transform -1 0 142580 0 -1 320426
box -738 -22 79994 49740
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 4 analog_io[0]
port 1 nsew
rlabel metal3 s 583520 474996 584960 475236 4 analog_io[10]
port 2 nsew
rlabel metal3 s 583520 521916 584960 522156 4 analog_io[11]
port 3 nsew
rlabel metal3 s 583520 568836 584960 569076 4 analog_io[12]
port 4 nsew
rlabel metal3 s 583520 615756 584960 615996 4 analog_io[13]
port 5 nsew
rlabel metal3 s 583520 662676 584960 662916 4 analog_io[14]
port 6 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[15]
port 7 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[16]
port 8 nsew
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[17]
port 9 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[18]
port 10 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 52716 584960 52956 4 analog_io[1]
port 12 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[20]
port 13 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[21]
port 14 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[22]
port 15 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 21 nsew
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 22 nsew
rlabel metal3 s 583520 99636 584960 99876 4 analog_io[2]
port 23 nsew
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 24 nsew
rlabel metal3 s 583520 146556 584960 146796 4 analog_io[3]
port 25 nsew
rlabel metal3 s 583520 193476 584960 193716 4 analog_io[4]
port 26 nsew
rlabel metal3 s 583520 240396 584960 240636 4 analog_io[5]
port 27 nsew
rlabel metal3 s 583520 287316 584960 287556 4 analog_io[6]
port 28 nsew
rlabel metal3 s 583520 334236 584960 334476 4 analog_io[7]
port 29 nsew
rlabel metal3 s 583520 381156 584960 381396 4 analog_io[8]
port 30 nsew
rlabel metal3 s 583520 428076 584960 428316 4 analog_io[9]
port 31 nsew
rlabel metal3 s 583520 17492 584960 17732 4 io_in[0]
port 32 nsew
rlabel metal3 s 583520 486692 584960 486932 4 io_in[10]
port 33 nsew
rlabel metal3 s 583520 533748 584960 533988 4 io_in[11]
port 34 nsew
rlabel metal3 s 583520 580668 584960 580908 4 io_in[12]
port 35 nsew
rlabel metal3 s 583520 627588 584960 627828 4 io_in[13]
port 36 nsew
rlabel metal3 s 583520 674508 584960 674748 4 io_in[14]
port 37 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 38 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 39 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 40 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 41 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 42 nsew
rlabel metal3 s 583520 64412 584960 64652 4 io_in[1]
port 43 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 44 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 45 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 46 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 47 nsew
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 48 nsew
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 49 nsew
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 50 nsew
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 51 nsew
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 52 nsew
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 53 nsew
rlabel metal3 s 583520 111332 584960 111572 4 io_in[2]
port 54 nsew
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 55 nsew
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 56 nsew
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 57 nsew
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 58 nsew
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 59 nsew
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 60 nsew
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 61 nsew
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 62 nsew
rlabel metal3 s 583520 158252 584960 158492 4 io_in[3]
port 63 nsew
rlabel metal3 s 583520 205172 584960 205412 4 io_in[4]
port 64 nsew
rlabel metal3 s 583520 252092 584960 252332 4 io_in[5]
port 65 nsew
rlabel metal3 s 583520 299012 584960 299252 4 io_in[6]
port 66 nsew
rlabel metal3 s 583520 345932 584960 346172 4 io_in[7]
port 67 nsew
rlabel metal3 s 583520 392852 584960 393092 4 io_in[8]
port 68 nsew
rlabel metal3 s 583520 439772 584960 440012 4 io_in[9]
port 69 nsew
rlabel metal3 s 583520 40884 584960 41124 4 io_oeb[0]
port 70 nsew
rlabel metal3 s 583520 510220 584960 510460 4 io_oeb[10]
port 71 nsew
rlabel metal3 s 583520 557140 584960 557380 4 io_oeb[11]
port 72 nsew
rlabel metal3 s 583520 604060 584960 604300 4 io_oeb[12]
port 73 nsew
rlabel metal3 s 583520 650980 584960 651220 4 io_oeb[13]
port 74 nsew
rlabel metal3 s 583520 697900 584960 698140 4 io_oeb[14]
port 75 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 76 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 77 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 78 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 79 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 80 nsew
rlabel metal3 s 583520 87804 584960 88044 4 io_oeb[1]
port 81 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 82 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 83 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 84 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 85 nsew
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 86 nsew
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 87 nsew
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 88 nsew
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 89 nsew
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 90 nsew
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 91 nsew
rlabel metal3 s 583520 134724 584960 134964 4 io_oeb[2]
port 92 nsew
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 93 nsew
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 94 nsew
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 95 nsew
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 96 nsew
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 97 nsew
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 98 nsew
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 99 nsew
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 100 nsew
rlabel metal3 s 583520 181780 584960 182020 4 io_oeb[3]
port 101 nsew
rlabel metal3 s 583520 228700 584960 228940 4 io_oeb[4]
port 102 nsew
rlabel metal3 s 583520 275620 584960 275860 4 io_oeb[5]
port 103 nsew
rlabel metal3 s 583520 322540 584960 322780 4 io_oeb[6]
port 104 nsew
rlabel metal3 s 583520 369460 584960 369700 4 io_oeb[7]
port 105 nsew
rlabel metal3 s 583520 416380 584960 416620 4 io_oeb[8]
port 106 nsew
rlabel metal3 s 583520 463300 584960 463540 4 io_oeb[9]
port 107 nsew
rlabel metal3 s 583520 29188 584960 29428 4 io_out[0]
port 108 nsew
rlabel metal3 s 583520 498524 584960 498764 4 io_out[10]
port 109 nsew
rlabel metal3 s 583520 545444 584960 545684 4 io_out[11]
port 110 nsew
rlabel metal3 s 583520 592364 584960 592604 4 io_out[12]
port 111 nsew
rlabel metal3 s 583520 639284 584960 639524 4 io_out[13]
port 112 nsew
rlabel metal3 s 583520 686204 584960 686444 4 io_out[14]
port 113 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 114 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 115 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 116 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 117 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 118 nsew
rlabel metal3 s 583520 76108 584960 76348 4 io_out[1]
port 119 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 120 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 121 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 122 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 123 nsew
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 124 nsew
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 125 nsew
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 126 nsew
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 127 nsew
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 128 nsew
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 129 nsew
rlabel metal3 s 583520 123028 584960 123268 4 io_out[2]
port 130 nsew
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 131 nsew
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 132 nsew
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 133 nsew
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 134 nsew
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 135 nsew
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 136 nsew
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 137 nsew
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 138 nsew
rlabel metal3 s 583520 169948 584960 170188 4 io_out[3]
port 139 nsew
rlabel metal3 s 583520 216868 584960 217108 4 io_out[4]
port 140 nsew
rlabel metal3 s 583520 263788 584960 264028 4 io_out[5]
port 141 nsew
rlabel metal3 s 583520 310708 584960 310948 4 io_out[6]
port 142 nsew
rlabel metal3 s 583520 357764 584960 358004 4 io_out[7]
port 143 nsew
rlabel metal3 s 583520 404684 584960 404924 4 io_out[8]
port 144 nsew
rlabel metal3 s 583520 451604 584960 451844 4 io_out[9]
port 145 nsew
rlabel metal2 s 126582 -960 126694 480 4 la_data_in[0]
port 146 nsew
rlabel metal2 s 483450 -960 483562 480 4 la_data_in[100]
port 147 nsew
rlabel metal2 s 486946 -960 487058 480 4 la_data_in[101]
port 148 nsew
rlabel metal2 s 490534 -960 490646 480 4 la_data_in[102]
port 149 nsew
rlabel metal2 s 494122 -960 494234 480 4 la_data_in[103]
port 150 nsew
rlabel metal2 s 497710 -960 497822 480 4 la_data_in[104]
port 151 nsew
rlabel metal2 s 501206 -960 501318 480 4 la_data_in[105]
port 152 nsew
rlabel metal2 s 504794 -960 504906 480 4 la_data_in[106]
port 153 nsew
rlabel metal2 s 508382 -960 508494 480 4 la_data_in[107]
port 154 nsew
rlabel metal2 s 511970 -960 512082 480 4 la_data_in[108]
port 155 nsew
rlabel metal2 s 515558 -960 515670 480 4 la_data_in[109]
port 156 nsew
rlabel metal2 s 162278 -960 162390 480 4 la_data_in[10]
port 157 nsew
rlabel metal2 s 519054 -960 519166 480 4 la_data_in[110]
port 158 nsew
rlabel metal2 s 522642 -960 522754 480 4 la_data_in[111]
port 159 nsew
rlabel metal2 s 526230 -960 526342 480 4 la_data_in[112]
port 160 nsew
rlabel metal2 s 529818 -960 529930 480 4 la_data_in[113]
port 161 nsew
rlabel metal2 s 533406 -960 533518 480 4 la_data_in[114]
port 162 nsew
rlabel metal2 s 536902 -960 537014 480 4 la_data_in[115]
port 163 nsew
rlabel metal2 s 540490 -960 540602 480 4 la_data_in[116]
port 164 nsew
rlabel metal2 s 544078 -960 544190 480 4 la_data_in[117]
port 165 nsew
rlabel metal2 s 547666 -960 547778 480 4 la_data_in[118]
port 166 nsew
rlabel metal2 s 551162 -960 551274 480 4 la_data_in[119]
port 167 nsew
rlabel metal2 s 165866 -960 165978 480 4 la_data_in[11]
port 168 nsew
rlabel metal2 s 554750 -960 554862 480 4 la_data_in[120]
port 169 nsew
rlabel metal2 s 558338 -960 558450 480 4 la_data_in[121]
port 170 nsew
rlabel metal2 s 561926 -960 562038 480 4 la_data_in[122]
port 171 nsew
rlabel metal2 s 565514 -960 565626 480 4 la_data_in[123]
port 172 nsew
rlabel metal2 s 569010 -960 569122 480 4 la_data_in[124]
port 173 nsew
rlabel metal2 s 572598 -960 572710 480 4 la_data_in[125]
port 174 nsew
rlabel metal2 s 576186 -960 576298 480 4 la_data_in[126]
port 175 nsew
rlabel metal2 s 579774 -960 579886 480 4 la_data_in[127]
port 176 nsew
rlabel metal2 s 169362 -960 169474 480 4 la_data_in[12]
port 177 nsew
rlabel metal2 s 172950 -960 173062 480 4 la_data_in[13]
port 178 nsew
rlabel metal2 s 176538 -960 176650 480 4 la_data_in[14]
port 179 nsew
rlabel metal2 s 180126 -960 180238 480 4 la_data_in[15]
port 180 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_in[16]
port 181 nsew
rlabel metal2 s 187210 -960 187322 480 4 la_data_in[17]
port 182 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_in[18]
port 183 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_in[19]
port 184 nsew
rlabel metal2 s 130170 -960 130282 480 4 la_data_in[1]
port 185 nsew
rlabel metal2 s 197974 -960 198086 480 4 la_data_in[20]
port 186 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_in[21]
port 187 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_in[22]
port 188 nsew
rlabel metal2 s 208646 -960 208758 480 4 la_data_in[23]
port 189 nsew
rlabel metal2 s 212234 -960 212346 480 4 la_data_in[24]
port 190 nsew
rlabel metal2 s 215822 -960 215934 480 4 la_data_in[25]
port 191 nsew
rlabel metal2 s 219318 -960 219430 480 4 la_data_in[26]
port 192 nsew
rlabel metal2 s 222906 -960 223018 480 4 la_data_in[27]
port 193 nsew
rlabel metal2 s 226494 -960 226606 480 4 la_data_in[28]
port 194 nsew
rlabel metal2 s 230082 -960 230194 480 4 la_data_in[29]
port 195 nsew
rlabel metal2 s 133758 -960 133870 480 4 la_data_in[2]
port 196 nsew
rlabel metal2 s 233670 -960 233782 480 4 la_data_in[30]
port 197 nsew
rlabel metal2 s 237166 -960 237278 480 4 la_data_in[31]
port 198 nsew
rlabel metal2 s 240754 -960 240866 480 4 la_data_in[32]
port 199 nsew
rlabel metal2 s 244342 -960 244454 480 4 la_data_in[33]
port 200 nsew
rlabel metal2 s 247930 -960 248042 480 4 la_data_in[34]
port 201 nsew
rlabel metal2 s 251426 -960 251538 480 4 la_data_in[35]
port 202 nsew
rlabel metal2 s 255014 -960 255126 480 4 la_data_in[36]
port 203 nsew
rlabel metal2 s 258602 -960 258714 480 4 la_data_in[37]
port 204 nsew
rlabel metal2 s 262190 -960 262302 480 4 la_data_in[38]
port 205 nsew
rlabel metal2 s 265778 -960 265890 480 4 la_data_in[39]
port 206 nsew
rlabel metal2 s 137254 -960 137366 480 4 la_data_in[3]
port 207 nsew
rlabel metal2 s 269274 -960 269386 480 4 la_data_in[40]
port 208 nsew
rlabel metal2 s 272862 -960 272974 480 4 la_data_in[41]
port 209 nsew
rlabel metal2 s 276450 -960 276562 480 4 la_data_in[42]
port 210 nsew
rlabel metal2 s 280038 -960 280150 480 4 la_data_in[43]
port 211 nsew
rlabel metal2 s 283626 -960 283738 480 4 la_data_in[44]
port 212 nsew
rlabel metal2 s 287122 -960 287234 480 4 la_data_in[45]
port 213 nsew
rlabel metal2 s 290710 -960 290822 480 4 la_data_in[46]
port 214 nsew
rlabel metal2 s 294298 -960 294410 480 4 la_data_in[47]
port 215 nsew
rlabel metal2 s 297886 -960 297998 480 4 la_data_in[48]
port 216 nsew
rlabel metal2 s 301382 -960 301494 480 4 la_data_in[49]
port 217 nsew
rlabel metal2 s 140842 -960 140954 480 4 la_data_in[4]
port 218 nsew
rlabel metal2 s 304970 -960 305082 480 4 la_data_in[50]
port 219 nsew
rlabel metal2 s 308558 -960 308670 480 4 la_data_in[51]
port 220 nsew
rlabel metal2 s 312146 -960 312258 480 4 la_data_in[52]
port 221 nsew
rlabel metal2 s 315734 -960 315846 480 4 la_data_in[53]
port 222 nsew
rlabel metal2 s 319230 -960 319342 480 4 la_data_in[54]
port 223 nsew
rlabel metal2 s 322818 -960 322930 480 4 la_data_in[55]
port 224 nsew
rlabel metal2 s 326406 -960 326518 480 4 la_data_in[56]
port 225 nsew
rlabel metal2 s 329994 -960 330106 480 4 la_data_in[57]
port 226 nsew
rlabel metal2 s 333582 -960 333694 480 4 la_data_in[58]
port 227 nsew
rlabel metal2 s 337078 -960 337190 480 4 la_data_in[59]
port 228 nsew
rlabel metal2 s 144430 -960 144542 480 4 la_data_in[5]
port 229 nsew
rlabel metal2 s 340666 -960 340778 480 4 la_data_in[60]
port 230 nsew
rlabel metal2 s 344254 -960 344366 480 4 la_data_in[61]
port 231 nsew
rlabel metal2 s 347842 -960 347954 480 4 la_data_in[62]
port 232 nsew
rlabel metal2 s 351338 -960 351450 480 4 la_data_in[63]
port 233 nsew
rlabel metal2 s 354926 -960 355038 480 4 la_data_in[64]
port 234 nsew
rlabel metal2 s 358514 -960 358626 480 4 la_data_in[65]
port 235 nsew
rlabel metal2 s 362102 -960 362214 480 4 la_data_in[66]
port 236 nsew
rlabel metal2 s 365690 -960 365802 480 4 la_data_in[67]
port 237 nsew
rlabel metal2 s 369186 -960 369298 480 4 la_data_in[68]
port 238 nsew
rlabel metal2 s 372774 -960 372886 480 4 la_data_in[69]
port 239 nsew
rlabel metal2 s 148018 -960 148130 480 4 la_data_in[6]
port 240 nsew
rlabel metal2 s 376362 -960 376474 480 4 la_data_in[70]
port 241 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_data_in[71]
port 242 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_data_in[72]
port 243 nsew
rlabel metal2 s 387034 -960 387146 480 4 la_data_in[73]
port 244 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_data_in[74]
port 245 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_data_in[75]
port 246 nsew
rlabel metal2 s 397798 -960 397910 480 4 la_data_in[76]
port 247 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_data_in[77]
port 248 nsew
rlabel metal2 s 404882 -960 404994 480 4 la_data_in[78]
port 249 nsew
rlabel metal2 s 408470 -960 408582 480 4 la_data_in[79]
port 250 nsew
rlabel metal2 s 151514 -960 151626 480 4 la_data_in[7]
port 251 nsew
rlabel metal2 s 412058 -960 412170 480 4 la_data_in[80]
port 252 nsew
rlabel metal2 s 415646 -960 415758 480 4 la_data_in[81]
port 253 nsew
rlabel metal2 s 419142 -960 419254 480 4 la_data_in[82]
port 254 nsew
rlabel metal2 s 422730 -960 422842 480 4 la_data_in[83]
port 255 nsew
rlabel metal2 s 426318 -960 426430 480 4 la_data_in[84]
port 256 nsew
rlabel metal2 s 429906 -960 430018 480 4 la_data_in[85]
port 257 nsew
rlabel metal2 s 433494 -960 433606 480 4 la_data_in[86]
port 258 nsew
rlabel metal2 s 436990 -960 437102 480 4 la_data_in[87]
port 259 nsew
rlabel metal2 s 440578 -960 440690 480 4 la_data_in[88]
port 260 nsew
rlabel metal2 s 444166 -960 444278 480 4 la_data_in[89]
port 261 nsew
rlabel metal2 s 155102 -960 155214 480 4 la_data_in[8]
port 262 nsew
rlabel metal2 s 447754 -960 447866 480 4 la_data_in[90]
port 263 nsew
rlabel metal2 s 451250 -960 451362 480 4 la_data_in[91]
port 264 nsew
rlabel metal2 s 454838 -960 454950 480 4 la_data_in[92]
port 265 nsew
rlabel metal2 s 458426 -960 458538 480 4 la_data_in[93]
port 266 nsew
rlabel metal2 s 462014 -960 462126 480 4 la_data_in[94]
port 267 nsew
rlabel metal2 s 465602 -960 465714 480 4 la_data_in[95]
port 268 nsew
rlabel metal2 s 469098 -960 469210 480 4 la_data_in[96]
port 269 nsew
rlabel metal2 s 472686 -960 472798 480 4 la_data_in[97]
port 270 nsew
rlabel metal2 s 476274 -960 476386 480 4 la_data_in[98]
port 271 nsew
rlabel metal2 s 479862 -960 479974 480 4 la_data_in[99]
port 272 nsew
rlabel metal2 s 158690 -960 158802 480 4 la_data_in[9]
port 273 nsew
rlabel metal2 s 127778 -960 127890 480 4 la_data_out[0]
port 274 nsew
rlabel metal2 s 484554 -960 484666 480 4 la_data_out[100]
port 275 nsew
rlabel metal2 s 488142 -960 488254 480 4 la_data_out[101]
port 276 nsew
rlabel metal2 s 491730 -960 491842 480 4 la_data_out[102]
port 277 nsew
rlabel metal2 s 495318 -960 495430 480 4 la_data_out[103]
port 278 nsew
rlabel metal2 s 498906 -960 499018 480 4 la_data_out[104]
port 279 nsew
rlabel metal2 s 502402 -960 502514 480 4 la_data_out[105]
port 280 nsew
rlabel metal2 s 505990 -960 506102 480 4 la_data_out[106]
port 281 nsew
rlabel metal2 s 509578 -960 509690 480 4 la_data_out[107]
port 282 nsew
rlabel metal2 s 513166 -960 513278 480 4 la_data_out[108]
port 283 nsew
rlabel metal2 s 516754 -960 516866 480 4 la_data_out[109]
port 284 nsew
rlabel metal2 s 163474 -960 163586 480 4 la_data_out[10]
port 285 nsew
rlabel metal2 s 520250 -960 520362 480 4 la_data_out[110]
port 286 nsew
rlabel metal2 s 523838 -960 523950 480 4 la_data_out[111]
port 287 nsew
rlabel metal2 s 527426 -960 527538 480 4 la_data_out[112]
port 288 nsew
rlabel metal2 s 531014 -960 531126 480 4 la_data_out[113]
port 289 nsew
rlabel metal2 s 534510 -960 534622 480 4 la_data_out[114]
port 290 nsew
rlabel metal2 s 538098 -960 538210 480 4 la_data_out[115]
port 291 nsew
rlabel metal2 s 541686 -960 541798 480 4 la_data_out[116]
port 292 nsew
rlabel metal2 s 545274 -960 545386 480 4 la_data_out[117]
port 293 nsew
rlabel metal2 s 548862 -960 548974 480 4 la_data_out[118]
port 294 nsew
rlabel metal2 s 552358 -960 552470 480 4 la_data_out[119]
port 295 nsew
rlabel metal2 s 167062 -960 167174 480 4 la_data_out[11]
port 296 nsew
rlabel metal2 s 555946 -960 556058 480 4 la_data_out[120]
port 297 nsew
rlabel metal2 s 559534 -960 559646 480 4 la_data_out[121]
port 298 nsew
rlabel metal2 s 563122 -960 563234 480 4 la_data_out[122]
port 299 nsew
rlabel metal2 s 566710 -960 566822 480 4 la_data_out[123]
port 300 nsew
rlabel metal2 s 570206 -960 570318 480 4 la_data_out[124]
port 301 nsew
rlabel metal2 s 573794 -960 573906 480 4 la_data_out[125]
port 302 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[126]
port 303 nsew
rlabel metal2 s 580970 -960 581082 480 4 la_data_out[127]
port 304 nsew
rlabel metal2 s 170558 -960 170670 480 4 la_data_out[12]
port 305 nsew
rlabel metal2 s 174146 -960 174258 480 4 la_data_out[13]
port 306 nsew
rlabel metal2 s 177734 -960 177846 480 4 la_data_out[14]
port 307 nsew
rlabel metal2 s 181322 -960 181434 480 4 la_data_out[15]
port 308 nsew
rlabel metal2 s 184818 -960 184930 480 4 la_data_out[16]
port 309 nsew
rlabel metal2 s 188406 -960 188518 480 4 la_data_out[17]
port 310 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_data_out[18]
port 311 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_data_out[19]
port 312 nsew
rlabel metal2 s 131366 -960 131478 480 4 la_data_out[1]
port 313 nsew
rlabel metal2 s 199170 -960 199282 480 4 la_data_out[20]
port 314 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_data_out[21]
port 315 nsew
rlabel metal2 s 206254 -960 206366 480 4 la_data_out[22]
port 316 nsew
rlabel metal2 s 209842 -960 209954 480 4 la_data_out[23]
port 317 nsew
rlabel metal2 s 213430 -960 213542 480 4 la_data_out[24]
port 318 nsew
rlabel metal2 s 217018 -960 217130 480 4 la_data_out[25]
port 319 nsew
rlabel metal2 s 220514 -960 220626 480 4 la_data_out[26]
port 320 nsew
rlabel metal2 s 224102 -960 224214 480 4 la_data_out[27]
port 321 nsew
rlabel metal2 s 227690 -960 227802 480 4 la_data_out[28]
port 322 nsew
rlabel metal2 s 231278 -960 231390 480 4 la_data_out[29]
port 323 nsew
rlabel metal2 s 134862 -960 134974 480 4 la_data_out[2]
port 324 nsew
rlabel metal2 s 234774 -960 234886 480 4 la_data_out[30]
port 325 nsew
rlabel metal2 s 238362 -960 238474 480 4 la_data_out[31]
port 326 nsew
rlabel metal2 s 241950 -960 242062 480 4 la_data_out[32]
port 327 nsew
rlabel metal2 s 245538 -960 245650 480 4 la_data_out[33]
port 328 nsew
rlabel metal2 s 249126 -960 249238 480 4 la_data_out[34]
port 329 nsew
rlabel metal2 s 252622 -960 252734 480 4 la_data_out[35]
port 330 nsew
rlabel metal2 s 256210 -960 256322 480 4 la_data_out[36]
port 331 nsew
rlabel metal2 s 259798 -960 259910 480 4 la_data_out[37]
port 332 nsew
rlabel metal2 s 263386 -960 263498 480 4 la_data_out[38]
port 333 nsew
rlabel metal2 s 266974 -960 267086 480 4 la_data_out[39]
port 334 nsew
rlabel metal2 s 138450 -960 138562 480 4 la_data_out[3]
port 335 nsew
rlabel metal2 s 270470 -960 270582 480 4 la_data_out[40]
port 336 nsew
rlabel metal2 s 274058 -960 274170 480 4 la_data_out[41]
port 337 nsew
rlabel metal2 s 277646 -960 277758 480 4 la_data_out[42]
port 338 nsew
rlabel metal2 s 281234 -960 281346 480 4 la_data_out[43]
port 339 nsew
rlabel metal2 s 284730 -960 284842 480 4 la_data_out[44]
port 340 nsew
rlabel metal2 s 288318 -960 288430 480 4 la_data_out[45]
port 341 nsew
rlabel metal2 s 291906 -960 292018 480 4 la_data_out[46]
port 342 nsew
rlabel metal2 s 295494 -960 295606 480 4 la_data_out[47]
port 343 nsew
rlabel metal2 s 299082 -960 299194 480 4 la_data_out[48]
port 344 nsew
rlabel metal2 s 302578 -960 302690 480 4 la_data_out[49]
port 345 nsew
rlabel metal2 s 142038 -960 142150 480 4 la_data_out[4]
port 346 nsew
rlabel metal2 s 306166 -960 306278 480 4 la_data_out[50]
port 347 nsew
rlabel metal2 s 309754 -960 309866 480 4 la_data_out[51]
port 348 nsew
rlabel metal2 s 313342 -960 313454 480 4 la_data_out[52]
port 349 nsew
rlabel metal2 s 316930 -960 317042 480 4 la_data_out[53]
port 350 nsew
rlabel metal2 s 320426 -960 320538 480 4 la_data_out[54]
port 351 nsew
rlabel metal2 s 324014 -960 324126 480 4 la_data_out[55]
port 352 nsew
rlabel metal2 s 327602 -960 327714 480 4 la_data_out[56]
port 353 nsew
rlabel metal2 s 331190 -960 331302 480 4 la_data_out[57]
port 354 nsew
rlabel metal2 s 334686 -960 334798 480 4 la_data_out[58]
port 355 nsew
rlabel metal2 s 338274 -960 338386 480 4 la_data_out[59]
port 356 nsew
rlabel metal2 s 145626 -960 145738 480 4 la_data_out[5]
port 357 nsew
rlabel metal2 s 341862 -960 341974 480 4 la_data_out[60]
port 358 nsew
rlabel metal2 s 345450 -960 345562 480 4 la_data_out[61]
port 359 nsew
rlabel metal2 s 349038 -960 349150 480 4 la_data_out[62]
port 360 nsew
rlabel metal2 s 352534 -960 352646 480 4 la_data_out[63]
port 361 nsew
rlabel metal2 s 356122 -960 356234 480 4 la_data_out[64]
port 362 nsew
rlabel metal2 s 359710 -960 359822 480 4 la_data_out[65]
port 363 nsew
rlabel metal2 s 363298 -960 363410 480 4 la_data_out[66]
port 364 nsew
rlabel metal2 s 366886 -960 366998 480 4 la_data_out[67]
port 365 nsew
rlabel metal2 s 370382 -960 370494 480 4 la_data_out[68]
port 366 nsew
rlabel metal2 s 373970 -960 374082 480 4 la_data_out[69]
port 367 nsew
rlabel metal2 s 149214 -960 149326 480 4 la_data_out[6]
port 368 nsew
rlabel metal2 s 377558 -960 377670 480 4 la_data_out[70]
port 369 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_out[71]
port 370 nsew
rlabel metal2 s 384642 -960 384754 480 4 la_data_out[72]
port 371 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_out[73]
port 372 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_out[74]
port 373 nsew
rlabel metal2 s 395406 -960 395518 480 4 la_data_out[75]
port 374 nsew
rlabel metal2 s 398994 -960 399106 480 4 la_data_out[76]
port 375 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_out[77]
port 376 nsew
rlabel metal2 s 406078 -960 406190 480 4 la_data_out[78]
port 377 nsew
rlabel metal2 s 409666 -960 409778 480 4 la_data_out[79]
port 378 nsew
rlabel metal2 s 152710 -960 152822 480 4 la_data_out[7]
port 379 nsew
rlabel metal2 s 413254 -960 413366 480 4 la_data_out[80]
port 380 nsew
rlabel metal2 s 416842 -960 416954 480 4 la_data_out[81]
port 381 nsew
rlabel metal2 s 420338 -960 420450 480 4 la_data_out[82]
port 382 nsew
rlabel metal2 s 423926 -960 424038 480 4 la_data_out[83]
port 383 nsew
rlabel metal2 s 427514 -960 427626 480 4 la_data_out[84]
port 384 nsew
rlabel metal2 s 431102 -960 431214 480 4 la_data_out[85]
port 385 nsew
rlabel metal2 s 434598 -960 434710 480 4 la_data_out[86]
port 386 nsew
rlabel metal2 s 438186 -960 438298 480 4 la_data_out[87]
port 387 nsew
rlabel metal2 s 441774 -960 441886 480 4 la_data_out[88]
port 388 nsew
rlabel metal2 s 445362 -960 445474 480 4 la_data_out[89]
port 389 nsew
rlabel metal2 s 156298 -960 156410 480 4 la_data_out[8]
port 390 nsew
rlabel metal2 s 448950 -960 449062 480 4 la_data_out[90]
port 391 nsew
rlabel metal2 s 452446 -960 452558 480 4 la_data_out[91]
port 392 nsew
rlabel metal2 s 456034 -960 456146 480 4 la_data_out[92]
port 393 nsew
rlabel metal2 s 459622 -960 459734 480 4 la_data_out[93]
port 394 nsew
rlabel metal2 s 463210 -960 463322 480 4 la_data_out[94]
port 395 nsew
rlabel metal2 s 466798 -960 466910 480 4 la_data_out[95]
port 396 nsew
rlabel metal2 s 470294 -960 470406 480 4 la_data_out[96]
port 397 nsew
rlabel metal2 s 473882 -960 473994 480 4 la_data_out[97]
port 398 nsew
rlabel metal2 s 477470 -960 477582 480 4 la_data_out[98]
port 399 nsew
rlabel metal2 s 481058 -960 481170 480 4 la_data_out[99]
port 400 nsew
rlabel metal2 s 159886 -960 159998 480 4 la_data_out[9]
port 401 nsew
rlabel metal2 s 128974 -960 129086 480 4 la_oen[0]
port 402 nsew
rlabel metal2 s 485750 -960 485862 480 4 la_oen[100]
port 403 nsew
rlabel metal2 s 489338 -960 489450 480 4 la_oen[101]
port 404 nsew
rlabel metal2 s 492926 -960 493038 480 4 la_oen[102]
port 405 nsew
rlabel metal2 s 496514 -960 496626 480 4 la_oen[103]
port 406 nsew
rlabel metal2 s 500102 -960 500214 480 4 la_oen[104]
port 407 nsew
rlabel metal2 s 503598 -960 503710 480 4 la_oen[105]
port 408 nsew
rlabel metal2 s 507186 -960 507298 480 4 la_oen[106]
port 409 nsew
rlabel metal2 s 510774 -960 510886 480 4 la_oen[107]
port 410 nsew
rlabel metal2 s 514362 -960 514474 480 4 la_oen[108]
port 411 nsew
rlabel metal2 s 517858 -960 517970 480 4 la_oen[109]
port 412 nsew
rlabel metal2 s 164670 -960 164782 480 4 la_oen[10]
port 413 nsew
rlabel metal2 s 521446 -960 521558 480 4 la_oen[110]
port 414 nsew
rlabel metal2 s 525034 -960 525146 480 4 la_oen[111]
port 415 nsew
rlabel metal2 s 528622 -960 528734 480 4 la_oen[112]
port 416 nsew
rlabel metal2 s 532210 -960 532322 480 4 la_oen[113]
port 417 nsew
rlabel metal2 s 535706 -960 535818 480 4 la_oen[114]
port 418 nsew
rlabel metal2 s 539294 -960 539406 480 4 la_oen[115]
port 419 nsew
rlabel metal2 s 542882 -960 542994 480 4 la_oen[116]
port 420 nsew
rlabel metal2 s 546470 -960 546582 480 4 la_oen[117]
port 421 nsew
rlabel metal2 s 550058 -960 550170 480 4 la_oen[118]
port 422 nsew
rlabel metal2 s 553554 -960 553666 480 4 la_oen[119]
port 423 nsew
rlabel metal2 s 168166 -960 168278 480 4 la_oen[11]
port 424 nsew
rlabel metal2 s 557142 -960 557254 480 4 la_oen[120]
port 425 nsew
rlabel metal2 s 560730 -960 560842 480 4 la_oen[121]
port 426 nsew
rlabel metal2 s 564318 -960 564430 480 4 la_oen[122]
port 427 nsew
rlabel metal2 s 567814 -960 567926 480 4 la_oen[123]
port 428 nsew
rlabel metal2 s 571402 -960 571514 480 4 la_oen[124]
port 429 nsew
rlabel metal2 s 574990 -960 575102 480 4 la_oen[125]
port 430 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oen[126]
port 431 nsew
rlabel metal2 s 582166 -960 582278 480 4 la_oen[127]
port 432 nsew
rlabel metal2 s 171754 -960 171866 480 4 la_oen[12]
port 433 nsew
rlabel metal2 s 175342 -960 175454 480 4 la_oen[13]
port 434 nsew
rlabel metal2 s 178930 -960 179042 480 4 la_oen[14]
port 435 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_oen[15]
port 436 nsew
rlabel metal2 s 186014 -960 186126 480 4 la_oen[16]
port 437 nsew
rlabel metal2 s 189602 -960 189714 480 4 la_oen[17]
port 438 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_oen[18]
port 439 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_oen[19]
port 440 nsew
rlabel metal2 s 132562 -960 132674 480 4 la_oen[1]
port 441 nsew
rlabel metal2 s 200366 -960 200478 480 4 la_oen[20]
port 442 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_oen[21]
port 443 nsew
rlabel metal2 s 207450 -960 207562 480 4 la_oen[22]
port 444 nsew
rlabel metal2 s 211038 -960 211150 480 4 la_oen[23]
port 445 nsew
rlabel metal2 s 214626 -960 214738 480 4 la_oen[24]
port 446 nsew
rlabel metal2 s 218122 -960 218234 480 4 la_oen[25]
port 447 nsew
rlabel metal2 s 221710 -960 221822 480 4 la_oen[26]
port 448 nsew
rlabel metal2 s 225298 -960 225410 480 4 la_oen[27]
port 449 nsew
rlabel metal2 s 228886 -960 228998 480 4 la_oen[28]
port 450 nsew
rlabel metal2 s 232474 -960 232586 480 4 la_oen[29]
port 451 nsew
rlabel metal2 s 136058 -960 136170 480 4 la_oen[2]
port 452 nsew
rlabel metal2 s 235970 -960 236082 480 4 la_oen[30]
port 453 nsew
rlabel metal2 s 239558 -960 239670 480 4 la_oen[31]
port 454 nsew
rlabel metal2 s 243146 -960 243258 480 4 la_oen[32]
port 455 nsew
rlabel metal2 s 246734 -960 246846 480 4 la_oen[33]
port 456 nsew
rlabel metal2 s 250322 -960 250434 480 4 la_oen[34]
port 457 nsew
rlabel metal2 s 253818 -960 253930 480 4 la_oen[35]
port 458 nsew
rlabel metal2 s 257406 -960 257518 480 4 la_oen[36]
port 459 nsew
rlabel metal2 s 260994 -960 261106 480 4 la_oen[37]
port 460 nsew
rlabel metal2 s 264582 -960 264694 480 4 la_oen[38]
port 461 nsew
rlabel metal2 s 268078 -960 268190 480 4 la_oen[39]
port 462 nsew
rlabel metal2 s 139646 -960 139758 480 4 la_oen[3]
port 463 nsew
rlabel metal2 s 271666 -960 271778 480 4 la_oen[40]
port 464 nsew
rlabel metal2 s 275254 -960 275366 480 4 la_oen[41]
port 465 nsew
rlabel metal2 s 278842 -960 278954 480 4 la_oen[42]
port 466 nsew
rlabel metal2 s 282430 -960 282542 480 4 la_oen[43]
port 467 nsew
rlabel metal2 s 285926 -960 286038 480 4 la_oen[44]
port 468 nsew
rlabel metal2 s 289514 -960 289626 480 4 la_oen[45]
port 469 nsew
rlabel metal2 s 293102 -960 293214 480 4 la_oen[46]
port 470 nsew
rlabel metal2 s 296690 -960 296802 480 4 la_oen[47]
port 471 nsew
rlabel metal2 s 300278 -960 300390 480 4 la_oen[48]
port 472 nsew
rlabel metal2 s 303774 -960 303886 480 4 la_oen[49]
port 473 nsew
rlabel metal2 s 143234 -960 143346 480 4 la_oen[4]
port 474 nsew
rlabel metal2 s 307362 -960 307474 480 4 la_oen[50]
port 475 nsew
rlabel metal2 s 310950 -960 311062 480 4 la_oen[51]
port 476 nsew
rlabel metal2 s 314538 -960 314650 480 4 la_oen[52]
port 477 nsew
rlabel metal2 s 318034 -960 318146 480 4 la_oen[53]
port 478 nsew
rlabel metal2 s 321622 -960 321734 480 4 la_oen[54]
port 479 nsew
rlabel metal2 s 325210 -960 325322 480 4 la_oen[55]
port 480 nsew
rlabel metal2 s 328798 -960 328910 480 4 la_oen[56]
port 481 nsew
rlabel metal2 s 332386 -960 332498 480 4 la_oen[57]
port 482 nsew
rlabel metal2 s 335882 -960 335994 480 4 la_oen[58]
port 483 nsew
rlabel metal2 s 339470 -960 339582 480 4 la_oen[59]
port 484 nsew
rlabel metal2 s 146822 -960 146934 480 4 la_oen[5]
port 485 nsew
rlabel metal2 s 343058 -960 343170 480 4 la_oen[60]
port 486 nsew
rlabel metal2 s 346646 -960 346758 480 4 la_oen[61]
port 487 nsew
rlabel metal2 s 350234 -960 350346 480 4 la_oen[62]
port 488 nsew
rlabel metal2 s 353730 -960 353842 480 4 la_oen[63]
port 489 nsew
rlabel metal2 s 357318 -960 357430 480 4 la_oen[64]
port 490 nsew
rlabel metal2 s 360906 -960 361018 480 4 la_oen[65]
port 491 nsew
rlabel metal2 s 364494 -960 364606 480 4 la_oen[66]
port 492 nsew
rlabel metal2 s 367990 -960 368102 480 4 la_oen[67]
port 493 nsew
rlabel metal2 s 371578 -960 371690 480 4 la_oen[68]
port 494 nsew
rlabel metal2 s 375166 -960 375278 480 4 la_oen[69]
port 495 nsew
rlabel metal2 s 150410 -960 150522 480 4 la_oen[6]
port 496 nsew
rlabel metal2 s 378754 -960 378866 480 4 la_oen[70]
port 497 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_oen[71]
port 498 nsew
rlabel metal2 s 385838 -960 385950 480 4 la_oen[72]
port 499 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_oen[73]
port 500 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_oen[74]
port 501 nsew
rlabel metal2 s 396602 -960 396714 480 4 la_oen[75]
port 502 nsew
rlabel metal2 s 400190 -960 400302 480 4 la_oen[76]
port 503 nsew
rlabel metal2 s 403686 -960 403798 480 4 la_oen[77]
port 504 nsew
rlabel metal2 s 407274 -960 407386 480 4 la_oen[78]
port 505 nsew
rlabel metal2 s 410862 -960 410974 480 4 la_oen[79]
port 506 nsew
rlabel metal2 s 153906 -960 154018 480 4 la_oen[7]
port 507 nsew
rlabel metal2 s 414450 -960 414562 480 4 la_oen[80]
port 508 nsew
rlabel metal2 s 417946 -960 418058 480 4 la_oen[81]
port 509 nsew
rlabel metal2 s 421534 -960 421646 480 4 la_oen[82]
port 510 nsew
rlabel metal2 s 425122 -960 425234 480 4 la_oen[83]
port 511 nsew
rlabel metal2 s 428710 -960 428822 480 4 la_oen[84]
port 512 nsew
rlabel metal2 s 432298 -960 432410 480 4 la_oen[85]
port 513 nsew
rlabel metal2 s 435794 -960 435906 480 4 la_oen[86]
port 514 nsew
rlabel metal2 s 439382 -960 439494 480 4 la_oen[87]
port 515 nsew
rlabel metal2 s 442970 -960 443082 480 4 la_oen[88]
port 516 nsew
rlabel metal2 s 446558 -960 446670 480 4 la_oen[89]
port 517 nsew
rlabel metal2 s 157494 -960 157606 480 4 la_oen[8]
port 518 nsew
rlabel metal2 s 450146 -960 450258 480 4 la_oen[90]
port 519 nsew
rlabel metal2 s 453642 -960 453754 480 4 la_oen[91]
port 520 nsew
rlabel metal2 s 457230 -960 457342 480 4 la_oen[92]
port 521 nsew
rlabel metal2 s 460818 -960 460930 480 4 la_oen[93]
port 522 nsew
rlabel metal2 s 464406 -960 464518 480 4 la_oen[94]
port 523 nsew
rlabel metal2 s 467902 -960 468014 480 4 la_oen[95]
port 524 nsew
rlabel metal2 s 471490 -960 471602 480 4 la_oen[96]
port 525 nsew
rlabel metal2 s 475078 -960 475190 480 4 la_oen[97]
port 526 nsew
rlabel metal2 s 478666 -960 478778 480 4 la_oen[98]
port 527 nsew
rlabel metal2 s 482254 -960 482366 480 4 la_oen[99]
port 528 nsew
rlabel metal2 s 161082 -960 161194 480 4 la_oen[9]
port 529 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_clock2
port 530 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 531 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 532 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 533 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 534 nsew
rlabel metal2 s 48106 -960 48218 480 4 wbs_adr_i[10]
port 535 nsew
rlabel metal2 s 51602 -960 51714 480 4 wbs_adr_i[11]
port 536 nsew
rlabel metal2 s 55190 -960 55302 480 4 wbs_adr_i[12]
port 537 nsew
rlabel metal2 s 58778 -960 58890 480 4 wbs_adr_i[13]
port 538 nsew
rlabel metal2 s 62366 -960 62478 480 4 wbs_adr_i[14]
port 539 nsew
rlabel metal2 s 65954 -960 66066 480 4 wbs_adr_i[15]
port 540 nsew
rlabel metal2 s 69450 -960 69562 480 4 wbs_adr_i[16]
port 541 nsew
rlabel metal2 s 73038 -960 73150 480 4 wbs_adr_i[17]
port 542 nsew
rlabel metal2 s 76626 -960 76738 480 4 wbs_adr_i[18]
port 543 nsew
rlabel metal2 s 80214 -960 80326 480 4 wbs_adr_i[19]
port 544 nsew
rlabel metal2 s 12410 -960 12522 480 4 wbs_adr_i[1]
port 545 nsew
rlabel metal2 s 83802 -960 83914 480 4 wbs_adr_i[20]
port 546 nsew
rlabel metal2 s 87298 -960 87410 480 4 wbs_adr_i[21]
port 547 nsew
rlabel metal2 s 90886 -960 90998 480 4 wbs_adr_i[22]
port 548 nsew
rlabel metal2 s 94474 -960 94586 480 4 wbs_adr_i[23]
port 549 nsew
rlabel metal2 s 98062 -960 98174 480 4 wbs_adr_i[24]
port 550 nsew
rlabel metal2 s 101558 -960 101670 480 4 wbs_adr_i[25]
port 551 nsew
rlabel metal2 s 105146 -960 105258 480 4 wbs_adr_i[26]
port 552 nsew
rlabel metal2 s 108734 -960 108846 480 4 wbs_adr_i[27]
port 553 nsew
rlabel metal2 s 112322 -960 112434 480 4 wbs_adr_i[28]
port 554 nsew
rlabel metal2 s 115910 -960 116022 480 4 wbs_adr_i[29]
port 555 nsew
rlabel metal2 s 17194 -960 17306 480 4 wbs_adr_i[2]
port 556 nsew
rlabel metal2 s 119406 -960 119518 480 4 wbs_adr_i[30]
port 557 nsew
rlabel metal2 s 122994 -960 123106 480 4 wbs_adr_i[31]
port 558 nsew
rlabel metal2 s 21886 -960 21998 480 4 wbs_adr_i[3]
port 559 nsew
rlabel metal2 s 26670 -960 26782 480 4 wbs_adr_i[4]
port 560 nsew
rlabel metal2 s 30258 -960 30370 480 4 wbs_adr_i[5]
port 561 nsew
rlabel metal2 s 33846 -960 33958 480 4 wbs_adr_i[6]
port 562 nsew
rlabel metal2 s 37342 -960 37454 480 4 wbs_adr_i[7]
port 563 nsew
rlabel metal2 s 40930 -960 41042 480 4 wbs_adr_i[8]
port 564 nsew
rlabel metal2 s 44518 -960 44630 480 4 wbs_adr_i[9]
port 565 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 566 nsew
rlabel metal2 s 8822 -960 8934 480 4 wbs_dat_i[0]
port 567 nsew
rlabel metal2 s 49302 -960 49414 480 4 wbs_dat_i[10]
port 568 nsew
rlabel metal2 s 52798 -960 52910 480 4 wbs_dat_i[11]
port 569 nsew
rlabel metal2 s 56386 -960 56498 480 4 wbs_dat_i[12]
port 570 nsew
rlabel metal2 s 59974 -960 60086 480 4 wbs_dat_i[13]
port 571 nsew
rlabel metal2 s 63562 -960 63674 480 4 wbs_dat_i[14]
port 572 nsew
rlabel metal2 s 67150 -960 67262 480 4 wbs_dat_i[15]
port 573 nsew
rlabel metal2 s 70646 -960 70758 480 4 wbs_dat_i[16]
port 574 nsew
rlabel metal2 s 74234 -960 74346 480 4 wbs_dat_i[17]
port 575 nsew
rlabel metal2 s 77822 -960 77934 480 4 wbs_dat_i[18]
port 576 nsew
rlabel metal2 s 81410 -960 81522 480 4 wbs_dat_i[19]
port 577 nsew
rlabel metal2 s 13606 -960 13718 480 4 wbs_dat_i[1]
port 578 nsew
rlabel metal2 s 84906 -960 85018 480 4 wbs_dat_i[20]
port 579 nsew
rlabel metal2 s 88494 -960 88606 480 4 wbs_dat_i[21]
port 580 nsew
rlabel metal2 s 92082 -960 92194 480 4 wbs_dat_i[22]
port 581 nsew
rlabel metal2 s 95670 -960 95782 480 4 wbs_dat_i[23]
port 582 nsew
rlabel metal2 s 99258 -960 99370 480 4 wbs_dat_i[24]
port 583 nsew
rlabel metal2 s 102754 -960 102866 480 4 wbs_dat_i[25]
port 584 nsew
rlabel metal2 s 106342 -960 106454 480 4 wbs_dat_i[26]
port 585 nsew
rlabel metal2 s 109930 -960 110042 480 4 wbs_dat_i[27]
port 586 nsew
rlabel metal2 s 113518 -960 113630 480 4 wbs_dat_i[28]
port 587 nsew
rlabel metal2 s 117106 -960 117218 480 4 wbs_dat_i[29]
port 588 nsew
rlabel metal2 s 18298 -960 18410 480 4 wbs_dat_i[2]
port 589 nsew
rlabel metal2 s 120602 -960 120714 480 4 wbs_dat_i[30]
port 590 nsew
rlabel metal2 s 124190 -960 124302 480 4 wbs_dat_i[31]
port 591 nsew
rlabel metal2 s 23082 -960 23194 480 4 wbs_dat_i[3]
port 592 nsew
rlabel metal2 s 27866 -960 27978 480 4 wbs_dat_i[4]
port 593 nsew
rlabel metal2 s 31454 -960 31566 480 4 wbs_dat_i[5]
port 594 nsew
rlabel metal2 s 34950 -960 35062 480 4 wbs_dat_i[6]
port 595 nsew
rlabel metal2 s 38538 -960 38650 480 4 wbs_dat_i[7]
port 596 nsew
rlabel metal2 s 42126 -960 42238 480 4 wbs_dat_i[8]
port 597 nsew
rlabel metal2 s 45714 -960 45826 480 4 wbs_dat_i[9]
port 598 nsew
rlabel metal2 s 10018 -960 10130 480 4 wbs_dat_o[0]
port 599 nsew
rlabel metal2 s 50498 -960 50610 480 4 wbs_dat_o[10]
port 600 nsew
rlabel metal2 s 53994 -960 54106 480 4 wbs_dat_o[11]
port 601 nsew
rlabel metal2 s 57582 -960 57694 480 4 wbs_dat_o[12]
port 602 nsew
rlabel metal2 s 61170 -960 61282 480 4 wbs_dat_o[13]
port 603 nsew
rlabel metal2 s 64758 -960 64870 480 4 wbs_dat_o[14]
port 604 nsew
rlabel metal2 s 68254 -960 68366 480 4 wbs_dat_o[15]
port 605 nsew
rlabel metal2 s 71842 -960 71954 480 4 wbs_dat_o[16]
port 606 nsew
rlabel metal2 s 75430 -960 75542 480 4 wbs_dat_o[17]
port 607 nsew
rlabel metal2 s 79018 -960 79130 480 4 wbs_dat_o[18]
port 608 nsew
rlabel metal2 s 82606 -960 82718 480 4 wbs_dat_o[19]
port 609 nsew
rlabel metal2 s 14802 -960 14914 480 4 wbs_dat_o[1]
port 610 nsew
rlabel metal2 s 86102 -960 86214 480 4 wbs_dat_o[20]
port 611 nsew
rlabel metal2 s 89690 -960 89802 480 4 wbs_dat_o[21]
port 612 nsew
rlabel metal2 s 93278 -960 93390 480 4 wbs_dat_o[22]
port 613 nsew
rlabel metal2 s 96866 -960 96978 480 4 wbs_dat_o[23]
port 614 nsew
rlabel metal2 s 100454 -960 100566 480 4 wbs_dat_o[24]
port 615 nsew
rlabel metal2 s 103950 -960 104062 480 4 wbs_dat_o[25]
port 616 nsew
rlabel metal2 s 107538 -960 107650 480 4 wbs_dat_o[26]
port 617 nsew
rlabel metal2 s 111126 -960 111238 480 4 wbs_dat_o[27]
port 618 nsew
rlabel metal2 s 114714 -960 114826 480 4 wbs_dat_o[28]
port 619 nsew
rlabel metal2 s 118210 -960 118322 480 4 wbs_dat_o[29]
port 620 nsew
rlabel metal2 s 19494 -960 19606 480 4 wbs_dat_o[2]
port 621 nsew
rlabel metal2 s 121798 -960 121910 480 4 wbs_dat_o[30]
port 622 nsew
rlabel metal2 s 125386 -960 125498 480 4 wbs_dat_o[31]
port 623 nsew
rlabel metal2 s 24278 -960 24390 480 4 wbs_dat_o[3]
port 624 nsew
rlabel metal2 s 29062 -960 29174 480 4 wbs_dat_o[4]
port 625 nsew
rlabel metal2 s 32650 -960 32762 480 4 wbs_dat_o[5]
port 626 nsew
rlabel metal2 s 36146 -960 36258 480 4 wbs_dat_o[6]
port 627 nsew
rlabel metal2 s 39734 -960 39846 480 4 wbs_dat_o[7]
port 628 nsew
rlabel metal2 s 43322 -960 43434 480 4 wbs_dat_o[8]
port 629 nsew
rlabel metal2 s 46910 -960 47022 480 4 wbs_dat_o[9]
port 630 nsew
rlabel metal2 s 11214 -960 11326 480 4 wbs_sel_i[0]
port 631 nsew
rlabel metal2 s 15998 -960 16110 480 4 wbs_sel_i[1]
port 632 nsew
rlabel metal2 s 20690 -960 20802 480 4 wbs_sel_i[2]
port 633 nsew
rlabel metal2 s 25474 -960 25586 480 4 wbs_sel_i[3]
port 634 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 635 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 636 nsew
rlabel metal5 s -1996 -924 585920 -324 4 vccd1
port 637 nsew
rlabel metal5 s -2916 -1844 586840 -1244 4 vssd1
port 638 nsew
rlabel metal5 s -3836 -2764 587760 -2164 4 vccd2
port 639 nsew
rlabel metal5 s -4756 -3684 588680 -3084 4 vssd2
port 640 nsew
rlabel metal5 s -5676 -4604 589600 -4004 4 vdda1
port 641 nsew
rlabel metal5 s -6596 -5524 590520 -4924 4 vssa1
port 642 nsew
rlabel metal5 s -7516 -6444 591440 -5844 4 vdda2
port 643 nsew
rlabel metal5 s -8436 -7364 592360 -6764 4 vssa2
port 644 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
