magic
tech sky130A
timestamp 1607536219
<< metal1 >>
rect 2106 8299 2213 8307
rect 2106 8285 2216 8299
rect 2189 5985 2216 8285
rect 1907 5965 2216 5985
rect 1907 5946 1958 5965
rect 2027 5485 2195 5504
rect 2166 3258 2195 5485
rect 2103 3236 2195 3258
rect 2166 3230 2195 3236
<< metal2 >>
rect 283 8377 1390 8403
rect 269 5938 296 6176
rect 269 5914 1501 5938
rect 269 5533 296 5914
rect 278 3327 1382 3351
<< metal3 >>
rect 1837 8263 1876 10360
rect 1154 8251 1876 8263
rect 1154 8216 1884 8251
rect 132 5537 170 6010
rect 935 5533 970 6805
rect 1593 6055 1631 7237
rect 1107 6054 1650 6055
rect 1100 6013 1650 6054
rect 1840 6040 1884 8216
rect 1100 5859 1144 6013
rect 1840 5981 1883 6040
rect 1195 5974 1883 5981
rect 1186 5947 1883 5974
rect 1186 5942 1858 5947
rect 1103 5390 1142 5859
rect 1186 5464 1220 5942
rect 1186 5427 1881 5464
rect 1192 5420 1881 5427
rect 1101 5375 1360 5390
rect 1837 5378 1878 5420
rect 1101 5356 1364 5375
rect 1329 5317 1364 5356
rect 1837 5347 1884 5378
rect 1322 5283 1640 5317
rect 1840 3211 1884 5347
rect 1148 3167 1884 3211
rect 1148 3164 1870 3167
<< metal4 >>
rect 479 5545 521 5732
rect 479 5506 1641 5545
rect 479 5503 521 5506
rect 516 2943 1528 2982
use Sw-1  Sw-1_0
timestamp 1607536219
transform 1 0 1336 0 1 5441
box -70 45 891 509
use 4good  4good_0
timestamp 1607536219
transform 1 0 48 0 1 614
box -1 2 2115 5105
use 4good  4good_1
timestamp 1607536219
transform 1 0 48 0 1 5663
box -1 2 2115 5105
<< end >>
