magic
tech sky130A
magscale 1 2
timestamp 1606237748
<< nwell >>
rect -111 -127 135 91
<< pmos >>
rect -11 -33 73 -3
<< pdiff >>
rect -11 43 73 55
rect -11 9 1 43
rect 61 9 73 43
rect -11 -3 73 9
rect -11 -45 73 -33
rect -11 -79 1 -45
rect 61 -79 73 -45
rect -11 -91 73 -79
<< pdiffc >>
rect 1 9 61 43
rect 1 -79 61 -45
<< poly >>
rect -108 -1 -42 15
rect -108 -35 -92 -1
rect -58 -3 -42 -1
rect -58 -33 -11 -3
rect 73 -33 99 -3
rect -58 -35 -42 -33
rect -108 -51 -42 -35
<< polycont >>
rect -92 -35 -58 -1
<< locali >>
rect -92 -1 -58 15
rect -15 9 1 43
rect 61 9 77 43
rect -92 -51 -58 -35
rect -15 -79 1 -45
rect 61 -79 77 -45
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.42 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
