magic
tech sky130A
magscale 1 2
timestamp 1608024784
<< dnwell >>
rect -430 -464 2462 2352
<< nwell >>
rect -510 2146 2542 2628
rect -510 -258 -224 2146
rect 2256 -258 2542 2146
rect -510 -544 2542 -258
<< nsubdiff >>
rect -300 2452 2284 2492
rect -300 2406 -254 2452
rect -198 2406 58 2452
rect 114 2406 370 2452
rect 426 2406 682 2452
rect 738 2406 994 2452
rect 1050 2406 1306 2452
rect 1362 2406 1618 2452
rect 1674 2406 1930 2452
rect 1986 2406 2284 2452
rect -300 2368 2284 2406
<< nsubdiffcont >>
rect -254 2406 -198 2452
rect 58 2406 114 2452
rect 370 2406 426 2452
rect 682 2406 738 2452
rect 994 2406 1050 2452
rect 1306 2406 1362 2452
rect 1618 2406 1674 2452
rect 1930 2406 1986 2452
<< locali >>
rect -349 2452 2070 2472
rect -349 2406 -254 2452
rect -198 2406 58 2452
rect 114 2406 370 2452
rect 426 2406 682 2452
rect 738 2406 994 2452
rect 1050 2406 1306 2452
rect 1362 2406 1618 2452
rect 1674 2406 1930 2452
rect 1986 2406 2070 2452
rect -349 2390 2070 2406
<< viali >>
rect -431 2390 -349 2472
<< metal1 >>
rect -437 2472 -343 2484
rect -925 2390 -431 2472
rect -349 2390 -343 2472
rect -437 2378 -343 2390
rect -968 1544 2980 1596
rect -956 1304 2992 1356
rect -938 490 3024 542
<< metal2 >>
rect 384 -840 436 2960
rect 776 -840 828 2974
rect 1156 -848 1208 2996
rect 1548 -870 1600 2996
use 1T-cell  1T-cell_0
array 0 1 772 0 1 814
timestamp 1606190511
transform 1 0 182 0 1 142
box -182 -142 1044 1024
<< labels >>
flabel metal1 -922 1320 -898 1338 0 FreeSans 800 0 0 0 WL0
port 0 nsew
flabel metal1 -918 508 -894 526 0 FreeSans 800 0 0 0 WL1
port 1 nsew
flabel metal2 396 2808 420 2826 0 FreeSans 800 0 0 0 BL0
port 2 nsew
flabel metal2 788 2628 812 2646 0 FreeSans 800 0 0 0 SL0
port 3 nsew
flabel metal2 1172 2834 1196 2852 0 FreeSans 800 0 0 0 BL1
port 4 nsew
flabel metal2 1558 2656 1582 2674 0 FreeSans 800 0 0 0 SL1
port 5 nsew
flabel metal1 -926 1556 -902 1574 0 FreeSans 800 0 0 0 body
port 7 nsew
flabel metal1 -898 2418 -856 2452 0 FreeSans 800 0 0 0 nwell
port 8 nsew
<< end >>
