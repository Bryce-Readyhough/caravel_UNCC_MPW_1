magic
tech sky130A
timestamp 1604306825
<< nmos >>
rect -20 -21 20 21
<< ndiff >>
rect -49 15 -20 21
rect -49 -15 -43 15
rect -26 -15 -20 15
rect -49 -21 -20 -15
rect 20 15 49 21
rect 20 -15 26 15
rect 43 -15 49 15
rect 20 -21 49 -15
<< ndiffc >>
rect -43 -15 -26 15
rect 26 -15 43 15
<< poly >>
rect -20 21 20 34
rect -20 -34 20 -21
<< locali >>
rect -43 15 -26 23
rect -43 -23 -26 -15
rect 26 15 43 23
rect 26 -23 43 -15
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 0.420 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0
string library sky130
<< end >>
