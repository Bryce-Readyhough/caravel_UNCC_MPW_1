magic
tech sky130A
magscale 1 2
timestamp 1606278851
<< locali >>
rect -280 8384 785 8444
rect -1000 8122 -482 8173
rect -280 7850 -220 8384
rect -1846 7720 -1232 7836
rect -964 7758 -505 7800
rect -425 7790 -220 7850
rect -262 2561 780 2621
rect -1025 2408 -547 2465
rect -1828 2018 -1256 2134
rect -262 2125 -202 2561
rect -980 2052 -582 2094
rect -502 2065 -202 2125
rect 19170 1011 19736 1051
rect 17885 447 18174 497
rect 19254 -755 20028 -715
rect 17851 -1291 18174 -1241
rect 19198 -2585 20536 -2545
rect 17945 -3117 18172 -3067
rect 19172 -4399 21036 -4359
rect 17807 -4935 18172 -4885
<< viali >>
rect -1962 7720 -1846 7836
rect -1944 2018 -1828 2134
rect 19736 1011 19776 1051
rect 17835 447 17885 497
rect 20028 -755 20068 -715
rect 17801 -1291 17851 -1241
rect 20536 -2585 20576 -2545
rect 17895 -3117 17945 -3067
rect 21036 -4399 21076 -4359
rect 17757 -4935 17807 -4885
<< metal1 >>
rect 5453 16323 10179 16433
rect 10289 16323 10295 16433
rect 5338 16079 9680 16191
rect 9792 16079 9798 16191
rect 5322 15835 6214 15947
rect 6326 15835 6332 15947
rect 5432 15585 6660 15697
rect 6772 15585 6778 15697
rect 5489 15335 7093 15445
rect 7203 15335 7209 15445
rect -3293 14894 -3287 15136
rect -3045 15015 806 15136
rect -3045 14981 839 15015
rect -3045 14894 806 14981
rect 5471 14701 10787 14787
rect 10873 14701 10879 14787
rect 5362 13382 11195 13447
rect 11260 13382 11266 13447
rect -2363 12404 -2357 12646
rect -2115 12404 1002 12646
rect 5453 12119 7531 12229
rect 7641 12119 7647 12229
rect 5496 11891 7940 12003
rect 8052 11891 8058 12003
rect 5464 11629 8356 11741
rect 8468 11629 8474 11741
rect 5429 10502 12867 10612
rect 12977 10502 12983 10612
rect 5166 10258 11762 10370
rect 11874 10258 11880 10370
rect 5326 10013 6214 10125
rect 6326 10013 6332 10125
rect 5456 9763 6660 9875
rect 6772 9763 6778 9875
rect 5469 9513 7083 9623
rect 7193 9513 7199 9623
rect -3277 9074 -3271 9316
rect -3029 9074 930 9316
rect -1140 8052 -1011 9074
rect 5419 8880 14129 8966
rect 14215 8880 14221 8966
rect -1968 7836 -1840 7848
rect -4208 7720 -4202 7836
rect -4086 7720 -1962 7836
rect -1846 7720 -1840 7836
rect -1968 7708 -1840 7720
rect 5324 7561 15163 7626
rect 15228 7561 15234 7626
rect -1112 6826 -983 7553
rect -2363 6584 -2357 6826
rect -2115 6584 968 6826
rect 5371 6297 7531 6407
rect 7641 6297 7647 6407
rect 5492 6069 7934 6181
rect 8046 6069 8052 6181
rect 5474 5807 8356 5919
rect 8468 5807 8474 5919
rect 5375 4679 13215 4789
rect 13325 4679 13331 4789
rect 5396 4435 12130 4547
rect 12242 4435 12248 4547
rect 5250 4191 6218 4303
rect 6330 4191 6336 4303
rect 5446 3941 6664 4053
rect 6776 3941 6782 4053
rect 5483 3691 7083 3801
rect 7193 3691 7199 3801
rect -3277 3250 -3271 3492
rect -3029 3375 840 3492
rect -3029 3341 895 3375
rect -3029 3250 840 3341
rect -1131 2357 -1001 3250
rect 5319 3057 14415 3143
rect 14501 3057 14507 3143
rect -1950 2134 -1822 2146
rect -4666 2018 -4660 2134
rect -4544 2018 -1944 2134
rect -1828 2018 -1822 2134
rect -1950 2006 -1822 2018
rect -1123 1002 -993 1846
rect 5364 1738 15479 1803
rect 15544 1738 15550 1803
rect 11787 1228 11793 1282
rect 11847 1228 18071 1282
rect 19730 1051 19782 1063
rect 19922 1051 19928 1057
rect 19730 1011 19736 1051
rect 19776 1011 19928 1051
rect -2379 760 -2373 1002
rect -2131 760 842 1002
rect 19730 999 19782 1011
rect 19922 1005 19928 1011
rect 19980 1005 19986 1057
rect 5411 475 7531 585
rect 7641 475 7647 585
rect 17538 446 17544 498
rect 17596 497 17602 498
rect 17829 497 17891 509
rect 17596 447 17835 497
rect 17885 447 17891 497
rect 17596 446 17602 447
rect 17829 435 17891 447
rect 5470 247 7940 359
rect 8052 247 8058 359
rect 12155 168 12161 222
rect 12215 168 18033 222
rect 5470 -15 8360 97
rect 8472 -15 8478 97
rect 12891 -538 12897 -484
rect 12951 -538 18093 -484
rect 20022 -715 20074 -703
rect 20386 -715 20392 -709
rect 20022 -755 20028 -715
rect 20068 -755 20392 -715
rect 20022 -767 20074 -755
rect 20386 -761 20392 -755
rect 20444 -761 20450 -709
rect 17542 -1292 17548 -1240
rect 17600 -1241 17606 -1240
rect 17795 -1241 17857 -1229
rect 17600 -1291 17801 -1241
rect 17851 -1291 17857 -1241
rect 17600 -1292 17606 -1291
rect 17795 -1303 17857 -1291
rect 13243 -1598 13249 -1544
rect 13303 -1598 18075 -1544
rect 14131 -2368 14137 -2314
rect 14191 -2368 18151 -2314
rect 20530 -2545 20582 -2533
rect 20812 -2545 20818 -2539
rect 20530 -2585 20536 -2545
rect 20576 -2585 20818 -2545
rect 20530 -2597 20582 -2585
rect 20812 -2591 20818 -2585
rect 20870 -2591 20876 -2539
rect 17540 -3118 17546 -3066
rect 17598 -3067 17604 -3066
rect 17889 -3067 17951 -3055
rect 17598 -3117 17895 -3067
rect 17945 -3117 17951 -3067
rect 17598 -3118 17604 -3117
rect 17889 -3129 17951 -3117
rect 14433 -3428 14439 -3374
rect 14493 -3428 18071 -3374
rect 15163 -4182 15169 -4128
rect 15223 -4182 18171 -4128
rect 21030 -4359 21082 -4347
rect 21278 -4359 21284 -4353
rect 21030 -4399 21036 -4359
rect 21076 -4399 21284 -4359
rect 21030 -4411 21082 -4399
rect 21278 -4405 21284 -4399
rect 21336 -4405 21342 -4353
rect 17538 -4936 17544 -4884
rect 17596 -4885 17602 -4884
rect 17751 -4885 17813 -4873
rect 17596 -4935 17757 -4885
rect 17807 -4935 17813 -4885
rect 17596 -4936 17602 -4935
rect 17751 -4947 17813 -4935
rect 15483 -5242 15489 -5188
rect 15543 -5242 18073 -5188
rect -3278 -5576 -2912 -5564
rect -3278 -5746 -3228 -5576
rect -3078 -5595 -2912 -5576
rect -3078 -5746 17951 -5595
rect -3278 -5761 17951 -5746
rect -3278 -5780 -2912 -5761
rect 17785 -5955 17951 -5761
rect 17779 -6121 17785 -5955
rect 17951 -6121 17957 -5955
rect -2362 -6264 -2050 -6258
rect -2362 -6430 -2312 -6264
rect -2146 -6267 -2050 -6264
rect -2146 -6430 18595 -6267
rect -2362 -6432 18595 -6430
rect 18760 -6432 18766 -6267
rect -2362 -6450 -2050 -6432
<< via1 >>
rect 10179 16323 10289 16433
rect 9680 16079 9792 16191
rect 6214 15835 6326 15947
rect 6660 15585 6772 15697
rect 7093 15335 7203 15445
rect -3287 14894 -3045 15136
rect 10787 14701 10873 14787
rect 11195 13382 11260 13447
rect -2357 12404 -2115 12646
rect 7531 12119 7641 12229
rect 7940 11891 8052 12003
rect 8356 11629 8468 11741
rect 12867 10502 12977 10612
rect 11762 10258 11874 10370
rect 6214 10013 6326 10125
rect 6660 9763 6772 9875
rect 7083 9513 7193 9623
rect -3271 9074 -3029 9316
rect 14129 8880 14215 8966
rect -4202 7720 -4086 7836
rect 15163 7561 15228 7626
rect -2357 6584 -2115 6826
rect 7531 6297 7641 6407
rect 7934 6069 8046 6181
rect 8356 5807 8468 5919
rect 13215 4679 13325 4789
rect 12130 4435 12242 4547
rect 6218 4191 6330 4303
rect 6664 3941 6776 4053
rect 7083 3691 7193 3801
rect -3271 3250 -3029 3492
rect 14415 3057 14501 3143
rect -4660 2018 -4544 2134
rect 15479 1738 15544 1803
rect 11793 1228 11847 1282
rect -2373 760 -2131 1002
rect 19928 1005 19980 1057
rect 7531 475 7641 585
rect 17544 446 17596 498
rect 7940 247 8052 359
rect 12161 168 12215 222
rect 8360 -15 8472 97
rect 12897 -538 12951 -484
rect 20392 -761 20444 -709
rect 17548 -1292 17600 -1240
rect 13249 -1598 13303 -1544
rect 14137 -2368 14191 -2314
rect 20818 -2591 20870 -2539
rect 17546 -3118 17598 -3066
rect 14439 -3428 14493 -3374
rect 15169 -4182 15223 -4128
rect 21284 -4405 21336 -4353
rect 17544 -4936 17596 -4884
rect 15489 -5242 15543 -5188
rect -3228 -5746 -3078 -5576
rect 17785 -6121 17951 -5955
rect -2312 -6430 -2146 -6264
rect 18595 -6432 18760 -6267
<< metal2 >>
rect -4660 2134 -4544 17848
rect -4660 -6690 -4544 2018
rect -4202 7836 -4086 17380
rect -3271 15142 -3029 17340
rect -3287 15136 -3029 15142
rect -3045 14894 -3029 15136
rect -3287 14888 -3029 14894
rect -4202 -6690 -4086 7720
rect -3271 9316 -3029 14888
rect -3271 3492 -3029 9074
rect -3271 -5576 -3029 3250
rect -2357 12646 -2115 17340
rect -2357 6826 -2115 12404
rect -2357 1008 -2115 6584
rect -2373 1002 -2115 1008
rect -2131 760 -2115 1002
rect -2373 754 -2115 760
rect -3271 -5746 -3228 -5576
rect -3078 -5746 -3029 -5576
rect -3271 -6690 -3029 -5746
rect -2357 -6264 -2115 754
rect -2357 -6430 -2312 -6264
rect -2146 -6430 -2115 -6264
rect -2357 -6690 -2115 -6430
rect 6214 15947 6326 17374
rect 6214 10125 6326 15835
rect 6214 4309 6326 10013
rect 6660 15697 6772 17340
rect 6660 9875 6772 15585
rect 6214 4303 6330 4309
rect 6214 4191 6218 4303
rect 6214 4185 6330 4191
rect 6214 -6690 6326 4185
rect 6660 4059 6772 9763
rect 7083 15451 7193 17340
rect 7083 15445 7203 15451
rect 7083 15335 7093 15445
rect 7083 15329 7203 15335
rect 7083 9623 7193 15329
rect 6660 4053 6776 4059
rect 6660 3941 6664 4053
rect 6660 3935 6776 3941
rect 6660 -6690 6772 3935
rect 7083 3801 7193 9513
rect 7083 -6690 7193 3691
rect 7527 12235 7637 17340
rect 7527 12229 7641 12235
rect 7527 12119 7531 12229
rect 7527 12113 7641 12119
rect 7527 6413 7637 12113
rect 7934 12009 8046 17340
rect 7934 12003 8052 12009
rect 7934 11891 7940 12003
rect 7934 11885 8052 11891
rect 7527 6407 7641 6413
rect 7527 6297 7531 6407
rect 7527 6291 7641 6297
rect 7527 591 7637 6291
rect 7934 6181 8046 11885
rect 7527 585 7641 591
rect 7527 475 7531 585
rect 7527 469 7641 475
rect 7527 -6690 7637 469
rect 7934 365 8046 6069
rect 8356 11741 8468 17340
rect 9680 16191 9792 17372
rect 10179 16433 10289 17339
rect 10179 16317 10289 16323
rect 9680 16073 9792 16079
rect 10787 14787 10873 17327
rect 10787 14695 10873 14701
rect 11195 13447 11260 17364
rect 11195 13376 11260 13382
rect 8356 5919 8468 11629
rect 12867 10612 12977 10618
rect 7934 359 8052 365
rect 7934 247 7940 359
rect 7934 241 8052 247
rect 7934 -6690 8046 241
rect 8356 103 8468 5807
rect 11762 10370 11874 10376
rect 11762 1282 11874 10258
rect 11762 1228 11793 1282
rect 11847 1228 11874 1282
rect 8356 97 8472 103
rect 8356 -15 8360 97
rect 8356 -21 8472 -15
rect 8356 -6690 8468 -21
rect 11762 -6182 11874 1228
rect 12130 4547 12242 4553
rect 12130 222 12242 4435
rect 12130 168 12161 222
rect 12215 168 12242 222
rect 12130 -6270 12242 168
rect 12867 -484 12977 10502
rect 14129 8966 14215 8972
rect 12867 -538 12897 -484
rect 12951 -538 12977 -484
rect 12867 -6287 12977 -538
rect 13215 4789 13325 4795
rect 13215 -1544 13325 4679
rect 13215 -1598 13249 -1544
rect 13303 -1598 13325 -1544
rect 13215 -6235 13325 -1598
rect 14129 -2314 14215 8880
rect 15163 7626 15228 7632
rect 14129 -2368 14137 -2314
rect 14191 -2368 14215 -2314
rect 14129 -6293 14215 -2368
rect 14415 3143 14501 3149
rect 14415 -3374 14501 3057
rect 14415 -3428 14439 -3374
rect 14493 -3428 14501 -3374
rect 14415 -6293 14501 -3428
rect 15163 -4128 15228 7561
rect 15163 -4182 15169 -4128
rect 15223 -4182 15228 -4128
rect 15163 -6282 15228 -4182
rect 15479 1803 15544 1809
rect 15479 -5188 15544 1738
rect 17545 504 17595 18217
rect 19934 1063 19974 18064
rect 19928 1057 19980 1063
rect 19928 999 19980 1005
rect 17544 498 17596 504
rect 17544 440 17596 446
rect 17545 -1234 17595 440
rect 17545 -1240 17600 -1234
rect 17545 -1292 17548 -1240
rect 17545 -1298 17600 -1292
rect 17545 -3060 17595 -1298
rect 17545 -3066 17598 -3060
rect 17545 -3118 17546 -3066
rect 17545 -3124 17598 -3118
rect 17545 -4878 17595 -3124
rect 17544 -4884 17596 -4878
rect 17544 -4942 17596 -4936
rect 15479 -5242 15489 -5188
rect 15543 -5242 15544 -5188
rect 15479 -6246 15544 -5242
rect 17545 -6515 17595 -4942
rect 17785 -5955 17951 -5949
rect 17951 -6121 18325 -5955
rect 18491 -6121 18500 -5955
rect 17785 -6127 17951 -6121
rect 18595 -6267 18760 -6261
rect 19429 -6267 19479 -5573
rect 18760 -6432 19479 -6267
rect 18595 -6438 18760 -6432
rect 19429 -7503 19479 -6432
rect 19934 -7622 19974 999
rect 20398 -703 20438 18006
rect 20392 -709 20444 -703
rect 20392 -767 20444 -761
rect 20398 -7908 20438 -767
rect 20824 -2533 20864 18234
rect 20818 -2539 20870 -2533
rect 20818 -2597 20870 -2591
rect 20824 -7892 20864 -2597
rect 21290 -4347 21330 18110
rect 21284 -4353 21336 -4347
rect 21284 -4411 21336 -4405
rect 21290 -8046 21330 -4411
<< via2 >>
rect 18325 -6121 18491 -5955
<< metal3 >>
rect 18320 -5955 18496 -5950
rect 19286 -5955 19358 -5650
rect 18320 -6121 18325 -5955
rect 18491 -6121 19358 -5955
rect 18320 -6126 18496 -6121
rect 19286 -7514 19358 -6121
use neuron-labeled-extended  neuron-labeled-extended_0
timestamp 1606259729
transform 1 0 630 0 1 623
box -683 -638 4978 4166
use inverter  inverter_0
timestamp 1604367083
transform 1 0 -1166 0 1 2098
box -126 -478 242 448
use one-way  one-way_0
timestamp 1606105257
transform 1 0 -618 0 1 1859
box -37 0 183 688
use neuron-labeled-extended  neuron-labeled-extended_1
timestamp 1606259729
transform 1 0 631 0 1 6446
box -683 -638 4978 4166
use inverter  inverter_1
timestamp 1604367083
transform 1 0 -1150 0 1 7804
box -126 -478 242 448
use one-way  one-way_1
timestamp 1606105257
transform 1 0 -543 0 1 7572
box -37 0 183 688
use neuron-labeled-extended  neuron-labeled-extended_2
timestamp 1606259729
transform 1 0 630 0 1 12267
box -683 -638 4978 4166
use pass-gate-inv-2  pass-gate-inv-2_2
timestamp 1605933175
transform 1 0 18580 0 1 -3752
box -610 -156 899 1683
use pass-gate-inv-2  pass-gate-inv-2_3
timestamp 1605933175
transform 1 0 18580 0 1 -5566
box -610 -156 899 1683
use pass-gate-inv-2  pass-gate-inv-2_1
timestamp 1605933175
transform 1 0 18582 0 1 -1922
box -610 -156 899 1683
use pass-gate-inv-2  pass-gate-inv-2_0
timestamp 1605933175
transform 1 0 18582 0 1 -156
box -610 -156 899 1683
<< labels >>
flabel metal2 6688 17108 6750 17190 0 FreeSans 800 0 0 0 vw
port 1 nsew
flabel metal2 7106 17118 7168 17200 0 FreeSans 800 0 0 0 vth
port 2 nsew
flabel metal2 7536 17148 7598 17230 0 FreeSans 800 0 0 0 vk
port 3 nsew
flabel metal2 7956 17138 8018 17220 0 FreeSans 800 0 0 0 vr
port 4 nsew
flabel metal2 8374 17148 8436 17230 0 FreeSans 800 0 0 0 vad
port 5 nsew
flabel metal2 9694 17180 9756 17262 0 FreeSans 800 0 0 0 v
port 6 nsew
flabel metal2 10196 17180 10258 17262 0 FreeSans 800 0 0 0 u
port 7 nsew
flabel metal2 10810 17158 10872 17240 0 FreeSans 800 0 0 0 a
port 8 nsew
flabel metal2 11212 17160 11234 17202 0 FreeSans 800 0 0 0 axon
port 9 nsew
flabel metal2 -4166 17140 -4144 17182 0 FreeSans 800 0 0 0 syn0
port 15 nsew
flabel metal2 -4618 17220 -4596 17262 0 FreeSans 800 0 0 0 syn1
port 16 nsew
flabel metal2 -3176 17008 -3154 17050 0 FreeSans 800 0 0 0 vdd
port 17 nsew
flabel metal2 -2270 16950 -2248 16992 0 FreeSans 800 0 0 0 vss
port 19 nsew
flabel metal2 6252 17166 6290 17216 0 FreeSans 800 0 0 0 vau
port 20 nsew
flabel metal2 17558 17744 17580 17786 0 FreeSans 800 0 0 0 sel
port 10 nsew
flabel metal2 19944 17708 19966 17750 0 FreeSans 800 0 0 0 v#
port 11 nsew
flabel metal2 20408 17732 20430 17774 0 FreeSans 800 0 0 0 u#
port 12 nsew
flabel metal2 20830 17764 20852 17806 0 FreeSans 800 0 0 0 a#
port 13 nsew
flabel metal2 21302 17782 21324 17824 0 FreeSans 800 0 0 0 axon#
port 14 nsew
<< end >>
