magic
tech sky130A
magscale 1 2
timestamp 1606535953
<< poly >>
rect 2418 4134 2490 4150
rect 2418 4082 2428 4134
rect 2480 4082 2490 4134
rect -209 3901 -119 3917
rect -209 3831 -199 3901
rect -129 3831 -119 3901
rect -209 1998 -119 3831
rect 2187 3652 2267 3668
rect 2187 3592 2197 3652
rect 2257 3592 2267 3652
rect 1778 3401 1858 3417
rect 1778 3341 1788 3401
rect 1848 3341 1858 3401
rect 1778 2913 1858 3341
rect 2187 2908 2267 3592
rect -209 1908 426 1998
rect 2418 1878 2490 4082
rect 2266 1806 2490 1878
rect -251 490 38 570
rect -251 -60 -171 490
rect -251 -120 -241 -60
rect -181 -120 -171 -60
rect -251 -136 -171 -120
rect 1936 -288 2016 52
rect 1936 -348 1946 -288
rect 2006 -348 2016 -288
rect 1936 -364 2016 -348
rect 2909 -547 2989 58
rect 2909 -607 2919 -547
rect 2979 -607 2989 -547
rect 2909 -623 2989 -607
<< polycont >>
rect 2428 4082 2480 4134
rect -199 3831 -129 3901
rect 2197 3592 2257 3652
rect 1788 3341 1848 3401
rect -241 -120 -181 -60
rect 1946 -348 2006 -288
rect 2919 -607 2979 -547
<< locali >>
rect 2414 4144 2494 4150
rect 2414 4074 2420 4144
rect 2490 4074 2494 4144
rect 2414 4066 2494 4074
rect -220 3902 -110 3918
rect -220 3832 -200 3902
rect -130 3901 -110 3902
rect -220 3831 -199 3832
rect -129 3831 -110 3901
rect -220 3816 -110 3831
rect 2178 3658 2276 3670
rect 2178 3588 2192 3658
rect 2262 3588 2276 3658
rect 2178 3576 2276 3588
rect 1766 3406 1864 3420
rect 1766 3336 1782 3406
rect 1852 3336 1864 3406
rect 1766 3326 1864 3336
rect -90 3150 -25 3178
rect -90 2294 -25 3088
rect 3628 2434 4171 2520
rect 4257 2434 4262 2520
rect -28 2277 -25 2294
rect 4284 1116 4294 1180
rect 4284 1115 4358 1116
rect -258 -56 -164 -48
rect -258 -126 -246 -56
rect -176 -126 -164 -56
rect -258 -138 -164 -126
rect 1924 -284 2024 -272
rect 1924 -354 1940 -284
rect 2010 -354 2024 -284
rect 1924 -370 2024 -354
rect 2898 -544 2998 -536
rect 2898 -614 2914 -544
rect 2984 -614 2998 -544
rect 2898 -626 2998 -614
<< viali >>
rect 2420 4134 2490 4144
rect 2420 4082 2428 4134
rect 2428 4082 2480 4134
rect 2480 4082 2490 4134
rect 2420 4074 2490 4082
rect -200 3901 -130 3902
rect -200 3832 -199 3901
rect -199 3832 -130 3901
rect 2192 3652 2262 3658
rect 2192 3592 2197 3652
rect 2197 3592 2257 3652
rect 2257 3592 2262 3652
rect 2192 3588 2262 3592
rect 1782 3401 1852 3406
rect 1782 3341 1788 3401
rect 1788 3341 1848 3401
rect 1848 3341 1852 3401
rect 1782 3336 1852 3341
rect -98 3088 -18 3150
rect 4171 2434 4257 2520
rect -90 2242 -28 2294
rect 4294 1116 4358 1180
rect -246 -60 -176 -56
rect -246 -120 -241 -60
rect -241 -120 -181 -60
rect -181 -120 -176 -60
rect -246 -126 -176 -120
rect 1940 -288 2010 -284
rect 1940 -348 1946 -288
rect 1946 -348 2006 -288
rect 2006 -348 2010 -288
rect 1940 -354 2010 -348
rect 2914 -547 2984 -544
rect 2914 -607 2919 -547
rect 2919 -607 2979 -547
rect 2979 -607 2984 -547
rect 2914 -614 2984 -607
<< metal1 >>
rect -649 4400 10399 4416
rect -649 4326 5626 4400
rect 5724 4398 8112 4400
rect 5724 4326 6882 4398
rect -649 4324 6882 4326
rect 6980 4326 8112 4398
rect 8210 4398 10399 4400
rect 8210 4326 9372 4398
rect 6980 4324 9372 4326
rect 9470 4324 10399 4398
rect -649 4306 10399 4324
rect -643 4152 9443 4166
rect -643 4144 6728 4152
rect -643 4074 2420 4144
rect 2490 4074 6728 4144
rect 6834 4074 9443 4152
rect -643 4056 9443 4074
rect -650 3910 9444 3924
rect -650 3902 5492 3910
rect -650 3832 -200 3902
rect -130 3832 5492 3902
rect -650 3830 5492 3832
rect 5590 3830 9444 3910
rect -650 3812 9444 3830
rect -1100 3658 10416 3680
rect -1100 3588 2192 3658
rect 2262 3588 10416 3658
rect -1100 3568 10416 3588
rect -1114 3406 10426 3430
rect -1114 3336 1782 3406
rect 1852 3336 10426 3406
rect -1114 3318 10426 3336
rect -1113 3150 10425 3178
rect -1113 3088 -98 3150
rect -18 3088 10425 3150
rect -1113 3068 10425 3088
rect 5103 2832 9507 2847
rect 804 2668 814 2818
rect 1120 2668 1130 2818
rect 2638 2670 2648 2820
rect 2954 2670 2964 2820
rect 3358 2670 3368 2820
rect 3674 2670 3684 2820
rect 5103 2772 7966 2832
rect 8054 2772 9507 2832
rect 5103 2761 9507 2772
rect 4165 2520 4263 2532
rect 5103 2520 5189 2761
rect 4165 2434 4171 2520
rect 4257 2434 5189 2520
rect 5355 2526 9226 2582
rect 9294 2526 9411 2582
rect 5355 2524 9411 2526
rect 4165 2422 4263 2434
rect -102 2294 -16 2300
rect -102 2242 -90 2294
rect -28 2242 -16 2294
rect -102 2236 -16 2242
rect -87 2086 -29 2236
rect -87 2028 92 2086
rect 5355 1895 5413 2524
rect 6546 2206 10595 2348
rect 5640 1946 5646 1998
rect 5698 1993 5704 1998
rect 5698 1951 5831 1993
rect 5698 1946 5704 1951
rect 6898 1946 6904 1998
rect 6956 1993 6962 1998
rect 6956 1951 7093 1993
rect 6956 1946 6962 1951
rect 8128 1946 8134 1998
rect 8186 1993 8192 1998
rect 8186 1951 8337 1993
rect 8186 1946 8192 1951
rect 9384 1946 9390 1998
rect 9442 1993 9448 1998
rect 9442 1951 9603 1993
rect 9442 1946 9448 1951
rect 4747 1837 5413 1895
rect 4282 1180 4372 1194
rect 4747 1180 4805 1837
rect 5508 1766 5514 1818
rect 5566 1813 5572 1818
rect 5566 1771 5833 1813
rect 5566 1766 5572 1771
rect 6746 1766 6752 1818
rect 6804 1813 6810 1818
rect 6804 1771 7089 1813
rect 6804 1766 6810 1771
rect 7978 1766 7984 1818
rect 8036 1813 8042 1818
rect 8036 1771 8341 1813
rect 8036 1766 8042 1771
rect 9228 1766 9234 1818
rect 9286 1813 9292 1818
rect 9286 1771 9595 1813
rect 9286 1766 9292 1771
rect 6473 1497 6515 1641
rect 6670 1539 6676 1544
rect 6522 1497 6676 1539
rect 6670 1492 6676 1497
rect 6728 1492 6734 1544
rect 7717 1497 7759 1655
rect 7946 1539 7952 1544
rect 7772 1497 7952 1539
rect 7946 1492 7952 1497
rect 8004 1492 8010 1544
rect 8939 1497 8981 1651
rect 9142 1539 9148 1544
rect 8995 1497 9148 1539
rect 9142 1492 9148 1497
rect 9200 1492 9206 1544
rect 10211 1497 10253 1647
rect 10318 1539 10324 1544
rect 10259 1497 10324 1539
rect 10318 1492 10324 1497
rect 10376 1492 10382 1544
rect 5147 1180 10633 1322
rect 4282 1116 4294 1180
rect 4358 1116 4830 1180
rect 4282 1115 4830 1116
rect 4282 1103 4372 1115
rect 5147 351 5289 1180
rect 6284 1030 10468 1042
rect 6284 942 6652 1030
rect 6754 942 10468 1030
rect 6284 930 10468 942
rect 7092 820 10462 830
rect 7092 732 7932 820
rect 8034 732 10462 820
rect 7092 718 10462 732
rect 8524 608 10468 617
rect 8524 520 9126 608
rect 9228 520 10468 608
rect 8524 505 10468 520
rect 3573 328 5289 351
rect 3573 209 3620 328
rect 3610 178 3620 209
rect 3926 209 5289 328
rect 10062 394 10476 405
rect 10062 306 10294 394
rect 10396 306 10476 394
rect 10062 293 10476 306
rect 3926 178 3936 209
rect -1011 -56 10491 -38
rect -1011 -126 -246 -56
rect -176 -126 10491 -56
rect -1011 -148 10491 -126
rect -998 -284 10504 -264
rect -998 -354 1940 -284
rect 2010 -354 10504 -284
rect -998 -376 10504 -354
rect -1012 -544 10492 -526
rect -1012 -614 2914 -544
rect 2984 -614 10492 -544
rect -1012 -638 10492 -614
<< via1 >>
rect 5626 4326 5724 4400
rect 6882 4324 6980 4398
rect 8112 4326 8210 4400
rect 9372 4324 9470 4398
rect 6728 4074 6834 4152
rect 5492 3830 5590 3910
rect 814 2668 1120 2818
rect 2648 2670 2954 2820
rect 3368 2670 3674 2820
rect 7966 2772 8054 2832
rect 9226 2526 9294 2582
rect 5646 1946 5698 1998
rect 6904 1946 6956 1998
rect 8134 1946 8186 1998
rect 9390 1946 9442 1998
rect 5514 1766 5566 1818
rect 6752 1766 6804 1818
rect 7984 1766 8036 1818
rect 9234 1766 9286 1818
rect 6676 1492 6728 1544
rect 7952 1492 8004 1544
rect 9148 1492 9200 1544
rect 10324 1492 10376 1544
rect 4294 1116 4358 1180
rect 6652 942 6754 1030
rect 7932 732 8034 820
rect 9126 520 9228 608
rect 3620 178 3926 328
rect 10294 306 10396 394
<< metal2 >>
rect 5626 4400 5724 4410
rect 5626 4316 5724 4326
rect 6882 4398 6980 4408
rect 5492 3910 5590 3920
rect 5492 3820 5590 3830
rect 814 2818 1120 2828
rect 814 2658 1120 2668
rect 2648 2820 2954 2830
rect 2648 2660 2954 2670
rect 3368 2820 3674 2830
rect 3368 2660 3674 2670
rect 5519 1824 5561 3820
rect 5651 2004 5693 4316
rect 6882 4314 6980 4324
rect 8112 4400 8210 4410
rect 8112 4316 8210 4326
rect 9372 4398 9470 4408
rect 6728 4152 6834 4162
rect 6728 4064 6834 4074
rect 5646 1998 5698 2004
rect 5646 1940 5698 1946
rect 6757 1824 6799 4064
rect 6909 2004 6951 4314
rect 7966 2832 8054 2842
rect 7966 2762 8054 2772
rect 6904 1998 6956 2004
rect 6904 1940 6956 1946
rect 7989 1824 8031 2762
rect 8139 2004 8181 4316
rect 9372 4314 9470 4324
rect 9226 2582 9294 2592
rect 9226 2516 9294 2526
rect 8134 1998 8186 2004
rect 8134 1940 8186 1946
rect 9239 1824 9281 2516
rect 9395 2004 9437 4314
rect 9390 1998 9442 2004
rect 9390 1940 9442 1946
rect 5514 1818 5566 1824
rect 5514 1760 5566 1766
rect 6752 1818 6804 1824
rect 6752 1760 6804 1766
rect 7984 1818 8036 1824
rect 7984 1760 8036 1766
rect 9234 1818 9286 1824
rect 9234 1760 9286 1766
rect 6676 1544 6728 1550
rect 6676 1486 6728 1492
rect 7952 1544 8004 1550
rect 7952 1486 8004 1492
rect 9148 1544 9200 1550
rect 9148 1486 9200 1492
rect 10324 1544 10376 1550
rect 10324 1486 10376 1492
rect 4294 1180 4358 1190
rect 1521 1116 4294 1180
rect 4294 1106 4358 1116
rect 6681 1040 6723 1486
rect 6652 1030 6754 1040
rect 6652 932 6754 942
rect 7957 830 7999 1486
rect 7932 820 8034 830
rect 7932 722 8034 732
rect 9153 618 9195 1486
rect 9126 608 9228 618
rect 9126 510 9228 520
rect 10329 404 10371 1486
rect 10294 394 10396 404
rect 3620 328 3926 338
rect 10294 296 10396 306
rect 3620 168 3926 178
<< via2 >>
rect 814 2668 1120 2818
rect 2648 2670 2954 2820
rect 3368 2670 3674 2820
rect 3620 178 3926 328
<< metal3 >>
rect -1107 2820 4928 2866
rect -1107 2818 2648 2820
rect -1107 2668 814 2818
rect 1120 2670 2648 2818
rect 2954 2670 3368 2820
rect 3674 2670 4928 2820
rect 1120 2668 4928 2670
rect -1107 2624 4928 2668
rect 3878 379 4120 380
rect -1011 328 4928 379
rect -1011 178 3620 328
rect 3926 178 4928 328
rect -1011 141 4928 178
rect 3878 138 4120 141
use neuron-labeled  neuron-labeled_0
timestamp 1604452313
transform 1 0 364 0 1 678
box -364 -678 3630 2294
use pmos-diff-amp  pmos-diff-amp_0
timestamp 1606516043
transform 1 0 6001 0 1 1657
box -231 -477 703 691
use pmos-diff-amp  pmos-diff-amp_1
timestamp 1606516043
transform 1 0 7251 0 1 1657
box -231 -477 703 691
use pmos-diff-amp  pmos-diff-amp_2
timestamp 1606516043
transform 1 0 8477 0 1 1657
box -231 -477 703 691
use pmos-diff-amp  pmos-diff-amp_3
timestamp 1606516043
transform 1 0 9749 0 1 1657
box -231 -477 703 691
<< labels >>
flabel metal1 -598 3840 -548 3886 0 FreeSans 800 0 0 0 v
port 0 nsew
flabel metal1 -596 4090 -546 4120 0 FreeSans 800 0 0 0 u
port 1 nsew
flabel metal1 -1064 3586 -1014 3630 0 FreeSans 800 0 0 0 vau
port 3 nsew
flabel metal1 -1064 3350 -1014 3380 0 FreeSans 800 0 0 0 vw
port 4 nsew
flabel metal1 -1070 3094 -1020 3124 0 FreeSans 800 0 0 0 vth
port 6 nsew
flabel metal1 -986 -122 -928 -80 0 FreeSans 800 0 0 0 vk
port 7 nsew
flabel metal1 -956 -350 -898 -308 0 FreeSans 800 0 0 0 vr
port 8 nsew
flabel metal1 -970 -600 -912 -558 0 FreeSans 800 0 0 0 vad
port 9 nsew
flabel metal3 -1042 2680 -936 2786 0 FreeSans 800 0 0 0 vdd
port 10 nsew
flabel metal1 8526 2774 8584 2824 0 FreeSans 800 0 0 0 a
port 2 nsew
flabel metal1 8422 2530 8472 2560 0 FreeSans 800 0 0 0 axon
port 12 nsew
flabel metal1 10218 4328 10298 4370 0 FreeSans 800 0 0 0 i_bias
port 13 nsew
flabel metal1 10004 970 10084 1012 0 FreeSans 800 0 0 0 v_buff
port 14 nsew
flabel metal1 10040 734 10120 776 0 FreeSans 800 0 0 0 u_buff
port 15 nsew
flabel metal1 10068 540 10148 582 0 FreeSans 800 0 0 0 a_buff
port 16 nsew
flabel metal1 10148 330 10228 372 0 FreeSans 800 0 0 0 axon_buff
port 17 nsew
flabel metal1 10464 2230 10534 2300 0 FreeSans 800 0 0 0 vdd_aux
port 18 nsew
flabel metal3 -928 206 -822 312 0 FreeSans 800 0 0 0 vss
port 11 nsew
<< end >>
