magic
tech sky130A
timestamp 1608000372
<< metal1 >>
rect 2051 2833 2083 3926
rect 1750 2814 2083 2833
rect 1750 2805 2070 2814
rect 1755 2747 1785 2805
rect 1843 2248 1877 2307
rect 2078 2248 2115 2250
rect 1843 2221 2115 2248
rect 1847 2210 2115 2221
rect 2078 1411 2115 2210
rect 2058 1374 2115 1411
<< metal2 >>
rect 222 2415 245 3013
<< metal3 >>
rect 1554 4059 1591 4677
rect 1554 4045 1603 4059
rect 1405 3997 1603 4045
rect 88 2411 121 2875
rect 888 2398 932 3671
rect 1005 2814 1043 2828
rect 1076 2823 1476 2825
rect 1561 2823 1603 3997
rect 1076 2814 1603 2823
rect 1005 2790 1603 2814
rect 1005 2781 1596 2790
rect 1005 2614 1043 2781
rect 1076 2778 1476 2781
rect 1003 2503 1043 2614
rect 1003 2279 1041 2503
rect 1003 2277 1132 2279
rect 1457 2277 1593 2279
rect 1003 2246 1593 2277
rect 1029 2242 1593 2246
rect 1059 2239 1593 2242
rect 1457 2237 1593 2239
rect 1544 1536 1587 2237
rect 1403 1522 1587 1536
rect 1403 1503 1582 1522
<< metal4 >>
rect 435 2401 473 2578
use Sw-1  Sw-1_0
timestamp 1608000372
transform 1 0 1173 0 1 2246
box -70 45 891 509
use 3good  3good_0
timestamp 1608000372
transform 1 0 -2 0 1 -1
box 1 3 2076 2588
use 3good  3good_1
timestamp 1608000372
transform 1 0 4 0 1 2517
box 1 3 2076 2588
<< end >>
