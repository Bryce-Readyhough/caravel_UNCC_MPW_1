magic
tech sky130A
magscale 1 2
timestamp 1606259729
<< poly >>
rect 2418 4134 2490 4150
rect 2418 4082 2428 4134
rect 2480 4082 2490 4134
rect -209 3901 -119 3917
rect -209 3831 -199 3901
rect -129 3831 -119 3901
rect -209 1998 -119 3831
rect 2187 3652 2267 3668
rect 2187 3592 2197 3652
rect 2257 3592 2267 3652
rect 1778 3401 1858 3417
rect 1778 3341 1788 3401
rect 1848 3341 1858 3401
rect 1778 2913 1858 3341
rect 2187 2908 2267 3592
rect -209 1908 426 1998
rect 2418 1878 2490 4082
rect 2266 1806 2490 1878
rect -251 490 38 570
rect -251 -60 -171 490
rect -251 -120 -241 -60
rect -181 -120 -171 -60
rect -251 -136 -171 -120
rect 1936 -288 2016 52
rect 1936 -348 1946 -288
rect 2006 -348 2016 -288
rect 1936 -364 2016 -348
rect 2909 -547 2989 58
rect 2909 -607 2919 -547
rect 2979 -607 2989 -547
rect 2909 -623 2989 -607
<< polycont >>
rect 2428 4082 2480 4134
rect -199 3831 -129 3901
rect 2197 3592 2257 3652
rect 1788 3341 1848 3401
rect -241 -120 -181 -60
rect 1946 -348 2006 -288
rect 2919 -607 2979 -547
<< locali >>
rect 2414 4144 2494 4150
rect 2414 4074 2420 4144
rect 2490 4074 2494 4144
rect 2414 4066 2494 4074
rect -220 3902 -110 3918
rect -220 3832 -200 3902
rect -130 3901 -110 3902
rect -220 3831 -199 3832
rect -129 3831 -110 3901
rect -220 3816 -110 3831
rect 2178 3658 2276 3670
rect 2178 3588 2192 3658
rect 2262 3588 2276 3658
rect 2178 3576 2276 3588
rect 1766 3406 1864 3420
rect 1766 3336 1782 3406
rect 1852 3336 1864 3406
rect 1766 3326 1864 3336
rect -90 3150 -25 3178
rect -90 2294 -25 3088
rect 3628 2434 4171 2520
rect 4257 2434 4262 2520
rect -28 2277 -25 2294
rect 4284 1116 4294 1180
rect 4284 1115 4358 1116
rect -258 -56 -164 -48
rect -258 -126 -246 -56
rect -176 -126 -164 -56
rect -258 -138 -164 -126
rect 1924 -284 2024 -272
rect 1924 -354 1940 -284
rect 2010 -354 2024 -284
rect 1924 -370 2024 -354
rect 2898 -544 2998 -536
rect 2898 -614 2914 -544
rect 2984 -614 2998 -544
rect 2898 -626 2998 -614
<< viali >>
rect 2420 4134 2490 4144
rect 2420 4082 2428 4134
rect 2428 4082 2480 4134
rect 2480 4082 2490 4134
rect 2420 4074 2490 4082
rect -200 3901 -130 3902
rect -200 3832 -199 3901
rect -199 3832 -130 3901
rect 2192 3652 2262 3658
rect 2192 3592 2197 3652
rect 2197 3592 2257 3652
rect 2257 3592 2262 3652
rect 2192 3588 2262 3592
rect 1782 3401 1852 3406
rect 1782 3341 1788 3401
rect 1788 3341 1848 3401
rect 1848 3341 1852 3401
rect 1782 3336 1852 3341
rect -98 3088 -18 3150
rect 4171 2434 4257 2520
rect -90 2242 -28 2294
rect 4294 1116 4358 1180
rect -246 -60 -176 -56
rect -246 -120 -241 -60
rect -241 -120 -181 -60
rect -181 -120 -176 -60
rect -246 -126 -176 -120
rect 1940 -288 2010 -284
rect 1940 -348 1946 -288
rect 1946 -348 2006 -288
rect 2006 -348 2010 -288
rect 1940 -354 2010 -348
rect 2914 -547 2984 -544
rect 2914 -607 2919 -547
rect 2919 -607 2979 -547
rect 2979 -607 2984 -547
rect 2914 -614 2984 -607
<< metal1 >>
rect -641 4144 4933 4166
rect -641 4074 2420 4144
rect 2490 4074 4933 4144
rect -641 4056 4933 4074
rect -646 3902 4936 3924
rect -646 3832 -200 3902
rect -130 3832 4936 3902
rect -646 3812 4936 3832
rect -652 3658 4928 3680
rect -652 3588 2192 3658
rect 2262 3588 4928 3658
rect -652 3568 4928 3588
rect -664 3406 4938 3430
rect -664 3336 1782 3406
rect 1852 3336 4938 3406
rect -664 3318 4938 3336
rect -683 3150 4969 3178
rect -683 3088 -98 3150
rect -18 3088 4969 3150
rect -683 3068 4969 3088
rect 804 2668 814 2818
rect 1120 2668 1130 2818
rect 2638 2670 2648 2820
rect 2954 2670 2964 2820
rect 3358 2670 3368 2820
rect 3674 2670 3684 2820
rect 4165 2520 4263 2532
rect 4165 2434 4171 2520
rect 4257 2434 4927 2520
rect 4165 2422 4263 2434
rect -102 2294 -16 2300
rect -102 2242 -90 2294
rect -28 2242 -16 2294
rect -102 2236 -16 2242
rect -87 2086 -29 2236
rect -87 2028 92 2086
rect 4282 1180 4372 1194
rect 4282 1116 4294 1180
rect 4358 1116 4928 1180
rect 4282 1115 4928 1116
rect 4282 1103 4372 1115
rect 3610 178 3620 328
rect 3926 178 3936 328
rect -629 -56 4953 -38
rect -629 -126 -246 -56
rect -176 -126 4953 -56
rect -629 -148 4953 -126
rect -642 -284 4978 -264
rect -642 -354 1940 -284
rect 2010 -354 4978 -284
rect -642 -376 4978 -354
rect -640 -544 4968 -526
rect -640 -614 2914 -544
rect 2984 -614 4968 -544
rect -640 -638 4968 -614
<< via1 >>
rect 814 2668 1120 2818
rect 2648 2670 2954 2820
rect 3368 2670 3674 2820
rect 4294 1116 4358 1180
rect 3620 178 3926 328
<< metal2 >>
rect 814 2818 1120 2828
rect 814 2658 1120 2668
rect 2648 2820 2954 2830
rect 2648 2660 2954 2670
rect 3368 2820 3674 2830
rect 3368 2660 3674 2670
rect 4294 1180 4358 1190
rect 1521 1116 4294 1180
rect 4294 1106 4358 1116
rect 3620 328 3926 338
rect 3620 168 3926 178
<< via2 >>
rect 814 2668 1120 2818
rect 2648 2670 2954 2820
rect 3368 2670 3674 2820
rect 3620 178 3926 328
<< metal3 >>
rect -630 2820 4928 2866
rect -630 2818 2648 2820
rect -630 2668 814 2818
rect 1120 2670 2648 2818
rect 2954 2670 3368 2820
rect 3674 2670 4928 2820
rect 1120 2668 4928 2670
rect -630 2624 4928 2668
rect 3878 379 4120 380
rect -630 328 4928 379
rect -630 178 3620 328
rect 3926 178 4928 328
rect -630 141 4928 178
rect 3878 138 4120 141
use neuron-labeled  neuron-labeled_0
timestamp 1604452313
transform 1 0 364 0 1 678
box -364 -678 3630 2294
<< labels >>
flabel metal3 -526 2692 -422 2786 0 FreeSans 800 0 0 0 vdd
port 10 nsew
flabel metal3 -546 210 -442 304 0 FreeSans 800 0 0 0 vss
port 12 nsew
flabel metal1 -594 -116 -556 -76 0 FreeSans 800 0 0 0 vk
port 5 nsew
flabel metal1 -614 -348 -568 -306 0 FreeSans 800 0 0 0 vr
port 13 nsew
flabel metal1 -606 -606 -570 -560 0 FreeSans 800 0 0 0 vad
port 14 nsew
flabel metal1 -582 4080 -540 4142 0 FreeSans 800 0 0 0 u
port 15 nsew
flabel metal1 -592 3836 -534 3896 0 FreeSans 800 0 0 0 v
port 16 nsew
flabel locali s -608 3594 -564 3644 0 FreeSans 800 0 0 0 vau
port 17 nsew
flabel locali s -618 3346 -580 3394 0 FreeSans 800 0 0 0 vw
port 18 nsew
flabel locali s -640 3094 -590 3144 0 FreeSans 800 0 0 0 vth
port 19 nsew
flabel locali s 4848 2450 4886 2496 0 FreeSans 800 0 0 0 a
port 20 nsew
flabel locali s 4882 1132 4904 1162 0 FreeSans 800 0 0 0 axon
port 21 nsew
<< end >>
