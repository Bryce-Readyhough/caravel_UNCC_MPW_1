magic
tech sky130A
magscale 1 2
timestamp 1608006408
<< checkpaint >>
rect -1260 -1260 718860 1038860
<< metal1 >>
rect 447760 1005711 447766 1005723
rect 437218 1005683 447766 1005711
rect 437218 1005575 437246 1005683
rect 447760 1005671 447766 1005683
rect 447818 1005671 447824 1005723
rect 469168 1005637 469174 1005649
rect 440482 1005609 469174 1005637
rect 95056 1005523 95062 1005575
rect 95114 1005563 95120 1005575
rect 95114 1005535 108734 1005563
rect 95114 1005523 95120 1005535
rect 108706 1005501 108734 1005535
rect 437200 1005523 437206 1005575
rect 437258 1005523 437264 1005575
rect 93616 1005449 93622 1005501
rect 93674 1005489 93680 1005501
rect 100720 1005489 100726 1005501
rect 93674 1005461 100726 1005489
rect 93674 1005449 93680 1005461
rect 100720 1005449 100726 1005461
rect 100778 1005449 100784 1005501
rect 108688 1005449 108694 1005501
rect 108746 1005449 108752 1005501
rect 433264 1005449 433270 1005501
rect 433322 1005489 433328 1005501
rect 440482 1005489 440510 1005609
rect 469168 1005597 469174 1005609
rect 469226 1005597 469232 1005649
rect 466480 1005563 466486 1005575
rect 441730 1005535 466486 1005563
rect 433322 1005461 440510 1005489
rect 433322 1005449 433328 1005461
rect 440560 1005449 440566 1005501
rect 440618 1005489 440624 1005501
rect 441616 1005489 441622 1005501
rect 440618 1005461 441622 1005489
rect 440618 1005449 440624 1005461
rect 441616 1005449 441622 1005461
rect 441674 1005449 441680 1005501
rect 93712 1005375 93718 1005427
rect 93770 1005415 93776 1005427
rect 115216 1005415 115222 1005427
rect 93770 1005387 115222 1005415
rect 93770 1005375 93776 1005387
rect 115216 1005375 115222 1005387
rect 115274 1005375 115280 1005427
rect 358672 1005375 358678 1005427
rect 358730 1005415 358736 1005427
rect 379120 1005415 379126 1005427
rect 358730 1005387 379126 1005415
rect 358730 1005375 358736 1005387
rect 379120 1005375 379126 1005387
rect 379178 1005375 379184 1005427
rect 431632 1005375 431638 1005427
rect 431690 1005415 431696 1005427
rect 441730 1005415 441758 1005535
rect 466480 1005523 466486 1005535
rect 466538 1005523 466544 1005575
rect 443440 1005449 443446 1005501
rect 443498 1005489 443504 1005501
rect 470992 1005489 470998 1005501
rect 443498 1005461 470998 1005489
rect 443498 1005449 443504 1005461
rect 470992 1005449 470998 1005461
rect 471050 1005449 471056 1005501
rect 504592 1005449 504598 1005501
rect 504650 1005489 504656 1005501
rect 504650 1005461 516926 1005489
rect 504650 1005449 504656 1005461
rect 431690 1005387 441758 1005415
rect 431690 1005375 431696 1005387
rect 441808 1005375 441814 1005427
rect 441866 1005415 441872 1005427
rect 471856 1005415 471862 1005427
rect 441866 1005387 471862 1005415
rect 441866 1005375 441872 1005387
rect 471856 1005375 471862 1005387
rect 471914 1005375 471920 1005427
rect 498736 1005375 498742 1005427
rect 498794 1005415 498800 1005427
rect 512656 1005415 512662 1005427
rect 498794 1005387 512662 1005415
rect 498794 1005375 498800 1005387
rect 512656 1005375 512662 1005387
rect 512714 1005375 512720 1005427
rect 92560 1005301 92566 1005353
rect 92618 1005341 92624 1005353
rect 109456 1005341 109462 1005353
rect 92618 1005313 109462 1005341
rect 92618 1005301 92624 1005313
rect 109456 1005301 109462 1005313
rect 109514 1005301 109520 1005353
rect 298288 1005301 298294 1005353
rect 298346 1005341 298352 1005353
rect 308752 1005341 308758 1005353
rect 298346 1005313 308758 1005341
rect 298346 1005301 298352 1005313
rect 308752 1005301 308758 1005313
rect 308810 1005301 308816 1005353
rect 365008 1005301 365014 1005353
rect 365066 1005341 365072 1005353
rect 383632 1005341 383638 1005353
rect 365066 1005313 383638 1005341
rect 365066 1005301 365072 1005313
rect 383632 1005301 383638 1005313
rect 383690 1005301 383696 1005353
rect 425296 1005301 425302 1005353
rect 425354 1005341 425360 1005353
rect 434704 1005341 434710 1005353
rect 425354 1005313 434710 1005341
rect 425354 1005301 425360 1005313
rect 434704 1005301 434710 1005313
rect 434762 1005301 434768 1005353
rect 434800 1005301 434806 1005353
rect 434858 1005341 434864 1005353
rect 437776 1005341 437782 1005353
rect 434858 1005313 437782 1005341
rect 434858 1005301 434864 1005313
rect 437776 1005301 437782 1005313
rect 437834 1005341 437840 1005353
rect 440560 1005341 440566 1005353
rect 437834 1005313 440566 1005341
rect 437834 1005301 437840 1005313
rect 440560 1005301 440566 1005313
rect 440618 1005301 440624 1005353
rect 452944 1005341 452950 1005353
rect 440962 1005313 452950 1005341
rect 92368 1005227 92374 1005279
rect 92426 1005267 92432 1005279
rect 106576 1005267 106582 1005279
rect 92426 1005239 106582 1005267
rect 92426 1005227 92432 1005239
rect 106576 1005227 106582 1005239
rect 106634 1005227 106640 1005279
rect 217264 1005227 217270 1005279
rect 217322 1005267 217328 1005279
rect 218896 1005267 218902 1005279
rect 217322 1005239 218902 1005267
rect 217322 1005227 217328 1005239
rect 218896 1005227 218902 1005239
rect 218954 1005227 218960 1005279
rect 299536 1005227 299542 1005279
rect 299594 1005267 299600 1005279
rect 309616 1005267 309622 1005279
rect 299594 1005239 309622 1005267
rect 299594 1005227 299600 1005239
rect 309616 1005227 309622 1005239
rect 309674 1005227 309680 1005279
rect 424528 1005227 424534 1005279
rect 424586 1005267 424592 1005279
rect 440848 1005267 440854 1005279
rect 424586 1005239 440854 1005267
rect 424586 1005227 424592 1005239
rect 440848 1005227 440854 1005239
rect 440906 1005227 440912 1005279
rect 198736 1005153 198742 1005205
rect 198794 1005193 198800 1005205
rect 207280 1005193 207286 1005205
rect 198794 1005165 207286 1005193
rect 198794 1005153 198800 1005165
rect 207280 1005153 207286 1005165
rect 207338 1005153 207344 1005205
rect 305296 1005153 305302 1005205
rect 305354 1005193 305360 1005205
rect 314224 1005193 314230 1005205
rect 305354 1005165 314230 1005193
rect 305354 1005153 305360 1005165
rect 314224 1005153 314230 1005165
rect 314282 1005153 314288 1005205
rect 325456 1005153 325462 1005205
rect 325514 1005193 325520 1005205
rect 331216 1005193 331222 1005205
rect 325514 1005165 331222 1005193
rect 325514 1005153 325520 1005165
rect 331216 1005153 331222 1005165
rect 331274 1005153 331280 1005205
rect 358000 1005153 358006 1005205
rect 358058 1005193 358064 1005205
rect 383536 1005193 383542 1005205
rect 358058 1005165 383542 1005193
rect 358058 1005153 358064 1005165
rect 383536 1005153 383542 1005165
rect 383594 1005153 383600 1005205
rect 426064 1005153 426070 1005205
rect 426122 1005193 426128 1005205
rect 440962 1005193 440990 1005313
rect 452944 1005301 452950 1005313
rect 453002 1005301 453008 1005353
rect 441040 1005227 441046 1005279
rect 441098 1005267 441104 1005279
rect 472048 1005267 472054 1005279
rect 441098 1005239 472054 1005267
rect 441098 1005227 441104 1005239
rect 472048 1005227 472054 1005239
rect 472106 1005227 472112 1005279
rect 502288 1005227 502294 1005279
rect 502346 1005267 502352 1005279
rect 516784 1005267 516790 1005279
rect 502346 1005239 516790 1005267
rect 502346 1005227 502352 1005239
rect 516784 1005227 516790 1005239
rect 516842 1005227 516848 1005279
rect 516898 1005267 516926 1005461
rect 572848 1005415 572854 1005427
rect 562306 1005387 572854 1005415
rect 521392 1005267 521398 1005279
rect 516898 1005239 521398 1005267
rect 521392 1005227 521398 1005239
rect 521450 1005227 521456 1005279
rect 554512 1005227 554518 1005279
rect 554570 1005267 554576 1005279
rect 562306 1005267 562334 1005387
rect 572848 1005375 572854 1005387
rect 572906 1005375 572912 1005427
rect 571888 1005267 571894 1005279
rect 554570 1005239 562334 1005267
rect 562402 1005239 571894 1005267
rect 554570 1005227 554576 1005239
rect 443440 1005193 443446 1005205
rect 426122 1005165 440990 1005193
rect 441058 1005165 443446 1005193
rect 426122 1005153 426128 1005165
rect 435568 1005079 435574 1005131
rect 435626 1005119 435632 1005131
rect 440752 1005119 440758 1005131
rect 435626 1005091 440758 1005119
rect 435626 1005079 435632 1005091
rect 440752 1005079 440758 1005091
rect 440810 1005119 440816 1005131
rect 441058 1005119 441086 1005165
rect 443440 1005153 443446 1005165
rect 443498 1005153 443504 1005205
rect 447760 1005153 447766 1005205
rect 447818 1005193 447824 1005205
rect 469360 1005193 469366 1005205
rect 447818 1005165 469366 1005193
rect 447818 1005153 447824 1005165
rect 469360 1005153 469366 1005165
rect 469418 1005153 469424 1005205
rect 508624 1005153 508630 1005205
rect 508682 1005193 508688 1005205
rect 523984 1005193 523990 1005205
rect 508682 1005165 523990 1005193
rect 508682 1005153 508688 1005165
rect 523984 1005153 523990 1005165
rect 524042 1005153 524048 1005205
rect 553744 1005153 553750 1005205
rect 553802 1005193 553808 1005205
rect 562402 1005193 562430 1005239
rect 571888 1005227 571894 1005239
rect 571946 1005227 571952 1005279
rect 553802 1005165 562430 1005193
rect 553802 1005153 553808 1005165
rect 562480 1005153 562486 1005205
rect 562538 1005193 562544 1005205
rect 572944 1005193 572950 1005205
rect 562538 1005165 572950 1005193
rect 562538 1005153 562544 1005165
rect 572944 1005153 572950 1005165
rect 573002 1005153 573008 1005205
rect 440810 1005091 441086 1005119
rect 440810 1005079 440816 1005091
rect 434704 1005005 434710 1005057
rect 434762 1005045 434768 1005057
rect 437200 1005045 437206 1005057
rect 434762 1005017 437206 1005045
rect 434762 1005005 434768 1005017
rect 437200 1005005 437206 1005017
rect 437258 1005005 437264 1005057
rect 100720 1004931 100726 1004983
rect 100778 1004971 100784 1004983
rect 114160 1004971 114166 1004983
rect 100778 1004943 114166 1004971
rect 100778 1004931 100784 1004943
rect 114160 1004931 114166 1004943
rect 114218 1004931 114224 1004983
rect 512656 1004857 512662 1004909
rect 512714 1004897 512720 1004909
rect 521200 1004897 521206 1004909
rect 512714 1004869 521206 1004897
rect 512714 1004857 512720 1004869
rect 521200 1004857 521206 1004869
rect 521258 1004857 521264 1004909
rect 356752 1003895 356758 1003947
rect 356810 1003935 356816 1003947
rect 377200 1003935 377206 1003947
rect 356810 1003907 377206 1003935
rect 356810 1003895 356816 1003907
rect 377200 1003895 377206 1003907
rect 377258 1003895 377264 1003947
rect 359056 1003821 359062 1003873
rect 359114 1003861 359120 1003873
rect 379984 1003861 379990 1003873
rect 359114 1003833 379990 1003861
rect 359114 1003821 359120 1003833
rect 379984 1003821 379990 1003833
rect 380042 1003821 380048 1003873
rect 428080 1003821 428086 1003873
rect 428138 1003861 428144 1003873
rect 466480 1003861 466486 1003873
rect 428138 1003833 466486 1003861
rect 428138 1003821 428144 1003833
rect 466480 1003821 466486 1003833
rect 466538 1003821 466544 1003873
rect 501136 1003821 501142 1003873
rect 501194 1003861 501200 1003873
rect 519472 1003861 519478 1003873
rect 501194 1003833 519478 1003861
rect 501194 1003821 501200 1003833
rect 519472 1003821 519478 1003833
rect 519530 1003821 519536 1003873
rect 551728 1003821 551734 1003873
rect 551786 1003861 551792 1003873
rect 570640 1003861 570646 1003873
rect 551786 1003833 570646 1003861
rect 551786 1003821 551792 1003833
rect 570640 1003821 570646 1003833
rect 570698 1003821 570704 1003873
rect 355984 1003747 355990 1003799
rect 356042 1003787 356048 1003799
rect 377104 1003787 377110 1003799
rect 356042 1003759 377110 1003787
rect 356042 1003747 356048 1003759
rect 377104 1003747 377110 1003759
rect 377162 1003747 377168 1003799
rect 423376 1003747 423382 1003799
rect 423434 1003787 423440 1003799
rect 469264 1003787 469270 1003799
rect 423434 1003759 469270 1003787
rect 423434 1003747 423440 1003759
rect 469264 1003747 469270 1003759
rect 469322 1003747 469328 1003799
rect 556528 1003747 556534 1003799
rect 556586 1003787 556592 1003799
rect 574480 1003787 574486 1003799
rect 556586 1003759 574486 1003787
rect 556586 1003747 556592 1003759
rect 574480 1003747 574486 1003759
rect 574538 1003747 574544 1003799
rect 195280 1003673 195286 1003725
rect 195338 1003713 195344 1003725
rect 211696 1003713 211702 1003725
rect 195338 1003685 211702 1003713
rect 195338 1003673 195344 1003685
rect 211696 1003673 211702 1003685
rect 211754 1003673 211760 1003725
rect 359920 1003673 359926 1003725
rect 359978 1003713 359984 1003725
rect 380080 1003713 380086 1003725
rect 359978 1003685 380086 1003713
rect 359978 1003673 359984 1003685
rect 380080 1003673 380086 1003685
rect 380138 1003673 380144 1003725
rect 426448 1003673 426454 1003725
rect 426506 1003713 426512 1003725
rect 470128 1003713 470134 1003725
rect 426506 1003685 470134 1003713
rect 426506 1003673 426512 1003685
rect 470128 1003673 470134 1003685
rect 470186 1003673 470192 1003725
rect 500368 1003673 500374 1003725
rect 500426 1003713 500432 1003725
rect 521008 1003713 521014 1003725
rect 500426 1003685 521014 1003713
rect 500426 1003673 500432 1003685
rect 521008 1003673 521014 1003685
rect 521066 1003673 521072 1003725
rect 552592 1003673 552598 1003725
rect 552650 1003713 552656 1003725
rect 573040 1003713 573046 1003725
rect 552650 1003685 573046 1003713
rect 552650 1003673 552656 1003685
rect 573040 1003673 573046 1003685
rect 573098 1003673 573104 1003725
rect 144208 1002563 144214 1002615
rect 144266 1002603 144272 1002615
rect 151504 1002603 151510 1002615
rect 144266 1002575 151510 1002603
rect 144266 1002563 144272 1002575
rect 151504 1002563 151510 1002575
rect 151562 1002563 151568 1002615
rect 143728 1002489 143734 1002541
rect 143786 1002529 143792 1002541
rect 152848 1002529 152854 1002541
rect 143786 1002501 152854 1002529
rect 143786 1002489 143792 1002501
rect 152848 1002489 152854 1002501
rect 152906 1002489 152912 1002541
rect 502768 1002489 502774 1002541
rect 502826 1002529 502832 1002541
rect 515440 1002529 515446 1002541
rect 502826 1002501 515446 1002529
rect 502826 1002489 502832 1002501
rect 515440 1002489 515446 1002501
rect 515498 1002489 515504 1002541
rect 559120 1002489 559126 1002541
rect 559178 1002529 559184 1002541
rect 566128 1002529 566134 1002541
rect 559178 1002501 566134 1002529
rect 559178 1002489 559184 1002501
rect 566128 1002489 566134 1002501
rect 566186 1002489 566192 1002541
rect 143920 1002415 143926 1002467
rect 143978 1002455 143984 1002467
rect 153616 1002455 153622 1002467
rect 143978 1002427 153622 1002455
rect 143978 1002415 143984 1002427
rect 153616 1002415 153622 1002427
rect 153674 1002415 153680 1002467
rect 489520 1002415 489526 1002467
rect 489578 1002455 489584 1002467
rect 489578 1002427 502142 1002455
rect 489578 1002415 489584 1002427
rect 144016 1002341 144022 1002393
rect 144074 1002381 144080 1002393
rect 150352 1002381 150358 1002393
rect 144074 1002353 150358 1002381
rect 144074 1002341 144080 1002353
rect 150352 1002341 150358 1002353
rect 150410 1002341 150416 1002393
rect 502114 1002381 502142 1002427
rect 503440 1002415 503446 1002467
rect 503498 1002455 503504 1002467
rect 513520 1002455 513526 1002467
rect 503498 1002427 513526 1002455
rect 503498 1002415 503504 1002427
rect 513520 1002415 513526 1002427
rect 513578 1002415 513584 1002467
rect 559888 1002415 559894 1002467
rect 559946 1002455 559952 1002467
rect 564496 1002455 564502 1002467
rect 559946 1002427 564502 1002455
rect 559946 1002415 559952 1002427
rect 564496 1002415 564502 1002427
rect 564554 1002415 564560 1002467
rect 518608 1002381 518614 1002393
rect 502114 1002353 518614 1002381
rect 518608 1002341 518614 1002353
rect 518666 1002341 518672 1002393
rect 560560 1002341 560566 1002393
rect 560618 1002381 560624 1002393
rect 564688 1002381 564694 1002393
rect 560618 1002353 564694 1002381
rect 560618 1002341 560624 1002353
rect 564688 1002341 564694 1002353
rect 564746 1002341 564752 1002393
rect 564784 1002341 564790 1002393
rect 564842 1002381 564848 1002393
rect 568720 1002381 568726 1002393
rect 564842 1002353 568726 1002381
rect 564842 1002341 564848 1002353
rect 568720 1002341 568726 1002353
rect 568778 1002341 568784 1002393
rect 144304 1002267 144310 1002319
rect 144362 1002307 144368 1002319
rect 178480 1002307 178486 1002319
rect 144362 1002279 178486 1002307
rect 144362 1002267 144368 1002279
rect 178480 1002267 178486 1002279
rect 178538 1002267 178544 1002319
rect 505072 1002267 505078 1002319
rect 505130 1002307 505136 1002319
rect 521488 1002307 521494 1002319
rect 505130 1002279 521494 1002307
rect 505130 1002267 505136 1002279
rect 521488 1002267 521494 1002279
rect 521546 1002267 521552 1002319
rect 561520 1002267 561526 1002319
rect 561578 1002307 561584 1002319
rect 565360 1002307 565366 1002319
rect 561578 1002279 565366 1002307
rect 561578 1002267 561584 1002279
rect 565360 1002267 565366 1002279
rect 565418 1002267 565424 1002319
rect 573040 1002193 573046 1002245
rect 573098 1002233 573104 1002245
rect 573328 1002233 573334 1002245
rect 573098 1002205 573334 1002233
rect 573098 1002193 573104 1002205
rect 573328 1002193 573334 1002205
rect 573386 1002193 573392 1002245
rect 452944 1002045 452950 1002097
rect 453002 1002085 453008 1002097
rect 461584 1002085 461590 1002097
rect 453002 1002057 461590 1002085
rect 453002 1002045 453008 1002057
rect 461584 1002045 461590 1002057
rect 461642 1002045 461648 1002097
rect 469360 1002045 469366 1002097
rect 469418 1002085 469424 1002097
rect 472144 1002085 472150 1002097
rect 469418 1002057 472150 1002085
rect 469418 1002045 469424 1002057
rect 472144 1002045 472150 1002057
rect 472202 1002045 472208 1002097
rect 566128 1001601 566134 1001653
rect 566186 1001641 566192 1001653
rect 570160 1001641 570166 1001653
rect 566186 1001613 570166 1001641
rect 566186 1001601 566192 1001613
rect 570160 1001601 570166 1001613
rect 570218 1001601 570224 1001653
rect 513520 1001453 513526 1001505
rect 513578 1001493 513584 1001505
rect 515728 1001493 515734 1001505
rect 513578 1001465 515734 1001493
rect 513578 1001453 513584 1001465
rect 515728 1001453 515734 1001465
rect 515786 1001453 515792 1001505
rect 572848 1001453 572854 1001505
rect 572906 1001493 572912 1001505
rect 574096 1001493 574102 1001505
rect 572906 1001465 574102 1001493
rect 572906 1001453 572912 1001465
rect 574096 1001453 574102 1001465
rect 574154 1001453 574160 1001505
rect 434032 1001083 434038 1001135
rect 434090 1001123 434096 1001135
rect 472624 1001123 472630 1001135
rect 434090 1001095 472630 1001123
rect 434090 1001083 434096 1001095
rect 472624 1001083 472630 1001095
rect 472682 1001083 472688 1001135
rect 432496 1001009 432502 1001061
rect 432554 1001049 432560 1001061
rect 472528 1001049 472534 1001061
rect 432554 1001021 472534 1001049
rect 432554 1001009 432560 1001021
rect 472528 1001009 472534 1001021
rect 472586 1001009 472592 1001061
rect 564496 1001009 564502 1001061
rect 564554 1001049 564560 1001061
rect 567760 1001049 567766 1001061
rect 564554 1001021 567766 1001049
rect 564554 1001009 564560 1001021
rect 567760 1001009 567766 1001021
rect 567818 1001009 567824 1001061
rect 571888 1001009 571894 1001061
rect 571946 1001049 571952 1001061
rect 573232 1001049 573238 1001061
rect 571946 1001021 573238 1001049
rect 571946 1001009 571952 1001021
rect 573232 1001009 573238 1001021
rect 573290 1001009 573296 1001061
rect 430864 1000935 430870 1000987
rect 430922 1000975 430928 1000987
rect 472336 1000975 472342 1000987
rect 430922 1000947 472342 1000975
rect 430922 1000935 430928 1000947
rect 472336 1000935 472342 1000947
rect 472394 1000935 472400 1000987
rect 510928 1000935 510934 1000987
rect 510986 1000975 510992 1000987
rect 516688 1000975 516694 1000987
rect 510986 1000947 516694 1000975
rect 510986 1000935 510992 1000947
rect 516688 1000935 516694 1000947
rect 516746 1000935 516752 1000987
rect 195088 1000861 195094 1000913
rect 195146 1000901 195152 1000913
rect 208144 1000901 208150 1000913
rect 195146 1000873 208150 1000901
rect 195146 1000861 195152 1000873
rect 208144 1000861 208150 1000873
rect 208202 1000861 208208 1000913
rect 428944 1000861 428950 1000913
rect 429002 1000901 429008 1000913
rect 472624 1000901 472630 1000913
rect 429002 1000873 472630 1000901
rect 429002 1000861 429008 1000873
rect 472624 1000861 472630 1000873
rect 472682 1000861 472688 1000913
rect 143824 1000787 143830 1000839
rect 143882 1000827 143888 1000839
rect 160240 1000827 160246 1000839
rect 143882 1000799 160246 1000827
rect 143882 1000787 143888 1000799
rect 160240 1000787 160246 1000799
rect 160298 1000787 160304 1000839
rect 361552 1000787 361558 1000839
rect 361610 1000827 361616 1000839
rect 383632 1000827 383638 1000839
rect 361610 1000799 383638 1000827
rect 361610 1000787 361616 1000799
rect 383632 1000787 383638 1000799
rect 383690 1000787 383696 1000839
rect 427312 1000787 427318 1000839
rect 427370 1000827 427376 1000839
rect 472432 1000827 472438 1000839
rect 427370 1000799 472438 1000827
rect 427370 1000787 427376 1000799
rect 472432 1000787 472438 1000799
rect 472490 1000787 472496 1000839
rect 509296 1000787 509302 1000839
rect 509354 1000827 509360 1000839
rect 516688 1000827 516694 1000839
rect 509354 1000799 516694 1000827
rect 509354 1000787 509360 1000799
rect 516688 1000787 516694 1000799
rect 516746 1000787 516752 1000839
rect 469168 1000713 469174 1000765
rect 469226 1000753 469232 1000765
rect 469552 1000753 469558 1000765
rect 469226 1000725 469558 1000753
rect 469226 1000713 469232 1000725
rect 469552 1000713 469558 1000725
rect 469610 1000713 469616 1000765
rect 298192 1000343 298198 1000395
rect 298250 1000383 298256 1000395
rect 305296 1000383 305302 1000395
rect 298250 1000355 305302 1000383
rect 298250 1000343 298256 1000355
rect 305296 1000343 305302 1000355
rect 305354 1000343 305360 1000395
rect 613456 999825 613462 999877
rect 613514 999865 613520 999877
rect 625552 999865 625558 999877
rect 613514 999837 625558 999865
rect 613514 999825 613520 999837
rect 625552 999825 625558 999837
rect 625610 999825 625616 999877
rect 610576 999751 610582 999803
rect 610634 999791 610640 999803
rect 625456 999791 625462 999803
rect 610634 999763 625462 999791
rect 610634 999751 610640 999763
rect 625456 999751 625462 999763
rect 625514 999751 625520 999803
rect 601840 999677 601846 999729
rect 601898 999717 601904 999729
rect 625840 999717 625846 999729
rect 601898 999689 625846 999717
rect 601898 999677 601904 999689
rect 625840 999677 625846 999689
rect 625898 999677 625904 999729
rect 379120 999603 379126 999655
rect 379178 999643 379184 999655
rect 381424 999643 381430 999655
rect 379178 999615 381430 999643
rect 379178 999603 379184 999615
rect 381424 999603 381430 999615
rect 381482 999603 381488 999655
rect 596176 999603 596182 999655
rect 596234 999643 596240 999655
rect 625744 999643 625750 999655
rect 596234 999615 625750 999643
rect 596234 999603 596240 999615
rect 625744 999603 625750 999615
rect 625802 999603 625808 999655
rect 246640 999529 246646 999581
rect 246698 999569 246704 999581
rect 260752 999569 260758 999581
rect 246698 999541 260758 999569
rect 246698 999529 246704 999541
rect 260752 999529 260758 999541
rect 260810 999529 260816 999581
rect 590704 999529 590710 999581
rect 590762 999569 590768 999581
rect 625360 999569 625366 999581
rect 590762 999541 625366 999569
rect 590762 999529 590768 999541
rect 625360 999529 625366 999541
rect 625418 999529 625424 999581
rect 144112 999455 144118 999507
rect 144170 999495 144176 999507
rect 155152 999495 155158 999507
rect 144170 999467 155158 999495
rect 144170 999455 144176 999467
rect 155152 999455 155158 999467
rect 155210 999455 155216 999507
rect 247696 999455 247702 999507
rect 247754 999495 247760 999507
rect 258832 999495 258838 999507
rect 247754 999467 258838 999495
rect 247754 999455 247760 999467
rect 258832 999455 258838 999467
rect 258890 999455 258896 999507
rect 497584 999455 497590 999507
rect 497642 999495 497648 999507
rect 516688 999495 516694 999507
rect 497642 999467 516694 999495
rect 497642 999455 497648 999467
rect 516688 999455 516694 999467
rect 516746 999455 516752 999507
rect 565360 999455 565366 999507
rect 565418 999495 565424 999507
rect 565418 999467 570398 999495
rect 565418 999455 565424 999467
rect 61840 999381 61846 999433
rect 61898 999421 61904 999433
rect 74704 999421 74710 999433
rect 61898 999393 74710 999421
rect 61898 999381 61904 999393
rect 74704 999381 74710 999393
rect 74762 999381 74768 999433
rect 92944 999381 92950 999433
rect 93002 999421 93008 999433
rect 123856 999421 123862 999433
rect 93002 999393 123862 999421
rect 93002 999381 93008 999393
rect 123856 999381 123862 999393
rect 123914 999381 123920 999433
rect 143728 999381 143734 999433
rect 143786 999421 143792 999433
rect 156880 999421 156886 999433
rect 143786 999393 156886 999421
rect 143786 999381 143792 999393
rect 156880 999381 156886 999393
rect 156938 999381 156944 999433
rect 195184 999381 195190 999433
rect 195242 999421 195248 999433
rect 226000 999421 226006 999433
rect 195242 999393 226006 999421
rect 195242 999381 195248 999393
rect 226000 999381 226006 999393
rect 226058 999381 226064 999433
rect 246544 999381 246550 999433
rect 246602 999421 246608 999433
rect 259600 999421 259606 999433
rect 246602 999393 259606 999421
rect 246602 999381 246608 999393
rect 259600 999381 259606 999393
rect 259658 999381 259664 999433
rect 298096 999381 298102 999433
rect 298154 999421 298160 999433
rect 311248 999421 311254 999433
rect 298154 999393 311254 999421
rect 298154 999381 298160 999393
rect 311248 999381 311254 999393
rect 311306 999381 311312 999433
rect 377104 999381 377110 999433
rect 377162 999421 377168 999433
rect 379024 999421 379030 999433
rect 377162 999393 379030 999421
rect 377162 999381 377168 999393
rect 379024 999381 379030 999393
rect 379082 999381 379088 999433
rect 466576 999381 466582 999433
rect 466634 999421 466640 999433
rect 472240 999421 472246 999433
rect 466634 999393 472246 999421
rect 466634 999381 466640 999393
rect 472240 999381 472246 999393
rect 472298 999381 472304 999433
rect 540304 999381 540310 999433
rect 540362 999421 540368 999433
rect 570256 999421 570262 999433
rect 540362 999393 570262 999421
rect 540362 999381 540368 999393
rect 570256 999381 570262 999393
rect 570314 999381 570320 999433
rect 506320 999307 506326 999359
rect 506378 999347 506384 999359
rect 516688 999347 516694 999359
rect 506378 999319 516694 999347
rect 506378 999307 506384 999319
rect 516688 999307 516694 999319
rect 516746 999307 516752 999359
rect 570370 999347 570398 999467
rect 590608 999455 590614 999507
rect 590666 999495 590672 999507
rect 625840 999495 625846 999507
rect 590666 999467 625846 999495
rect 590666 999455 590672 999467
rect 625840 999455 625846 999467
rect 625898 999455 625904 999507
rect 590512 999381 590518 999433
rect 590570 999421 590576 999433
rect 625648 999421 625654 999433
rect 590570 999393 625654 999421
rect 590570 999381 590576 999393
rect 625648 999381 625654 999393
rect 625706 999381 625712 999433
rect 571024 999347 571030 999359
rect 570370 999319 571030 999347
rect 571024 999307 571030 999319
rect 571082 999307 571088 999359
rect 461584 998715 461590 998767
rect 461642 998755 461648 998767
rect 466576 998755 466582 998767
rect 461642 998727 466582 998755
rect 461642 998715 461648 998727
rect 466576 998715 466582 998727
rect 466634 998715 466640 998767
rect 567760 998567 567766 998619
rect 567818 998607 567824 998619
rect 570832 998607 570838 998619
rect 567818 998579 570838 998607
rect 567818 998567 567824 998579
rect 570832 998567 570838 998579
rect 570890 998567 570896 998619
rect 195376 997901 195382 997953
rect 195434 997941 195440 997953
rect 209392 997941 209398 997953
rect 195434 997913 209398 997941
rect 195434 997901 195440 997913
rect 209392 997901 209398 997913
rect 209450 997901 209456 997953
rect 328336 997901 328342 997953
rect 328394 997941 328400 997953
rect 367888 997941 367894 997953
rect 328394 997913 367894 997941
rect 328394 997901 328400 997913
rect 367888 997901 367894 997913
rect 367946 997941 367952 997953
rect 371440 997941 371446 997953
rect 367946 997913 371446 997941
rect 367946 997901 367952 997913
rect 371440 997901 371446 997913
rect 371498 997901 371504 997953
rect 555184 997901 555190 997953
rect 555242 997941 555248 997953
rect 559888 997941 559894 997953
rect 555242 997913 559894 997941
rect 555242 997901 555248 997913
rect 559888 997901 559894 997913
rect 559946 997901 559952 997953
rect 570256 997901 570262 997953
rect 570314 997941 570320 997953
rect 610672 997941 610678 997953
rect 570314 997913 610678 997941
rect 570314 997901 570320 997913
rect 610672 997901 610678 997913
rect 610730 997901 610736 997953
rect 325456 997827 325462 997879
rect 325514 997867 325520 997879
rect 350128 997867 350134 997879
rect 325514 997839 350134 997867
rect 325514 997827 325520 997839
rect 350128 997827 350134 997839
rect 350186 997827 350192 997879
rect 557296 997827 557302 997879
rect 557354 997867 557360 997879
rect 596176 997867 596182 997879
rect 557354 997839 596182 997867
rect 557354 997827 557360 997839
rect 596176 997827 596182 997839
rect 596234 997827 596240 997879
rect 318448 997753 318454 997805
rect 318506 997793 318512 997805
rect 369040 997793 369046 997805
rect 318506 997765 369046 997793
rect 318506 997753 318512 997765
rect 369040 997753 369046 997765
rect 369098 997753 369104 997805
rect 556144 997753 556150 997805
rect 556202 997793 556208 997805
rect 590512 997793 590518 997805
rect 556202 997765 590518 997793
rect 556202 997753 556208 997765
rect 590512 997753 590518 997765
rect 590570 997753 590576 997805
rect 564688 997679 564694 997731
rect 564746 997719 564752 997731
rect 590608 997719 590614 997731
rect 564746 997691 590614 997719
rect 564746 997679 564752 997691
rect 590608 997679 590614 997691
rect 590666 997679 590672 997731
rect 573328 997605 573334 997657
rect 573386 997645 573392 997657
rect 590704 997645 590710 997657
rect 573386 997617 590710 997645
rect 573386 997605 573392 997617
rect 590704 997605 590710 997617
rect 590762 997605 590768 997657
rect 573232 997531 573238 997583
rect 573290 997571 573296 997583
rect 610576 997571 610582 997583
rect 573290 997543 610582 997571
rect 573290 997531 573296 997543
rect 610576 997531 610582 997543
rect 610634 997531 610640 997583
rect 559888 997457 559894 997509
rect 559946 997497 559952 997509
rect 570544 997497 570550 997509
rect 559946 997469 570550 997497
rect 559946 997457 559952 997469
rect 570544 997457 570550 997469
rect 570602 997457 570608 997509
rect 572944 997457 572950 997509
rect 573002 997497 573008 997509
rect 601840 997497 601846 997509
rect 573002 997469 601846 997497
rect 573002 997457 573008 997469
rect 601840 997457 601846 997469
rect 601898 997457 601904 997509
rect 574480 997383 574486 997435
rect 574538 997423 574544 997435
rect 613456 997423 613462 997435
rect 574538 997395 613462 997423
rect 574538 997383 574544 997395
rect 613456 997383 613462 997395
rect 613514 997383 613520 997435
rect 377200 997087 377206 997139
rect 377258 997127 377264 997139
rect 382000 997127 382006 997139
rect 377258 997099 382006 997127
rect 377258 997087 377264 997099
rect 382000 997087 382006 997099
rect 382058 997087 382064 997139
rect 510256 996569 510262 996621
rect 510314 996609 510320 996621
rect 521104 996609 521110 996621
rect 510314 996581 521110 996609
rect 510314 996569 510320 996581
rect 521104 996569 521110 996581
rect 521162 996569 521168 996621
rect 259120 996495 259126 996547
rect 259178 996535 259184 996547
rect 263920 996535 263926 996547
rect 259178 996507 263926 996535
rect 259178 996495 259184 996507
rect 263920 996495 263926 996507
rect 263978 996495 263984 996547
rect 379984 996495 379990 996547
rect 380042 996535 380048 996547
rect 380272 996535 380278 996547
rect 380042 996507 380278 996535
rect 380042 996495 380048 996507
rect 380272 996495 380278 996507
rect 380330 996495 380336 996547
rect 507856 996495 507862 996547
rect 507914 996535 507920 996547
rect 521200 996535 521206 996547
rect 507914 996507 521206 996535
rect 507914 996495 507920 996507
rect 521200 996495 521206 996507
rect 521258 996495 521264 996547
rect 316336 996421 316342 996473
rect 316394 996461 316400 996473
rect 316394 996433 328382 996461
rect 316394 996421 316400 996433
rect 328354 996387 328382 996433
rect 328354 996359 348446 996387
rect 162640 996125 162646 996177
rect 162698 996165 162704 996177
rect 213328 996165 213334 996177
rect 162698 996137 213334 996165
rect 162698 996125 162704 996137
rect 213328 996125 213334 996137
rect 213386 996165 213392 996177
rect 265072 996165 265078 996177
rect 213386 996137 265078 996165
rect 213386 996125 213392 996137
rect 265072 996125 265078 996137
rect 265130 996165 265136 996177
rect 276496 996165 276502 996177
rect 265130 996137 276502 996165
rect 265130 996125 265136 996137
rect 276496 996125 276502 996137
rect 276554 996125 276560 996177
rect 302320 996125 302326 996177
rect 302378 996165 302384 996177
rect 316336 996165 316342 996177
rect 302378 996137 316342 996165
rect 302378 996125 302384 996137
rect 316336 996125 316342 996137
rect 316394 996125 316400 996177
rect 348418 996165 348446 996359
rect 423280 996347 423286 996399
rect 423338 996387 423344 996399
rect 440752 996387 440758 996399
rect 423338 996359 440758 996387
rect 423338 996347 423344 996359
rect 440752 996347 440758 996359
rect 440810 996347 440816 996399
rect 511888 996199 511894 996251
rect 511946 996239 511952 996251
rect 511946 996211 513566 996239
rect 511946 996199 511952 996211
rect 348418 996137 367166 996165
rect 367138 996103 367166 996137
rect 399856 996125 399862 996177
rect 399914 996165 399920 996177
rect 408880 996165 408886 996177
rect 399914 996137 408886 996165
rect 399914 996125 399920 996137
rect 408880 996125 408886 996137
rect 408938 996125 408944 996177
rect 408976 996125 408982 996177
rect 409034 996165 409040 996177
rect 423280 996165 423286 996177
rect 409034 996137 423286 996165
rect 409034 996125 409040 996137
rect 423280 996125 423286 996137
rect 423338 996125 423344 996177
rect 436432 996125 436438 996177
rect 436490 996165 436496 996177
rect 513424 996165 513430 996177
rect 436490 996137 513430 996165
rect 436490 996125 436496 996137
rect 513424 996125 513430 996137
rect 513482 996125 513488 996177
rect 513538 996165 513566 996211
rect 563728 996165 563734 996177
rect 513538 996137 563734 996165
rect 563728 996125 563734 996137
rect 563786 996125 563792 996177
rect 164080 996051 164086 996103
rect 164138 996091 164144 996103
rect 215632 996091 215638 996103
rect 164138 996063 215638 996091
rect 164138 996051 164144 996063
rect 215632 996051 215638 996063
rect 215690 996051 215696 996103
rect 218896 996051 218902 996103
rect 218954 996091 218960 996103
rect 266896 996091 266902 996103
rect 218954 996063 266902 996091
rect 218954 996051 218960 996063
rect 266896 996051 266902 996063
rect 266954 996051 266960 996103
rect 266992 996051 266998 996103
rect 267050 996091 267056 996103
rect 318640 996091 318646 996103
rect 267050 996063 318646 996091
rect 267050 996051 267056 996063
rect 318640 996051 318646 996063
rect 318698 996051 318704 996103
rect 367120 996051 367126 996103
rect 367178 996091 367184 996103
rect 437776 996091 437782 996103
rect 367178 996063 437782 996091
rect 367178 996051 367184 996063
rect 437776 996051 437782 996063
rect 437834 996051 437840 996103
rect 471856 996051 471862 996103
rect 471914 996091 471920 996103
rect 511120 996091 511126 996103
rect 471914 996063 511126 996091
rect 471914 996051 471920 996063
rect 511120 996051 511126 996063
rect 511178 996091 511184 996103
rect 562768 996091 562774 996103
rect 511178 996063 562774 996091
rect 511178 996051 511184 996063
rect 562768 996051 562774 996063
rect 562826 996051 562832 996103
rect 103888 996017 103894 996029
rect 81058 995989 103894 996017
rect 81058 995807 81086 995989
rect 103888 995977 103894 995989
rect 103946 995977 103952 996029
rect 115216 995977 115222 996029
rect 115274 996017 115280 996029
rect 164176 996017 164182 996029
rect 115274 995989 164182 996017
rect 115274 995977 115280 995989
rect 164176 995977 164182 995989
rect 164234 995977 164240 996029
rect 276496 995977 276502 996029
rect 276554 996017 276560 996029
rect 436432 996017 436438 996029
rect 276554 995989 282302 996017
rect 276554 995977 276560 995989
rect 92368 995943 92374 995955
rect 84802 995915 92374 995943
rect 84802 995807 84830 995915
rect 92368 995903 92374 995915
rect 92426 995903 92432 995955
rect 92464 995903 92470 995955
rect 92522 995943 92528 995955
rect 101488 995943 101494 995955
rect 92522 995915 101494 995943
rect 92522 995903 92528 995915
rect 101488 995903 101494 995915
rect 101546 995903 101552 995955
rect 106480 995903 106486 995955
rect 106538 995943 106544 995955
rect 113392 995943 113398 995955
rect 106538 995915 113398 995943
rect 106538 995903 106544 995915
rect 113392 995903 113398 995915
rect 113450 995903 113456 995955
rect 144112 995943 144118 995955
rect 132418 995915 144118 995943
rect 132418 995807 132446 995915
rect 144112 995903 144118 995915
rect 144170 995903 144176 995955
rect 144400 995903 144406 995955
rect 144458 995943 144464 995955
rect 151984 995943 151990 995955
rect 144458 995915 151990 995943
rect 144458 995903 144464 995915
rect 151984 995903 151990 995915
rect 152042 995903 152048 995955
rect 195664 995903 195670 995955
rect 195722 995943 195728 995955
rect 200272 995943 200278 995955
rect 195722 995915 200278 995943
rect 195722 995903 195728 995915
rect 200272 995903 200278 995915
rect 200330 995943 200336 995955
rect 200944 995943 200950 995955
rect 200330 995915 200950 995943
rect 200330 995903 200336 995915
rect 200944 995903 200950 995915
rect 201002 995903 201008 995955
rect 213040 995903 213046 995955
rect 213098 995943 213104 995955
rect 216784 995943 216790 995955
rect 213098 995915 216790 995943
rect 213098 995903 213104 995915
rect 216784 995903 216790 995915
rect 216842 995903 216848 995955
rect 246448 995903 246454 995955
rect 246506 995943 246512 995955
rect 282274 995943 282302 995989
rect 377890 995989 436438 996017
rect 246506 995915 255134 995943
rect 282274 995915 282494 995943
rect 246506 995903 246512 995915
rect 254896 995869 254902 995881
rect 236482 995841 254902 995869
rect 236482 995807 236510 995841
rect 254896 995829 254902 995841
rect 254954 995829 254960 995881
rect 255106 995869 255134 995915
rect 257296 995869 257302 995881
rect 255106 995841 257302 995869
rect 257296 995829 257302 995841
rect 257354 995829 257360 995881
rect 81040 995755 81046 995807
rect 81098 995755 81104 995807
rect 84784 995755 84790 995807
rect 84842 995755 84848 995807
rect 91504 995755 91510 995807
rect 91562 995795 91568 995807
rect 105424 995795 105430 995807
rect 91562 995767 105430 995795
rect 91562 995755 91568 995767
rect 105424 995755 105430 995767
rect 105482 995755 105488 995807
rect 113392 995755 113398 995807
rect 113450 995795 113456 995807
rect 118096 995795 118102 995807
rect 113450 995767 118102 995795
rect 113450 995755 113456 995767
rect 118096 995755 118102 995767
rect 118154 995755 118160 995807
rect 132400 995755 132406 995807
rect 132458 995755 132464 995807
rect 142960 995755 142966 995807
rect 143018 995795 143024 995807
rect 143728 995795 143734 995807
rect 143018 995767 143734 995795
rect 143018 995755 143024 995767
rect 143728 995755 143734 995767
rect 143786 995755 143792 995807
rect 164080 995755 164086 995807
rect 164138 995795 164144 995807
rect 165616 995795 165622 995807
rect 164138 995767 165622 995795
rect 164138 995755 164144 995767
rect 165616 995755 165622 995767
rect 165674 995755 165680 995807
rect 188080 995755 188086 995807
rect 188138 995795 188144 995807
rect 202864 995795 202870 995807
rect 188138 995767 202870 995795
rect 188138 995755 188144 995767
rect 202864 995755 202870 995767
rect 202922 995755 202928 995807
rect 236464 995755 236470 995807
rect 236522 995755 236528 995807
rect 245680 995755 245686 995807
rect 245738 995795 245744 995807
rect 246544 995795 246550 995807
rect 245738 995767 246550 995795
rect 245738 995755 245744 995767
rect 246544 995755 246550 995767
rect 246602 995755 246608 995807
rect 250480 995755 250486 995807
rect 250538 995795 250544 995807
rect 254032 995795 254038 995807
rect 250538 995767 254038 995795
rect 250538 995755 250544 995767
rect 254032 995755 254038 995767
rect 254090 995755 254096 995807
rect 268528 995755 268534 995807
rect 268586 995795 268592 995807
rect 273712 995795 273718 995807
rect 268586 995767 273718 995795
rect 268586 995755 268592 995767
rect 273712 995755 273718 995767
rect 273770 995755 273776 995807
rect 74896 995681 74902 995733
rect 74954 995721 74960 995733
rect 82480 995721 82486 995733
rect 74954 995693 82486 995721
rect 74954 995681 74960 995693
rect 82480 995681 82486 995693
rect 82538 995681 82544 995733
rect 85360 995681 85366 995733
rect 85418 995721 85424 995733
rect 99760 995721 99766 995733
rect 85418 995693 99766 995721
rect 85418 995681 85424 995693
rect 99760 995681 99766 995693
rect 99818 995681 99824 995733
rect 141040 995681 141046 995733
rect 141098 995721 141104 995733
rect 143824 995721 143830 995733
rect 141098 995693 143830 995721
rect 141098 995681 141104 995693
rect 143824 995681 143830 995693
rect 143882 995681 143888 995733
rect 163984 995681 163990 995733
rect 164042 995721 164048 995733
rect 166192 995721 166198 995733
rect 164042 995693 166198 995721
rect 164042 995681 164048 995693
rect 166192 995681 166198 995693
rect 166250 995681 166256 995733
rect 188848 995681 188854 995733
rect 188906 995721 188912 995733
rect 204208 995721 204214 995733
rect 188906 995693 204214 995721
rect 188906 995681 188912 995693
rect 204208 995681 204214 995693
rect 204266 995681 204272 995733
rect 250384 995681 250390 995733
rect 250442 995721 250448 995733
rect 255664 995721 255670 995733
rect 250442 995693 255670 995721
rect 250442 995681 250448 995693
rect 255664 995681 255670 995693
rect 255722 995681 255728 995733
rect 133072 995607 133078 995659
rect 133130 995647 133136 995659
rect 146800 995647 146806 995659
rect 133130 995619 146806 995647
rect 133130 995607 133136 995619
rect 146800 995607 146806 995619
rect 146858 995607 146864 995659
rect 194416 995607 194422 995659
rect 194474 995647 194480 995659
rect 195088 995647 195094 995659
rect 194474 995619 195094 995647
rect 194474 995607 194480 995619
rect 195088 995607 195094 995619
rect 195146 995607 195152 995659
rect 139312 995533 139318 995585
rect 139370 995573 139376 995585
rect 143920 995573 143926 995585
rect 139370 995545 143926 995573
rect 139370 995533 139376 995545
rect 143920 995533 143926 995545
rect 143978 995533 143984 995585
rect 191920 995533 191926 995585
rect 191978 995573 191984 995585
rect 195184 995573 195190 995585
rect 191978 995545 195190 995573
rect 191978 995533 191984 995545
rect 195184 995533 195190 995545
rect 195242 995533 195248 995585
rect 82288 995459 82294 995511
rect 82346 995499 82352 995511
rect 99664 995499 99670 995511
rect 82346 995471 99670 995499
rect 82346 995459 82352 995471
rect 99664 995459 99670 995471
rect 99722 995459 99728 995511
rect 184336 995459 184342 995511
rect 184394 995499 184400 995511
rect 201520 995499 201526 995511
rect 184394 995471 201526 995499
rect 184394 995459 184400 995471
rect 201520 995459 201526 995471
rect 201578 995459 201584 995511
rect 282466 995499 282494 995915
rect 370192 995903 370198 995955
rect 370250 995943 370256 995955
rect 374512 995943 374518 995955
rect 370250 995915 374518 995943
rect 370250 995903 370256 995915
rect 374512 995903 374518 995915
rect 374570 995903 374576 995955
rect 298288 995869 298294 995881
rect 291106 995841 298294 995869
rect 287440 995607 287446 995659
rect 287498 995647 287504 995659
rect 291106 995647 291134 995841
rect 298288 995829 298294 995841
rect 298346 995829 298352 995881
rect 299440 995829 299446 995881
rect 299498 995869 299504 995881
rect 304720 995869 304726 995881
rect 299498 995841 304726 995869
rect 299498 995829 299504 995841
rect 304720 995829 304726 995841
rect 304778 995829 304784 995881
rect 368848 995829 368854 995881
rect 368906 995869 368912 995881
rect 377890 995869 377918 995989
rect 436432 995977 436438 995989
rect 436490 995977 436496 996029
rect 470992 995977 470998 996029
rect 471050 996017 471056 996029
rect 511888 996017 511894 996029
rect 471050 995989 511894 996017
rect 471050 995977 471056 995989
rect 511888 995977 511894 995989
rect 511946 995977 511952 996029
rect 513424 995977 513430 996029
rect 513482 996017 513488 996029
rect 564784 996017 564790 996029
rect 513482 995989 564790 996017
rect 513482 995977 513488 995989
rect 564784 995977 564790 995989
rect 564842 995977 564848 996029
rect 625360 995977 625366 996029
rect 625418 996017 625424 996029
rect 625418 995989 633278 996017
rect 625418 995977 625424 995989
rect 399856 995943 399862 995955
rect 368906 995841 377918 995869
rect 377986 995915 399862 995943
rect 368906 995829 368912 995841
rect 291184 995755 291190 995807
rect 291242 995795 291248 995807
rect 305680 995795 305686 995807
rect 291242 995767 305686 995795
rect 291242 995755 291248 995767
rect 305680 995755 305686 995767
rect 305738 995755 305744 995807
rect 310288 995795 310294 995807
rect 305794 995767 310294 995795
rect 297328 995681 297334 995733
rect 297386 995721 297392 995733
rect 298096 995721 298102 995733
rect 297386 995693 298102 995721
rect 297386 995681 297392 995693
rect 298096 995681 298102 995693
rect 298154 995681 298160 995733
rect 302416 995681 302422 995733
rect 302474 995721 302480 995733
rect 305794 995721 305822 995767
rect 310288 995755 310294 995767
rect 310346 995755 310352 995807
rect 360976 995755 360982 995807
rect 361034 995795 361040 995807
rect 365776 995795 365782 995807
rect 361034 995767 365782 995795
rect 361034 995755 361040 995767
rect 365776 995755 365782 995767
rect 365834 995755 365840 995807
rect 371440 995755 371446 995807
rect 371498 995795 371504 995807
rect 377986 995795 378014 995915
rect 399856 995903 399862 995915
rect 399914 995903 399920 995955
rect 472336 995903 472342 995955
rect 472394 995943 472400 995955
rect 472394 995915 481022 995943
rect 472394 995903 472400 995915
rect 383536 995829 383542 995881
rect 383594 995869 383600 995881
rect 383594 995841 389438 995869
rect 383594 995829 383600 995841
rect 389410 995807 389438 995841
rect 472432 995829 472438 995881
rect 472490 995869 472496 995881
rect 472490 995841 477758 995869
rect 472490 995829 472496 995841
rect 477730 995807 477758 995841
rect 480994 995807 481022 995915
rect 523504 995903 523510 995955
rect 523562 995943 523568 995955
rect 523562 995915 529886 995943
rect 523562 995903 523568 995915
rect 523888 995829 523894 995881
rect 523946 995869 523952 995881
rect 523946 995841 529022 995869
rect 523946 995829 523952 995841
rect 528994 995807 529022 995841
rect 529858 995807 529886 995915
rect 625456 995903 625462 995955
rect 625514 995943 625520 995955
rect 625514 995915 631454 995943
rect 625514 995903 625520 995915
rect 610672 995829 610678 995881
rect 610730 995869 610736 995881
rect 616336 995869 616342 995881
rect 610730 995841 616342 995869
rect 610730 995829 610736 995841
rect 616336 995829 616342 995841
rect 616394 995829 616400 995881
rect 625648 995829 625654 995881
rect 625706 995869 625712 995881
rect 625706 995841 630974 995869
rect 625706 995829 625712 995841
rect 630946 995807 630974 995841
rect 371498 995767 378014 995795
rect 371498 995755 371504 995767
rect 383632 995755 383638 995807
rect 383690 995795 383696 995807
rect 384976 995795 384982 995807
rect 383690 995767 384982 995795
rect 383690 995755 383696 995767
rect 384976 995755 384982 995767
rect 385034 995755 385040 995807
rect 389392 995755 389398 995807
rect 389450 995755 389456 995807
rect 472624 995755 472630 995807
rect 472682 995795 472688 995807
rect 474064 995795 474070 995807
rect 472682 995767 474070 995795
rect 472682 995755 472688 995767
rect 474064 995755 474070 995767
rect 474122 995755 474128 995807
rect 477712 995755 477718 995807
rect 477770 995755 477776 995807
rect 480976 995755 480982 995807
rect 481034 995755 481040 995807
rect 523984 995755 523990 995807
rect 524042 995795 524048 995807
rect 527824 995795 527830 995807
rect 524042 995767 527830 995795
rect 524042 995755 524048 995767
rect 527824 995755 527830 995767
rect 527882 995755 527888 995807
rect 528976 995755 528982 995807
rect 529034 995755 529040 995807
rect 529840 995755 529846 995807
rect 529898 995755 529904 995807
rect 537136 995755 537142 995807
rect 537194 995795 537200 995807
rect 540304 995795 540310 995807
rect 537194 995767 540310 995795
rect 537194 995755 537200 995767
rect 540304 995755 540310 995767
rect 540362 995755 540368 995807
rect 563728 995755 563734 995807
rect 563786 995795 563792 995807
rect 567472 995795 567478 995807
rect 563786 995767 567478 995795
rect 563786 995755 563792 995767
rect 567472 995755 567478 995767
rect 567530 995755 567536 995807
rect 625840 995755 625846 995807
rect 625898 995795 625904 995807
rect 626512 995795 626518 995807
rect 625898 995767 626518 995795
rect 625898 995755 625904 995767
rect 626512 995755 626518 995767
rect 626570 995755 626576 995807
rect 630928 995755 630934 995807
rect 630986 995755 630992 995807
rect 631426 995795 631454 995915
rect 631504 995795 631510 995807
rect 631426 995767 631510 995795
rect 631504 995755 631510 995767
rect 631562 995755 631568 995807
rect 633250 995795 633278 995989
rect 634576 995795 634582 995807
rect 633250 995767 634582 995795
rect 634576 995755 634582 995767
rect 634634 995755 634640 995807
rect 302474 995693 305822 995721
rect 302474 995681 302480 995693
rect 365872 995681 365878 995733
rect 365930 995721 365936 995733
rect 377296 995721 377302 995733
rect 365930 995693 377302 995721
rect 365930 995681 365936 995693
rect 377296 995681 377302 995693
rect 377354 995681 377360 995733
rect 383728 995681 383734 995733
rect 383786 995721 383792 995733
rect 384400 995721 384406 995733
rect 383786 995693 384406 995721
rect 383786 995681 383792 995693
rect 384400 995681 384406 995693
rect 384458 995681 384464 995733
rect 472528 995681 472534 995733
rect 472586 995721 472592 995733
rect 473296 995721 473302 995733
rect 472586 995693 473302 995721
rect 472586 995681 472592 995693
rect 473296 995681 473302 995693
rect 473354 995681 473360 995733
rect 524080 995681 524086 995733
rect 524138 995721 524144 995733
rect 528400 995721 528406 995733
rect 524138 995693 528406 995721
rect 524138 995681 524144 995693
rect 528400 995681 528406 995693
rect 528458 995681 528464 995733
rect 625744 995681 625750 995733
rect 625802 995721 625808 995733
rect 627088 995721 627094 995733
rect 625802 995693 627094 995721
rect 625802 995681 625808 995693
rect 627088 995681 627094 995693
rect 627146 995681 627152 995733
rect 287498 995619 291134 995647
rect 287498 995607 287504 995619
rect 291760 995607 291766 995659
rect 291818 995647 291824 995659
rect 307312 995647 307318 995659
rect 291818 995619 307318 995647
rect 291818 995607 291824 995619
rect 307312 995607 307318 995619
rect 307370 995607 307376 995659
rect 472720 995607 472726 995659
rect 472778 995647 472784 995659
rect 474640 995647 474646 995659
rect 472778 995619 474646 995647
rect 472778 995607 472784 995619
rect 474640 995607 474646 995619
rect 474698 995607 474704 995659
rect 523792 995607 523798 995659
rect 523850 995647 523856 995659
rect 525328 995647 525334 995659
rect 523850 995619 525334 995647
rect 523850 995607 523856 995619
rect 525328 995607 525334 995619
rect 525386 995607 525392 995659
rect 562768 995607 562774 995659
rect 562826 995647 562832 995659
rect 567376 995647 567382 995659
rect 562826 995619 567382 995647
rect 562826 995607 562832 995619
rect 567376 995607 567382 995619
rect 567434 995607 567440 995659
rect 625936 995607 625942 995659
rect 625994 995647 626000 995659
rect 627856 995647 627862 995659
rect 625994 995619 627862 995647
rect 625994 995607 626000 995619
rect 627856 995607 627862 995619
rect 627914 995607 627920 995659
rect 287920 995533 287926 995585
rect 287978 995573 287984 995585
rect 302320 995573 302326 995585
rect 287978 995545 302326 995573
rect 287978 995533 287984 995545
rect 302320 995533 302326 995545
rect 302378 995533 302384 995585
rect 472240 995533 472246 995585
rect 472298 995573 472304 995585
rect 476368 995573 476374 995585
rect 472298 995545 476374 995573
rect 472298 995533 472304 995545
rect 476368 995533 476374 995545
rect 476426 995533 476432 995585
rect 482032 995573 482038 995585
rect 476482 995545 482038 995573
rect 302224 995499 302230 995511
rect 282466 995471 302230 995499
rect 302224 995459 302230 995471
rect 302282 995459 302288 995511
rect 466576 995459 466582 995511
rect 466634 995499 466640 995511
rect 476482 995499 476510 995545
rect 482032 995533 482038 995545
rect 482090 995533 482096 995585
rect 523696 995533 523702 995585
rect 523754 995573 523760 995585
rect 524752 995573 524758 995585
rect 523754 995545 524758 995573
rect 523754 995533 523760 995545
rect 524752 995533 524758 995545
rect 524810 995533 524816 995585
rect 625552 995533 625558 995585
rect 625610 995573 625616 995585
rect 630160 995573 630166 995585
rect 625610 995545 630166 995573
rect 625610 995533 625616 995545
rect 630160 995533 630166 995545
rect 630218 995533 630224 995585
rect 478288 995499 478294 995511
rect 466634 995471 476510 995499
rect 476674 995471 478294 995499
rect 466634 995459 466640 995471
rect 81616 995385 81622 995437
rect 81674 995425 81680 995437
rect 103120 995425 103126 995437
rect 81674 995397 103126 995425
rect 81674 995385 81680 995397
rect 103120 995385 103126 995397
rect 103178 995385 103184 995437
rect 129328 995385 129334 995437
rect 129386 995425 129392 995437
rect 146800 995425 146806 995437
rect 129386 995397 146806 995425
rect 129386 995385 129392 995397
rect 146800 995385 146806 995397
rect 146858 995385 146864 995437
rect 183760 995385 183766 995437
rect 183818 995425 183824 995437
rect 206608 995425 206614 995437
rect 183818 995397 206614 995425
rect 183818 995385 183824 995397
rect 206608 995385 206614 995397
rect 206666 995385 206672 995437
rect 472144 995385 472150 995437
rect 472202 995425 472208 995437
rect 476674 995425 476702 995471
rect 478288 995459 478294 995471
rect 478346 995459 478352 995511
rect 523600 995459 523606 995511
rect 523658 995499 523664 995511
rect 526096 995499 526102 995511
rect 523658 995471 526102 995499
rect 523658 995459 523664 995471
rect 526096 995459 526102 995471
rect 526154 995459 526160 995511
rect 482704 995425 482710 995437
rect 472202 995397 476702 995425
rect 476770 995397 482710 995425
rect 472202 995385 472208 995397
rect 85696 995311 85702 995363
rect 85754 995351 85760 995363
rect 92464 995351 92470 995363
rect 85754 995323 92470 995351
rect 85754 995311 85760 995323
rect 92464 995311 92470 995323
rect 92522 995311 92528 995363
rect 133984 995311 133990 995363
rect 134042 995351 134048 995363
rect 144304 995351 144310 995363
rect 134042 995323 144310 995351
rect 134042 995311 134048 995323
rect 144304 995311 144310 995323
rect 144362 995311 144368 995363
rect 133408 995237 133414 995289
rect 133466 995277 133472 995289
rect 144400 995277 144406 995289
rect 133466 995249 144406 995277
rect 133466 995237 133472 995249
rect 144400 995237 144406 995249
rect 144458 995237 144464 995289
rect 469456 995237 469462 995289
rect 469514 995277 469520 995289
rect 476770 995277 476798 995397
rect 482704 995385 482710 995397
rect 482762 995385 482768 995437
rect 521104 995385 521110 995437
rect 521162 995425 521168 995437
rect 537136 995425 537142 995437
rect 521162 995397 537142 995425
rect 521162 995385 521168 995397
rect 537136 995385 537142 995397
rect 537194 995385 537200 995437
rect 518608 995311 518614 995363
rect 518666 995351 518672 995363
rect 530560 995351 530566 995363
rect 518666 995323 530566 995351
rect 518666 995311 518672 995323
rect 530560 995311 530566 995323
rect 530618 995311 530624 995363
rect 469514 995249 476798 995277
rect 469514 995237 469520 995249
rect 521296 995163 521302 995215
rect 521354 995203 521360 995215
rect 633712 995203 633718 995215
rect 521354 995175 633718 995203
rect 521354 995163 521360 995175
rect 633712 995163 633718 995175
rect 633770 995163 633776 995215
rect 485584 995089 485590 995141
rect 485642 995129 485648 995141
rect 643984 995129 643990 995141
rect 485642 995101 643990 995129
rect 485642 995089 485648 995101
rect 643984 995089 643990 995101
rect 644042 995089 644048 995141
rect 226000 995015 226006 995067
rect 226058 995055 226064 995067
rect 642448 995055 642454 995067
rect 226058 995027 642454 995055
rect 226058 995015 226064 995027
rect 642448 995015 642454 995027
rect 642506 995015 642512 995067
rect 320752 994719 320758 994771
rect 320810 994759 320816 994771
rect 325456 994759 325462 994771
rect 320810 994731 325462 994759
rect 320810 994719 320816 994731
rect 325456 994719 325462 994731
rect 325514 994719 325520 994771
rect 227536 994423 227542 994475
rect 227594 994463 227600 994475
rect 236752 994463 236758 994475
rect 227594 994435 236758 994463
rect 227594 994423 227600 994435
rect 236752 994423 236758 994435
rect 236810 994463 236816 994475
rect 238960 994463 238966 994475
rect 236810 994435 238966 994463
rect 236810 994423 236816 994435
rect 238960 994423 238966 994435
rect 239018 994423 239024 994475
rect 630832 994349 630838 994401
rect 630890 994389 630896 994401
rect 632368 994389 632374 994401
rect 630890 994361 632374 994389
rect 630890 994349 630896 994361
rect 632368 994349 632374 994361
rect 632426 994349 632432 994401
rect 247792 994127 247798 994179
rect 247850 994167 247856 994179
rect 250480 994167 250486 994179
rect 247850 994139 250486 994167
rect 247850 994127 247856 994139
rect 250480 994127 250486 994139
rect 250538 994127 250544 994179
rect 82576 994053 82582 994105
rect 82634 994093 82640 994105
rect 133936 994093 133942 994105
rect 82634 994065 133942 994093
rect 82634 994053 82640 994065
rect 133936 994053 133942 994065
rect 133994 994053 134000 994105
rect 259120 994093 259126 994105
rect 247810 994065 259126 994093
rect 243088 993979 243094 994031
rect 243146 994019 243152 994031
rect 247696 994019 247702 994031
rect 243146 993991 247702 994019
rect 243146 993979 243152 993991
rect 247696 993979 247702 993991
rect 247754 993979 247760 994031
rect 235792 993905 235798 993957
rect 235850 993945 235856 993957
rect 246448 993945 246454 993957
rect 235850 993917 246454 993945
rect 235850 993905 235856 993917
rect 246448 993905 246454 993917
rect 246506 993905 246512 993957
rect 180496 993831 180502 993883
rect 180554 993871 180560 993883
rect 198736 993871 198742 993883
rect 180554 993843 198742 993871
rect 180554 993831 180560 993843
rect 198736 993831 198742 993843
rect 198794 993831 198800 993883
rect 234928 993831 234934 993883
rect 234986 993871 234992 993883
rect 247696 993871 247702 993883
rect 234986 993843 247702 993871
rect 234986 993831 234992 993843
rect 247696 993831 247702 993843
rect 247754 993831 247760 993883
rect 77680 993757 77686 993809
rect 77738 993797 77744 993809
rect 100720 993797 100726 993809
rect 77738 993769 100726 993797
rect 77738 993757 77744 993769
rect 100720 993757 100726 993769
rect 100778 993757 100784 993809
rect 131824 993757 131830 993809
rect 131882 993797 131888 993809
rect 158608 993797 158614 993809
rect 131882 993769 158614 993797
rect 131882 993757 131888 993769
rect 158608 993757 158614 993769
rect 158666 993757 158672 993809
rect 182992 993757 182998 993809
rect 183050 993797 183056 993809
rect 210160 993797 210166 993809
rect 183050 993769 210166 993797
rect 183050 993757 183056 993769
rect 210160 993757 210166 993769
rect 210218 993757 210224 993809
rect 232144 993757 232150 993809
rect 232202 993797 232208 993809
rect 243088 993797 243094 993809
rect 232202 993769 243094 993797
rect 232202 993757 232208 993769
rect 243088 993757 243094 993769
rect 243146 993757 243152 993809
rect 247810 993797 247838 994065
rect 259120 994053 259126 994065
rect 259178 994053 259184 994105
rect 574096 993979 574102 994031
rect 574154 994019 574160 994031
rect 635248 994019 635254 994031
rect 574154 993991 635254 994019
rect 574154 993979 574160 993991
rect 635248 993979 635254 993991
rect 635306 993979 635312 994031
rect 570640 993831 570646 993883
rect 570698 993871 570704 993883
rect 636112 993871 636118 993883
rect 570698 993843 636118 993871
rect 570698 993831 570704 993843
rect 636112 993831 636118 993843
rect 636170 993831 636176 993883
rect 243202 993769 247838 993797
rect 77296 993683 77302 993735
rect 77354 993723 77360 993735
rect 108208 993723 108214 993735
rect 77354 993695 108214 993723
rect 77354 993683 77360 993695
rect 108208 993683 108214 993695
rect 108266 993683 108272 993735
rect 128464 993683 128470 993735
rect 128522 993723 128528 993735
rect 159472 993723 159478 993735
rect 128522 993695 159478 993723
rect 128522 993683 128528 993695
rect 159472 993683 159478 993695
rect 159530 993683 159536 993735
rect 181360 993683 181366 993735
rect 181418 993723 181424 993735
rect 212656 993723 212662 993735
rect 181418 993695 212662 993723
rect 181418 993683 181424 993695
rect 212656 993683 212662 993695
rect 212714 993683 212720 993735
rect 232528 993683 232534 993735
rect 232586 993723 232592 993735
rect 243202 993723 243230 993769
rect 470128 993757 470134 993809
rect 470186 993797 470192 993809
rect 484144 993797 484150 993809
rect 470186 993769 484150 993797
rect 470186 993757 470192 993769
rect 484144 993757 484150 993769
rect 484202 993757 484208 993809
rect 515728 993757 515734 993809
rect 515786 993797 515792 993809
rect 535312 993797 535318 993809
rect 515786 993769 535318 993797
rect 515786 993757 515792 993769
rect 535312 993757 535318 993769
rect 535370 993757 535376 993809
rect 570544 993757 570550 993809
rect 570602 993797 570608 993809
rect 637360 993797 637366 993809
rect 570602 993769 637366 993797
rect 570602 993757 570608 993769
rect 637360 993757 637366 993769
rect 637418 993757 637424 993809
rect 232586 993695 243230 993723
rect 232586 993683 232592 993695
rect 243280 993683 243286 993735
rect 243338 993723 243344 993735
rect 247600 993723 247606 993735
rect 243338 993695 247606 993723
rect 243338 993683 243344 993695
rect 247600 993683 247606 993695
rect 247658 993683 247664 993735
rect 283504 993683 283510 993735
rect 283562 993723 283568 993735
rect 302416 993723 302422 993735
rect 283562 993695 302422 993723
rect 283562 993683 283568 993695
rect 302416 993683 302422 993695
rect 302474 993683 302480 993735
rect 506608 993683 506614 993735
rect 506666 993723 506672 993735
rect 538960 993723 538966 993735
rect 506666 993695 538966 993723
rect 506666 993683 506672 993695
rect 538960 993683 538966 993695
rect 539018 993683 539024 993735
rect 557968 993683 557974 993735
rect 558026 993723 558032 993735
rect 641008 993723 641014 993735
rect 558026 993695 641014 993723
rect 558026 993683 558032 993695
rect 641008 993683 641014 993695
rect 641066 993683 641072 993735
rect 179824 993609 179830 993661
rect 179882 993649 179888 993661
rect 211024 993649 211030 993661
rect 179882 993621 211030 993649
rect 179882 993609 179888 993621
rect 211024 993609 211030 993621
rect 211082 993609 211088 993661
rect 238960 993609 238966 993661
rect 239018 993649 239024 993661
rect 279280 993649 279286 993661
rect 239018 993621 279286 993649
rect 239018 993609 239024 993621
rect 279280 993609 279286 993621
rect 279338 993609 279344 993661
rect 282832 993609 282838 993661
rect 282890 993649 282896 993661
rect 313840 993649 313846 993661
rect 282890 993621 313846 993649
rect 282890 993609 282896 993621
rect 313840 993609 313846 993621
rect 313898 993609 313904 993661
rect 362320 993609 362326 993661
rect 362378 993649 362384 993661
rect 398800 993649 398806 993661
rect 362378 993621 398806 993649
rect 362378 993609 362384 993621
rect 398800 993609 398806 993621
rect 398858 993609 398864 993661
rect 429712 993609 429718 993661
rect 429770 993649 429776 993661
rect 487792 993649 487798 993661
rect 429770 993621 487798 993649
rect 429770 993609 429776 993621
rect 487792 993609 487798 993621
rect 487850 993609 487856 993661
rect 530608 993609 530614 993661
rect 530666 993649 530672 993661
rect 630832 993649 630838 993661
rect 530666 993621 630838 993649
rect 530666 993609 530672 993621
rect 630832 993609 630838 993621
rect 630890 993609 630896 993661
rect 638896 993609 638902 993661
rect 638954 993649 638960 993661
rect 643600 993649 643606 993661
rect 638954 993621 643606 993649
rect 638954 993609 638960 993621
rect 643600 993609 643606 993621
rect 643658 993609 643664 993661
rect 214384 993575 214390 993587
rect 187234 993547 214390 993575
rect 115312 993461 115318 993513
rect 115370 993501 115376 993513
rect 126736 993501 126742 993513
rect 115370 993473 126742 993501
rect 115370 993461 115376 993473
rect 126736 993461 126742 993473
rect 126794 993461 126800 993513
rect 162928 993501 162934 993513
rect 162754 993473 162934 993501
rect 115216 993387 115222 993439
rect 115274 993427 115280 993439
rect 162640 993427 162646 993439
rect 115274 993399 162646 993427
rect 115274 993387 115280 993399
rect 162640 993387 162646 993399
rect 162698 993387 162704 993439
rect 126736 993313 126742 993365
rect 126794 993353 126800 993365
rect 162754 993353 162782 993473
rect 162928 993461 162934 993473
rect 162986 993501 162992 993513
rect 187234 993501 187262 993547
rect 214384 993535 214390 993547
rect 214442 993575 214448 993587
rect 265744 993575 265750 993587
rect 214442 993547 265750 993575
rect 214442 993535 214448 993547
rect 265744 993535 265750 993547
rect 265802 993575 265808 993587
rect 317488 993575 317494 993587
rect 265802 993547 317494 993575
rect 265802 993535 265808 993547
rect 317488 993535 317494 993547
rect 317546 993575 317552 993587
rect 328336 993575 328342 993587
rect 317546 993547 328342 993575
rect 317546 993535 317552 993547
rect 328336 993535 328342 993547
rect 328394 993535 328400 993587
rect 469456 993535 469462 993587
rect 469514 993575 469520 993587
rect 479152 993575 479158 993587
rect 469514 993547 479158 993575
rect 469514 993535 469520 993547
rect 479152 993535 479158 993547
rect 479210 993575 479216 993587
rect 489520 993575 489526 993587
rect 479210 993547 489526 993575
rect 479210 993535 479216 993547
rect 489520 993535 489526 993547
rect 489578 993535 489584 993587
rect 162986 993473 187262 993501
rect 162986 993461 162992 993473
rect 126794 993325 162782 993353
rect 126794 993313 126800 993325
rect 331216 992129 331222 992181
rect 331274 992169 331280 992181
rect 332560 992169 332566 992181
rect 331274 992141 332566 992169
rect 331274 992129 331280 992141
rect 332560 992129 332566 992141
rect 332618 992129 332624 992181
rect 547120 992129 547126 992181
rect 547178 992169 547184 992181
rect 650896 992169 650902 992181
rect 547178 992141 650902 992169
rect 547178 992129 547184 992141
rect 650896 992129 650902 992141
rect 650954 992129 650960 992181
rect 633712 990649 633718 990701
rect 633770 990689 633776 990701
rect 640432 990689 640438 990701
rect 633770 990661 640438 990689
rect 633770 990649 633776 990661
rect 640432 990649 640438 990661
rect 640490 990649 640496 990701
rect 643984 990649 643990 990701
rect 644042 990689 644048 990701
rect 649840 990689 649846 990701
rect 644042 990661 649846 990689
rect 644042 990649 644048 990661
rect 649840 990649 649846 990661
rect 649898 990649 649904 990701
rect 640720 989761 640726 989813
rect 640778 989801 640784 989813
rect 649552 989801 649558 989813
rect 640778 989773 649558 989801
rect 640778 989761 640784 989773
rect 649552 989761 649558 989773
rect 649610 989761 649616 989813
rect 638512 989317 638518 989369
rect 638570 989357 638576 989369
rect 649936 989357 649942 989369
rect 638570 989329 649942 989357
rect 638570 989317 638576 989329
rect 649936 989317 649942 989329
rect 649994 989317 650000 989369
rect 616336 989243 616342 989295
rect 616394 989283 616400 989295
rect 643216 989283 643222 989295
rect 616394 989255 643222 989283
rect 616394 989243 616400 989255
rect 643216 989243 643222 989255
rect 643274 989243 643280 989295
rect 223120 987763 223126 987815
rect 223178 987803 223184 987815
rect 235600 987803 235606 987815
rect 223178 987775 235606 987803
rect 223178 987763 223184 987775
rect 235600 987763 235606 987775
rect 235658 987763 235664 987815
rect 518416 987763 518422 987815
rect 518474 987803 518480 987815
rect 527536 987803 527542 987815
rect 518474 987775 527542 987803
rect 518474 987763 518480 987775
rect 527536 987763 527542 987775
rect 527594 987763 527600 987815
rect 642448 987763 642454 987815
rect 642506 987803 642512 987815
rect 647344 987803 647350 987815
rect 642506 987775 647350 987803
rect 642506 987763 642512 987775
rect 647344 987763 647350 987775
rect 647402 987763 647408 987815
rect 219376 987097 219382 987149
rect 219434 987137 219440 987149
rect 221872 987137 221878 987149
rect 219434 987109 221878 987137
rect 219434 987097 219440 987109
rect 221872 987097 221878 987109
rect 221930 987097 221936 987149
rect 154480 986727 154486 986779
rect 154538 986767 154544 986779
rect 163984 986767 163990 986779
rect 154538 986739 163990 986767
rect 154538 986727 154544 986739
rect 163984 986727 163990 986739
rect 164042 986727 164048 986779
rect 374416 986505 374422 986557
rect 374474 986545 374480 986557
rect 397744 986545 397750 986557
rect 374474 986517 397750 986545
rect 374474 986505 374480 986517
rect 397744 986505 397750 986517
rect 397802 986505 397808 986557
rect 570256 986505 570262 986557
rect 570314 986545 570320 986557
rect 592432 986545 592438 986557
rect 570314 986517 592438 986545
rect 570314 986505 570320 986517
rect 592432 986505 592438 986517
rect 592490 986505 592496 986557
rect 273616 986431 273622 986483
rect 273674 986471 273680 986483
rect 284272 986471 284278 986483
rect 273674 986443 284278 986471
rect 273674 986431 273680 986443
rect 284272 986431 284278 986443
rect 284330 986431 284336 986483
rect 316912 986431 316918 986483
rect 316970 986471 316976 986483
rect 320752 986471 320758 986483
rect 316970 986443 320758 986471
rect 316970 986431 316976 986443
rect 320752 986431 320758 986443
rect 320810 986431 320816 986483
rect 326800 986431 326806 986483
rect 326858 986471 326864 986483
rect 349072 986471 349078 986483
rect 326858 986443 349078 986471
rect 326858 986431 326864 986443
rect 349072 986431 349078 986443
rect 349130 986431 349136 986483
rect 377488 986431 377494 986483
rect 377546 986471 377552 986483
rect 414064 986471 414070 986483
rect 377546 986443 414070 986471
rect 377546 986431 377552 986443
rect 414064 986431 414070 986443
rect 414122 986431 414128 986483
rect 445072 986431 445078 986483
rect 445130 986471 445136 986483
rect 478960 986471 478966 986483
rect 445130 986443 478966 986471
rect 445130 986431 445136 986443
rect 478960 986431 478966 986443
rect 479018 986431 479024 986483
rect 521392 986431 521398 986483
rect 521450 986471 521456 986483
rect 543760 986471 543766 986483
rect 521450 986443 543766 986471
rect 521450 986431 521456 986443
rect 543760 986431 543766 986443
rect 543818 986431 543824 986483
rect 573136 986431 573142 986483
rect 573194 986471 573200 986483
rect 608752 986471 608758 986483
rect 573194 986443 608758 986471
rect 573194 986431 573200 986443
rect 608752 986431 608758 986443
rect 608810 986431 608816 986483
rect 73360 986357 73366 986409
rect 73418 986397 73424 986409
rect 93616 986397 93622 986409
rect 73418 986369 93622 986397
rect 73418 986357 73424 986369
rect 93616 986357 93622 986369
rect 93674 986357 93680 986409
rect 138256 986357 138262 986409
rect 138314 986397 138320 986409
rect 164080 986397 164086 986409
rect 138314 986369 164086 986397
rect 138314 986357 138320 986369
rect 164080 986357 164086 986369
rect 164138 986357 164144 986409
rect 273712 986357 273718 986409
rect 273770 986397 273776 986409
rect 300400 986397 300406 986409
rect 273770 986369 300406 986397
rect 273770 986357 273776 986369
rect 300400 986357 300406 986369
rect 300458 986357 300464 986409
rect 323920 986357 323926 986409
rect 323978 986397 323984 986409
rect 365392 986397 365398 986409
rect 323978 986369 365398 986397
rect 323978 986357 323984 986369
rect 365392 986357 365398 986369
rect 365450 986357 365456 986409
rect 374512 986357 374518 986409
rect 374570 986397 374576 986409
rect 430288 986397 430294 986409
rect 374570 986369 430294 986397
rect 374570 986357 374576 986369
rect 430288 986357 430294 986369
rect 430346 986357 430352 986409
rect 440656 986357 440662 986409
rect 440714 986397 440720 986409
rect 495088 986397 495094 986409
rect 440714 986369 495094 986397
rect 440714 986357 440720 986369
rect 495088 986357 495094 986369
rect 495146 986357 495152 986409
rect 518512 986357 518518 986409
rect 518570 986397 518576 986409
rect 560080 986397 560086 986409
rect 518570 986369 560086 986397
rect 518570 986357 518576 986369
rect 560080 986357 560086 986369
rect 560138 986357 560144 986409
rect 570448 986357 570454 986409
rect 570506 986397 570512 986409
rect 624880 986397 624886 986409
rect 570506 986369 624886 986397
rect 570506 986357 570512 986369
rect 624880 986357 624886 986369
rect 624938 986357 624944 986409
rect 203152 986283 203158 986335
rect 203210 986323 203216 986335
rect 213040 986323 213046 986335
rect 203210 986295 213046 986323
rect 203210 986283 203216 986295
rect 213040 986283 213046 986295
rect 213098 986283 213104 986335
rect 640432 986283 640438 986335
rect 640490 986323 640496 986335
rect 646096 986323 646102 986335
rect 640490 986295 646102 986323
rect 640490 986283 640496 986295
rect 646096 986283 646102 986295
rect 646154 986283 646160 986335
rect 89584 985839 89590 985891
rect 89642 985879 89648 985891
rect 93712 985879 93718 985891
rect 89642 985851 93718 985879
rect 89642 985839 89648 985851
rect 93712 985839 93718 985851
rect 93770 985839 93776 985891
rect 90640 985765 90646 985817
rect 90698 985805 90704 985817
rect 90698 985777 100862 985805
rect 90698 985765 90704 985777
rect 100834 985731 100862 985777
rect 100834 985703 100958 985731
rect 100930 985657 100958 985703
rect 100930 985629 126590 985657
rect 45136 985469 45142 985521
rect 45194 985509 45200 985521
rect 63280 985509 63286 985521
rect 45194 985481 63286 985509
rect 45194 985469 45200 985481
rect 63280 985469 63286 985481
rect 63338 985469 63344 985521
rect 50512 985395 50518 985447
rect 50570 985435 50576 985447
rect 122032 985435 122038 985447
rect 50570 985407 122038 985435
rect 50570 985395 50576 985407
rect 122032 985395 122038 985407
rect 122090 985395 122096 985447
rect 126562 985435 126590 985629
rect 166882 985555 167198 985583
rect 166882 985435 166910 985555
rect 167170 985509 167198 985555
rect 181456 985509 181462 985521
rect 167170 985481 181462 985509
rect 181456 985469 181462 985481
rect 181514 985469 181520 985521
rect 126562 985407 166910 985435
rect 47728 985321 47734 985373
rect 47786 985361 47792 985373
rect 186928 985361 186934 985373
rect 47786 985333 186934 985361
rect 47786 985321 47792 985333
rect 186928 985321 186934 985333
rect 186986 985321 186992 985373
rect 187312 985321 187318 985373
rect 187370 985361 187376 985373
rect 187370 985333 227582 985361
rect 187370 985321 187376 985333
rect 63280 985247 63286 985299
rect 63338 985287 63344 985299
rect 90640 985287 90646 985299
rect 63338 985259 90646 985287
rect 63338 985247 63344 985259
rect 90640 985247 90646 985259
rect 90698 985247 90704 985299
rect 227554 985287 227582 985333
rect 251728 985287 251734 985299
rect 227554 985259 251734 985287
rect 251728 985247 251734 985259
rect 251786 985247 251792 985299
rect 45040 985173 45046 985225
rect 45098 985213 45104 985225
rect 316720 985213 316726 985225
rect 45098 985185 316726 985213
rect 45098 985173 45104 985185
rect 316720 985173 316726 985185
rect 316778 985173 316784 985225
rect 44944 985099 44950 985151
rect 45002 985139 45008 985151
rect 381616 985139 381622 985151
rect 45002 985111 381622 985139
rect 45002 985099 45008 985111
rect 381616 985099 381622 985111
rect 381674 985099 381680 985151
rect 444880 985099 444886 985151
rect 444938 985139 444944 985151
rect 462736 985139 462742 985151
rect 444938 985111 462742 985139
rect 444938 985099 444944 985111
rect 462736 985099 462742 985111
rect 462794 985099 462800 985151
rect 44848 985025 44854 985077
rect 44906 985065 44912 985077
rect 446416 985065 446422 985077
rect 44906 985037 446422 985065
rect 44906 985025 44912 985037
rect 446416 985025 446422 985037
rect 446474 985025 446480 985077
rect 42544 984951 42550 985003
rect 42602 984991 42608 985003
rect 511408 984991 511414 985003
rect 42602 984963 511414 984991
rect 42602 984951 42608 984963
rect 511408 984951 511414 984963
rect 511466 984951 511472 985003
rect 633616 984951 633622 985003
rect 633674 984991 633680 985003
rect 641104 984991 641110 985003
rect 633674 984963 641110 984991
rect 633674 984951 633680 984963
rect 641104 984951 641110 984963
rect 641162 984951 641168 985003
rect 643216 984877 643222 984929
rect 643274 984917 643280 984929
rect 650128 984917 650134 984929
rect 643274 984889 650134 984917
rect 643274 984877 643280 984889
rect 650128 984877 650134 984889
rect 650186 984877 650192 984929
rect 65200 983841 65206 983893
rect 65258 983881 65264 983893
rect 94960 983881 94966 983893
rect 65258 983853 94966 983881
rect 65258 983841 65264 983853
rect 94960 983841 94966 983853
rect 95018 983841 95024 983893
rect 44752 983767 44758 983819
rect 44810 983807 44816 983819
rect 115312 983807 115318 983819
rect 44810 983779 115318 983807
rect 44810 983767 44816 983779
rect 115312 983767 115318 983779
rect 115370 983767 115376 983819
rect 44560 983693 44566 983745
rect 44618 983733 44624 983745
rect 115216 983733 115222 983745
rect 44618 983705 115222 983733
rect 44618 983693 44624 983705
rect 115216 983693 115222 983705
rect 115274 983693 115280 983745
rect 44656 983619 44662 983671
rect 44714 983659 44720 983671
rect 118096 983659 118102 983671
rect 44714 983631 118102 983659
rect 44714 983619 44720 983631
rect 118096 983619 118102 983631
rect 118154 983619 118160 983671
rect 567376 983619 567382 983671
rect 567434 983659 567440 983671
rect 652240 983659 652246 983671
rect 567434 983631 652246 983659
rect 567434 983619 567440 983631
rect 652240 983619 652246 983631
rect 652298 983619 652304 983671
rect 65104 983545 65110 983597
rect 65162 983585 65168 983597
rect 145264 983585 145270 983597
rect 65162 983557 145270 983585
rect 65162 983545 65168 983557
rect 145264 983545 145270 983557
rect 145322 983545 145328 983597
rect 567472 983545 567478 983597
rect 567530 983585 567536 983597
rect 652336 983585 652342 983597
rect 567530 983557 652342 983585
rect 567530 983545 567536 983557
rect 652336 983545 652342 983557
rect 652394 983545 652400 983597
rect 65008 983471 65014 983523
rect 65066 983511 65072 983523
rect 195664 983511 195670 983523
rect 65066 983483 195670 983511
rect 65066 983471 65072 983483
rect 195664 983471 195670 983483
rect 195722 983471 195728 983523
rect 568720 983471 568726 983523
rect 568778 983511 568784 983523
rect 652432 983511 652438 983523
rect 568778 983483 652438 983511
rect 568778 983471 568784 983483
rect 652432 983471 652438 983483
rect 652490 983471 652496 983523
rect 64912 980807 64918 980859
rect 64970 980847 64976 980859
rect 243280 980847 243286 980859
rect 64970 980819 243286 980847
rect 64970 980807 64976 980819
rect 243280 980807 243286 980819
rect 243338 980807 243344 980859
rect 643600 980807 643606 980859
rect 643658 980847 643664 980859
rect 649744 980847 649750 980859
rect 643658 980819 649750 980847
rect 643658 980807 643664 980819
rect 649744 980807 649750 980819
rect 649802 980807 649808 980859
rect 64816 980733 64822 980785
rect 64874 980773 64880 980785
rect 298480 980773 298486 980785
rect 64874 980745 298486 980773
rect 64874 980733 64880 980745
rect 298480 980733 298486 980745
rect 298538 980733 298544 980785
rect 647344 980733 647350 980785
rect 647402 980773 647408 980785
rect 649456 980773 649462 980785
rect 647402 980745 649462 980773
rect 647402 980733 647408 980745
rect 649456 980733 649462 980745
rect 649514 980733 649520 980785
rect 64624 980659 64630 980711
rect 64682 980699 64688 980711
rect 316912 980699 316918 980711
rect 64682 980671 316918 980699
rect 64682 980659 64688 980671
rect 316912 980659 316918 980671
rect 316970 980659 316976 980711
rect 630832 980659 630838 980711
rect 630890 980699 630896 980711
rect 673936 980699 673942 980711
rect 630890 980671 673942 980699
rect 630890 980659 630896 980671
rect 673936 980659 673942 980671
rect 673994 980659 674000 980711
rect 64720 980585 64726 980637
rect 64778 980625 64784 980637
rect 410320 980625 410326 980637
rect 64778 980597 410326 980625
rect 64778 980585 64784 980597
rect 410320 980585 410326 980597
rect 410378 980585 410384 980637
rect 630736 980585 630742 980637
rect 630794 980625 630800 980637
rect 674512 980625 674518 980637
rect 630794 980597 674518 980625
rect 630794 980585 630800 980597
rect 674512 980585 674518 980597
rect 674570 980585 674576 980637
rect 646096 980511 646102 980563
rect 646154 980551 646160 980563
rect 649360 980551 649366 980563
rect 646154 980523 649366 980551
rect 646154 980511 646160 980523
rect 649360 980511 649366 980523
rect 649418 980511 649424 980563
rect 53296 970595 53302 970647
rect 53354 970635 53360 970647
rect 59536 970635 59542 970647
rect 53354 970607 59542 970635
rect 53354 970595 53360 970607
rect 59536 970595 59542 970607
rect 59594 970595 59600 970647
rect 42160 967265 42166 967317
rect 42218 967305 42224 967317
rect 42544 967305 42550 967317
rect 42218 967277 42550 967305
rect 42218 967265 42224 967277
rect 42544 967265 42550 967277
rect 42602 967265 42608 967317
rect 42160 960975 42166 961027
rect 42218 961015 42224 961027
rect 42352 961015 42358 961027
rect 42218 960987 42358 961015
rect 42218 960975 42224 960987
rect 42352 960975 42358 960987
rect 42410 960975 42416 961027
rect 673936 958977 673942 959029
rect 673994 959017 674000 959029
rect 675472 959017 675478 959029
rect 673994 958989 675478 959017
rect 673994 958977 674000 958989
rect 675472 958977 675478 958989
rect 675530 958977 675536 959029
rect 675088 958385 675094 958437
rect 675146 958425 675152 958437
rect 675376 958425 675382 958437
rect 675146 958397 675382 958425
rect 675146 958385 675152 958397
rect 675376 958385 675382 958397
rect 675434 958385 675440 958437
rect 675184 956979 675190 957031
rect 675242 957019 675248 957031
rect 675472 957019 675478 957031
rect 675242 956991 675478 957019
rect 675242 956979 675248 956991
rect 675472 956979 675478 956991
rect 675530 956979 675536 957031
rect 42352 956165 42358 956217
rect 42410 956205 42416 956217
rect 59344 956205 59350 956217
rect 42410 956177 59350 956205
rect 42410 956165 42416 956177
rect 59344 956165 59350 956177
rect 59402 956165 59408 956217
rect 42064 955203 42070 955255
rect 42122 955243 42128 955255
rect 42928 955243 42934 955255
rect 42122 955215 42934 955243
rect 42122 955203 42128 955215
rect 42928 955203 42934 955215
rect 42986 955203 42992 955255
rect 669520 954685 669526 954737
rect 669578 954725 669584 954737
rect 675376 954725 675382 954737
rect 669578 954697 675382 954725
rect 669578 954685 669584 954697
rect 675376 954685 675382 954697
rect 675434 954685 675440 954737
rect 42160 954611 42166 954663
rect 42218 954651 42224 954663
rect 43024 954651 43030 954663
rect 42218 954623 43030 954651
rect 42218 954611 42224 954623
rect 43024 954611 43030 954623
rect 43082 954611 43088 954663
rect 674032 953871 674038 953923
rect 674090 953911 674096 953923
rect 675472 953911 675478 953923
rect 674090 953883 675478 953911
rect 674090 953871 674096 953883
rect 675472 953871 675478 953883
rect 675530 953871 675536 953923
rect 649456 953279 649462 953331
rect 649514 953319 649520 953331
rect 653680 953319 653686 953331
rect 649514 953291 653686 953319
rect 649514 953279 649520 953291
rect 653680 953279 653686 953291
rect 653738 953279 653744 953331
rect 674128 952021 674134 952073
rect 674186 952061 674192 952073
rect 675472 952061 675478 952073
rect 674186 952033 675478 952061
rect 674186 952021 674192 952033
rect 675472 952021 675478 952033
rect 675530 952021 675536 952073
rect 655216 944843 655222 944895
rect 655274 944883 655280 944895
rect 674704 944883 674710 944895
rect 655274 944855 674710 944883
rect 655274 944843 655280 944855
rect 674704 944843 674710 944855
rect 674762 944843 674768 944895
rect 655120 944621 655126 944673
rect 655178 944661 655184 944673
rect 674704 944661 674710 944673
rect 655178 944633 674710 944661
rect 655178 944621 655184 944633
rect 674704 944621 674710 944633
rect 674762 944621 674768 944673
rect 652336 943141 652342 943193
rect 652394 943181 652400 943193
rect 672880 943181 672886 943193
rect 652394 943153 672886 943181
rect 652394 943141 652400 943153
rect 672880 943141 672886 943153
rect 672938 943141 672944 943193
rect 672304 942549 672310 942601
rect 672362 942589 672368 942601
rect 674416 942589 674422 942601
rect 672362 942561 674422 942589
rect 672362 942549 672368 942561
rect 674416 942549 674422 942561
rect 674474 942549 674480 942601
rect 654352 942031 654358 942083
rect 654410 942071 654416 942083
rect 674704 942071 674710 942083
rect 654410 942043 674710 942071
rect 654410 942031 654416 942043
rect 674704 942031 674710 942043
rect 674762 942031 674768 942083
rect 652432 941883 652438 941935
rect 652490 941923 652496 941935
rect 674608 941923 674614 941935
rect 652490 941895 674614 941923
rect 652490 941883 652496 941895
rect 674608 941883 674614 941895
rect 674666 941883 674672 941935
rect 672880 941809 672886 941861
rect 672938 941849 672944 941861
rect 673840 941849 673846 941861
rect 672938 941821 673846 941849
rect 672938 941809 672944 941821
rect 673840 941809 673846 941821
rect 673898 941809 673904 941861
rect 53200 941735 53206 941787
rect 53258 941775 53264 941787
rect 59536 941775 59542 941787
rect 53258 941747 59542 941775
rect 53258 941735 53264 941747
rect 59536 941735 59542 941747
rect 59594 941735 59600 941787
rect 652240 939071 652246 939123
rect 652298 939111 652304 939123
rect 674896 939111 674902 939123
rect 652298 939083 674902 939111
rect 652298 939071 652304 939083
rect 674896 939071 674902 939083
rect 674954 939071 674960 939123
rect 654448 927453 654454 927505
rect 654506 927493 654512 927505
rect 666736 927493 666742 927505
rect 654506 927465 666742 927493
rect 654506 927453 654512 927465
rect 666736 927453 666742 927465
rect 666794 927453 666800 927505
rect 50320 927379 50326 927431
rect 50378 927419 50384 927431
rect 59536 927419 59542 927431
rect 50378 927391 59542 927419
rect 50378 927379 50384 927391
rect 59536 927379 59542 927391
rect 59594 927379 59600 927431
rect 649456 927379 649462 927431
rect 649514 927419 649520 927431
rect 679792 927419 679798 927431
rect 649514 927391 679798 927419
rect 649514 927379 649520 927391
rect 679792 927379 679798 927391
rect 679850 927379 679856 927431
rect 47440 912949 47446 913001
rect 47498 912989 47504 913001
rect 59536 912989 59542 913001
rect 47498 912961 59542 912989
rect 47498 912949 47504 912961
rect 59536 912949 59542 912961
rect 59594 912949 59600 913001
rect 654448 912949 654454 913001
rect 654506 912989 654512 913001
rect 660976 912989 660982 913001
rect 654506 912961 660982 912989
rect 654506 912949 654512 912961
rect 660976 912949 660982 912961
rect 661034 912949 661040 913001
rect 42640 908065 42646 908117
rect 42698 908105 42704 908117
rect 53200 908105 53206 908117
rect 42698 908077 53206 908105
rect 42698 908065 42704 908077
rect 53200 908065 53206 908077
rect 53258 908065 53264 908117
rect 42256 907473 42262 907525
rect 42314 907513 42320 907525
rect 50320 907513 50326 907525
rect 42314 907485 50326 907513
rect 42314 907473 42320 907485
rect 50320 907473 50326 907485
rect 50378 907473 50384 907525
rect 42640 904809 42646 904861
rect 42698 904849 42704 904861
rect 44656 904849 44662 904861
rect 42698 904821 44662 904849
rect 42698 904809 42704 904821
rect 44656 904809 44662 904821
rect 44714 904809 44720 904861
rect 654448 901479 654454 901531
rect 654506 901519 654512 901531
rect 663952 901519 663958 901531
rect 654506 901491 663958 901519
rect 654506 901479 654512 901491
rect 663952 901479 663958 901491
rect 664010 901479 664016 901531
rect 53200 898593 53206 898645
rect 53258 898633 53264 898645
rect 59536 898633 59542 898645
rect 53258 898605 59542 898633
rect 53258 898593 53264 898605
rect 59536 898593 59542 898605
rect 59594 898593 59600 898645
rect 42352 889639 42358 889691
rect 42410 889679 42416 889691
rect 44560 889679 44566 889691
rect 42410 889651 44566 889679
rect 42410 889639 42416 889651
rect 44560 889639 44566 889651
rect 44618 889639 44624 889691
rect 50416 884163 50422 884215
rect 50474 884203 50480 884215
rect 59536 884203 59542 884215
rect 50474 884175 59542 884203
rect 50474 884163 50480 884175
rect 59536 884163 59542 884175
rect 59594 884163 59600 884215
rect 654448 878391 654454 878443
rect 654506 878431 654512 878443
rect 660880 878431 660886 878443
rect 654506 878403 660886 878431
rect 654506 878391 654512 878403
rect 660880 878391 660886 878403
rect 660938 878391 660944 878443
rect 40048 872619 40054 872671
rect 40106 872659 40112 872671
rect 40432 872659 40438 872671
rect 40106 872631 40438 872659
rect 40106 872619 40112 872631
rect 40432 872619 40438 872631
rect 40490 872619 40496 872671
rect 674224 872101 674230 872153
rect 674282 872141 674288 872153
rect 675472 872141 675478 872153
rect 674282 872113 675478 872141
rect 674282 872101 674288 872113
rect 675472 872101 675478 872113
rect 675530 872101 675536 872153
rect 674896 871879 674902 871931
rect 674954 871919 674960 871931
rect 675568 871919 675574 871931
rect 674954 871891 675574 871919
rect 674954 871879 674960 871891
rect 675568 871879 675574 871891
rect 675626 871879 675632 871931
rect 39952 869807 39958 869859
rect 40010 869847 40016 869859
rect 40432 869847 40438 869859
rect 40010 869819 40438 869847
rect 40010 869807 40016 869819
rect 40432 869807 40438 869819
rect 40490 869807 40496 869859
rect 674992 868993 674998 869045
rect 675050 869033 675056 869045
rect 675472 869033 675478 869045
rect 675050 869005 675478 869033
rect 675050 868993 675056 869005
rect 675472 868993 675478 869005
rect 675530 868993 675536 869045
rect 674320 868327 674326 868379
rect 674378 868367 674384 868379
rect 675376 868367 675382 868379
rect 674378 868339 675382 868367
rect 674378 868327 674384 868339
rect 675376 868327 675382 868339
rect 675434 868327 675440 868379
rect 673648 867809 673654 867861
rect 673706 867849 673712 867861
rect 675376 867849 675382 867861
rect 673706 867821 675382 867849
rect 673706 867809 673712 867821
rect 675376 867809 675382 867821
rect 675434 867809 675440 867861
rect 654448 867291 654454 867343
rect 654506 867331 654512 867343
rect 663760 867331 663766 867343
rect 654506 867303 663766 867331
rect 654506 867291 654512 867303
rect 663760 867291 663766 867303
rect 663818 867291 663824 867343
rect 674896 866847 674902 866899
rect 674954 866887 674960 866899
rect 675088 866887 675094 866899
rect 674954 866859 675094 866887
rect 674954 866847 674960 866859
rect 675088 866847 675094 866859
rect 675146 866847 675152 866899
rect 666640 865293 666646 865345
rect 666698 865333 666704 865345
rect 675376 865333 675382 865345
rect 666698 865305 675382 865333
rect 666698 865293 666704 865305
rect 675376 865293 675382 865305
rect 675434 865293 675440 865345
rect 675376 862925 675382 862977
rect 675434 862925 675440 862977
rect 675394 862607 675422 862925
rect 675376 862555 675382 862607
rect 675434 862555 675440 862607
rect 50320 855377 50326 855429
rect 50378 855417 50384 855429
rect 59536 855417 59542 855429
rect 50378 855389 59542 855417
rect 50378 855377 50384 855389
rect 59536 855377 59542 855389
rect 59594 855377 59600 855429
rect 654448 855377 654454 855429
rect 654506 855417 654512 855429
rect 661168 855417 661174 855429
rect 654506 855389 661174 855417
rect 654506 855377 654512 855389
rect 661168 855377 661174 855389
rect 661226 855377 661232 855429
rect 39952 852491 39958 852543
rect 40010 852491 40016 852543
rect 39970 852383 39998 852491
rect 40048 852383 40054 852395
rect 39970 852355 40054 852383
rect 40048 852343 40054 852355
rect 40106 852343 40112 852395
rect 674800 846719 674806 846771
rect 674858 846759 674864 846771
rect 675088 846759 675094 846771
rect 674858 846731 675094 846759
rect 674858 846719 674864 846731
rect 675088 846719 675094 846731
rect 675146 846719 675152 846771
rect 675376 846719 675382 846771
rect 675434 846759 675440 846771
rect 675568 846759 675574 846771
rect 675434 846731 675574 846759
rect 675434 846719 675440 846731
rect 675568 846719 675574 846731
rect 675626 846719 675632 846771
rect 40048 846645 40054 846697
rect 40106 846685 40112 846697
rect 40144 846685 40150 846697
rect 40106 846657 40150 846685
rect 40106 846645 40112 846657
rect 40144 846645 40150 846657
rect 40202 846645 40208 846697
rect 53392 840947 53398 840999
rect 53450 840987 53456 840999
rect 59536 840987 59542 840999
rect 53450 840959 59542 840987
rect 53450 840947 53456 840959
rect 59536 840947 59542 840959
rect 59594 840947 59600 840999
rect 654448 832363 654454 832415
rect 654506 832403 654512 832415
rect 669712 832403 669718 832415
rect 654506 832375 669718 832403
rect 654506 832363 654512 832375
rect 669712 832363 669718 832375
rect 669770 832363 669776 832415
rect 50608 829477 50614 829529
rect 50666 829517 50672 829529
rect 58192 829517 58198 829529
rect 50666 829489 58198 829517
rect 50666 829477 50672 829489
rect 58192 829477 58198 829489
rect 58250 829477 58256 829529
rect 39952 826591 39958 826643
rect 40010 826631 40016 826643
rect 40144 826631 40150 826643
rect 40010 826603 40150 826631
rect 40010 826591 40016 826603
rect 40144 826591 40150 826603
rect 40202 826591 40208 826643
rect 674416 826517 674422 826569
rect 674474 826557 674480 826569
rect 674704 826557 674710 826569
rect 674474 826529 674710 826557
rect 674474 826517 674480 826529
rect 674704 826517 674710 826529
rect 674762 826517 674768 826569
rect 675472 826517 675478 826569
rect 675530 826557 675536 826569
rect 675664 826557 675670 826569
rect 675530 826529 675670 826557
rect 675530 826517 675536 826529
rect 675664 826517 675670 826529
rect 675722 826517 675728 826569
rect 42352 823853 42358 823905
rect 42410 823893 42416 823905
rect 50416 823893 50422 823905
rect 42410 823865 50422 823893
rect 42410 823853 42416 823865
rect 50416 823853 50422 823865
rect 50474 823853 50480 823905
rect 42352 822225 42358 822277
rect 42410 822265 42416 822277
rect 53200 822265 53206 822277
rect 42410 822237 53206 822265
rect 42410 822225 42416 822237
rect 53200 822225 53206 822237
rect 53258 822225 53264 822277
rect 42448 821855 42454 821907
rect 42506 821895 42512 821907
rect 58960 821895 58966 821907
rect 42506 821867 58966 821895
rect 42506 821855 42512 821867
rect 58960 821855 58966 821867
rect 59018 821855 59024 821907
rect 654448 820819 654454 820871
rect 654506 820859 654512 820871
rect 667024 820859 667030 820871
rect 654506 820831 667030 820859
rect 654506 820819 654512 820831
rect 667024 820819 667030 820831
rect 667082 820819 667088 820871
rect 40144 817859 40150 817911
rect 40202 817899 40208 817911
rect 43312 817899 43318 817911
rect 40202 817871 43318 817899
rect 40202 817859 40208 817871
rect 43312 817859 43318 817871
rect 43370 817859 43376 817911
rect 47536 812161 47542 812213
rect 47594 812201 47600 812213
rect 59536 812201 59542 812213
rect 47594 812173 59542 812201
rect 47594 812161 47600 812173
rect 59536 812161 59542 812173
rect 59594 812161 59600 812213
rect 654448 809275 654454 809327
rect 654506 809315 654512 809327
rect 664048 809315 664054 809327
rect 654506 809287 664054 809315
rect 654506 809275 654512 809287
rect 664048 809275 664054 809287
rect 664106 809275 664112 809327
rect 674416 806389 674422 806441
rect 674474 806429 674480 806441
rect 674608 806429 674614 806441
rect 674474 806401 674614 806429
rect 674474 806389 674480 806401
rect 674608 806389 674614 806401
rect 674666 806389 674672 806441
rect 675280 806389 675286 806441
rect 675338 806429 675344 806441
rect 675664 806429 675670 806441
rect 675338 806401 675670 806429
rect 675338 806389 675344 806401
rect 675664 806389 675670 806401
rect 675722 806389 675728 806441
rect 42256 805131 42262 805183
rect 42314 805171 42320 805183
rect 44752 805171 44758 805183
rect 42314 805143 44758 805171
rect 42314 805131 42320 805143
rect 44752 805131 44758 805143
rect 44810 805131 44816 805183
rect 42448 803577 42454 803629
rect 42506 803617 42512 803629
rect 42928 803617 42934 803629
rect 42506 803589 42934 803617
rect 42506 803577 42512 803589
rect 42928 803577 42934 803589
rect 42986 803577 42992 803629
rect 40240 803429 40246 803481
rect 40298 803469 40304 803481
rect 42448 803469 42454 803481
rect 40298 803441 42454 803469
rect 40298 803429 40304 803441
rect 42448 803429 42454 803441
rect 42506 803429 42512 803481
rect 41968 802393 41974 802445
rect 42026 802433 42032 802445
rect 43024 802433 43030 802445
rect 42026 802405 43030 802433
rect 42026 802393 42032 802405
rect 43024 802393 43030 802405
rect 43082 802393 43088 802445
rect 43504 800839 43510 800891
rect 43562 800879 43568 800891
rect 44848 800879 44854 800891
rect 43562 800851 44854 800879
rect 43562 800839 43568 800851
rect 44848 800839 44854 800851
rect 44906 800839 44912 800891
rect 42256 800247 42262 800299
rect 42314 800287 42320 800299
rect 43408 800287 43414 800299
rect 42314 800259 43414 800287
rect 42314 800247 42320 800259
rect 43408 800247 43414 800259
rect 43466 800247 43472 800299
rect 41872 800173 41878 800225
rect 41930 800173 41936 800225
rect 41890 799781 41918 800173
rect 41872 799729 41878 799781
rect 41930 799729 41936 799781
rect 42160 798027 42166 798079
rect 42218 798067 42224 798079
rect 42448 798067 42454 798079
rect 42218 798039 42454 798067
rect 42218 798027 42224 798039
rect 42448 798027 42454 798039
rect 42506 798027 42512 798079
rect 53200 797805 53206 797857
rect 53258 797845 53264 797857
rect 59536 797845 59542 797857
rect 53258 797817 59542 797845
rect 53258 797805 53264 797817
rect 59536 797805 59542 797817
rect 59594 797805 59600 797857
rect 42064 797287 42070 797339
rect 42122 797327 42128 797339
rect 43504 797327 43510 797339
rect 42122 797299 43510 797327
rect 42122 797287 42128 797299
rect 43504 797287 43510 797299
rect 43562 797287 43568 797339
rect 42160 796251 42166 796303
rect 42218 796291 42224 796303
rect 43120 796291 43126 796303
rect 42218 796263 43126 796291
rect 42218 796251 42224 796263
rect 43120 796251 43126 796263
rect 43178 796251 43184 796303
rect 43120 796103 43126 796155
rect 43178 796143 43184 796155
rect 43408 796143 43414 796155
rect 43178 796115 43414 796143
rect 43178 796103 43184 796115
rect 43408 796103 43414 796115
rect 43466 796103 43472 796155
rect 42160 794993 42166 795045
rect 42218 795033 42224 795045
rect 42736 795033 42742 795045
rect 42218 795005 42742 795033
rect 42218 794993 42224 795005
rect 42736 794993 42742 795005
rect 42794 794993 42800 795045
rect 42160 793809 42166 793861
rect 42218 793849 42224 793861
rect 42448 793849 42454 793861
rect 42218 793821 42454 793849
rect 42218 793809 42224 793821
rect 42448 793809 42454 793821
rect 42506 793809 42512 793861
rect 42160 793143 42166 793195
rect 42218 793183 42224 793195
rect 43024 793183 43030 793195
rect 42218 793155 43030 793183
rect 42218 793143 42224 793155
rect 43024 793143 43030 793155
rect 43082 793143 43088 793195
rect 43120 792107 43126 792159
rect 43178 792147 43184 792159
rect 43600 792147 43606 792159
rect 43178 792119 43606 792147
rect 43178 792107 43184 792119
rect 43600 792107 43606 792119
rect 43658 792107 43664 792159
rect 43024 791959 43030 792011
rect 43082 791999 43088 792011
rect 43600 791999 43606 792011
rect 43082 791971 43606 791999
rect 43082 791959 43088 791971
rect 43600 791959 43606 791971
rect 43658 791959 43664 792011
rect 42256 790035 42262 790087
rect 42314 790075 42320 790087
rect 42832 790075 42838 790087
rect 42314 790047 42838 790075
rect 42314 790035 42320 790047
rect 42832 790035 42838 790047
rect 42890 790035 42896 790087
rect 42160 789887 42166 789939
rect 42218 789927 42224 789939
rect 43120 789927 43126 789939
rect 42218 789899 43126 789927
rect 42218 789887 42224 789899
rect 43120 789887 43126 789899
rect 43178 789887 43184 789939
rect 42256 788851 42262 788903
rect 42314 788891 42320 788903
rect 42928 788891 42934 788903
rect 42314 788863 42934 788891
rect 42314 788851 42320 788863
rect 42928 788851 42934 788863
rect 42986 788851 42992 788903
rect 42160 787001 42166 787053
rect 42218 787041 42224 787053
rect 43024 787041 43030 787053
rect 42218 787013 43030 787041
rect 42218 787001 42224 787013
rect 43024 787001 43030 787013
rect 43082 787001 43088 787053
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42448 786449 42454 786461
rect 42218 786421 42454 786449
rect 42218 786409 42224 786421
rect 42448 786409 42454 786421
rect 42506 786409 42512 786461
rect 654448 786261 654454 786313
rect 654506 786301 654512 786313
rect 666832 786301 666838 786313
rect 654506 786273 666838 786301
rect 654506 786261 654512 786273
rect 666832 786261 666838 786273
rect 666890 786261 666896 786313
rect 42064 785595 42070 785647
rect 42122 785635 42128 785647
rect 42736 785635 42742 785647
rect 42122 785607 42742 785635
rect 42122 785595 42128 785607
rect 42736 785595 42742 785607
rect 42794 785595 42800 785647
rect 674512 784929 674518 784981
rect 674570 784969 674576 784981
rect 675376 784969 675382 784981
rect 674570 784941 675382 784969
rect 674570 784929 674576 784941
rect 675376 784929 675382 784941
rect 675434 784929 675440 784981
rect 672208 783449 672214 783501
rect 672266 783489 672272 783501
rect 675376 783489 675382 783501
rect 672266 783461 675382 783489
rect 672266 783449 672272 783461
rect 675376 783449 675382 783461
rect 675434 783449 675440 783501
rect 674992 783005 674998 783057
rect 675050 783045 675056 783057
rect 675376 783045 675382 783057
rect 675050 783017 675382 783045
rect 675050 783005 675056 783017
rect 675376 783005 675382 783017
rect 675434 783005 675440 783057
rect 672496 782265 672502 782317
rect 672554 782305 672560 782317
rect 674608 782305 674614 782317
rect 672554 782277 674614 782305
rect 672554 782265 672560 782277
rect 674608 782265 674614 782277
rect 674666 782305 674672 782317
rect 675376 782305 675382 782317
rect 674666 782277 675382 782305
rect 674666 782265 674672 782277
rect 675376 782265 675382 782277
rect 675434 782265 675440 782317
rect 663856 780489 663862 780541
rect 663914 780529 663920 780541
rect 675088 780529 675094 780541
rect 663914 780501 675094 780529
rect 663914 780489 663920 780501
rect 675088 780489 675094 780501
rect 675146 780489 675152 780541
rect 42736 780415 42742 780467
rect 42794 780455 42800 780467
rect 50608 780455 50614 780467
rect 42794 780427 50614 780455
rect 42794 780415 42800 780427
rect 50608 780415 50614 780427
rect 50666 780415 50672 780467
rect 674416 780415 674422 780467
rect 674474 780455 674480 780467
rect 675472 780455 675478 780467
rect 674474 780427 675478 780455
rect 674474 780415 674480 780427
rect 675472 780415 675478 780427
rect 675530 780415 675536 780467
rect 42448 779897 42454 779949
rect 42506 779937 42512 779949
rect 47536 779937 47542 779949
rect 42506 779909 47542 779937
rect 42506 779897 42512 779909
rect 47536 779897 47542 779909
rect 47594 779897 47600 779949
rect 672688 779749 672694 779801
rect 672746 779789 672752 779801
rect 675376 779789 675382 779801
rect 672746 779761 675382 779789
rect 672746 779749 672752 779761
rect 675376 779749 675382 779761
rect 675434 779749 675440 779801
rect 672016 779305 672022 779357
rect 672074 779345 672080 779357
rect 675472 779345 675478 779357
rect 672074 779317 675478 779345
rect 672074 779305 672080 779317
rect 675472 779305 675478 779317
rect 675530 779305 675536 779357
rect 42736 778861 42742 778913
rect 42794 778901 42800 778913
rect 53392 778901 53398 778913
rect 42794 778873 53398 778901
rect 42794 778861 42800 778873
rect 53392 778861 53398 778873
rect 53450 778861 53456 778913
rect 672112 778565 672118 778617
rect 672170 778605 672176 778617
rect 675376 778605 675382 778617
rect 672170 778577 675382 778605
rect 672170 778565 672176 778577
rect 675376 778565 675382 778577
rect 675434 778565 675440 778617
rect 672400 777603 672406 777655
rect 672458 777643 672464 777655
rect 675472 777643 675478 777655
rect 672458 777615 675478 777643
rect 672458 777603 672464 777615
rect 675472 777603 675478 777615
rect 675530 777603 675536 777655
rect 675088 777011 675094 777063
rect 675146 777051 675152 777063
rect 675376 777051 675382 777063
rect 675146 777023 675382 777051
rect 675146 777011 675152 777023
rect 675376 777011 675382 777023
rect 675434 777011 675440 777063
rect 674800 775457 674806 775509
rect 674858 775497 674864 775509
rect 675376 775497 675382 775509
rect 674858 775469 675382 775497
rect 674858 775457 674864 775469
rect 675376 775457 675382 775469
rect 675434 775457 675440 775509
rect 654448 774717 654454 774769
rect 654506 774757 654512 774769
rect 669808 774757 669814 774769
rect 654506 774729 669814 774757
rect 654506 774717 654512 774729
rect 669808 774717 669814 774729
rect 669866 774717 669872 774769
rect 674224 773607 674230 773659
rect 674282 773647 674288 773659
rect 675376 773647 675382 773659
rect 674282 773619 675382 773647
rect 674282 773607 674288 773619
rect 675376 773607 675382 773619
rect 675434 773607 675440 773659
rect 53392 771831 53398 771883
rect 53450 771871 53456 771883
rect 59536 771871 59542 771883
rect 53450 771843 59542 771871
rect 53450 771831 53456 771843
rect 59536 771831 59542 771843
rect 59594 771831 59600 771883
rect 660976 767761 660982 767813
rect 661034 767801 661040 767813
rect 674704 767801 674710 767813
rect 661034 767773 674710 767801
rect 661034 767761 661040 767773
rect 674704 767761 674710 767773
rect 674762 767761 674768 767813
rect 666736 766873 666742 766925
rect 666794 766913 666800 766925
rect 674704 766913 674710 766925
rect 666794 766885 674710 766913
rect 666794 766873 666800 766885
rect 674704 766873 674710 766885
rect 674762 766873 674768 766925
rect 663952 765837 663958 765889
rect 664010 765877 664016 765889
rect 674320 765877 674326 765889
rect 664010 765849 674326 765877
rect 664010 765837 664016 765849
rect 674320 765837 674326 765849
rect 674378 765837 674384 765889
rect 672304 765245 672310 765297
rect 672362 765285 672368 765297
rect 674704 765285 674710 765297
rect 672362 765257 674710 765285
rect 672362 765245 672368 765257
rect 674704 765245 674710 765257
rect 674762 765245 674768 765297
rect 672592 763987 672598 764039
rect 672650 764027 672656 764039
rect 674704 764027 674710 764039
rect 672650 763999 674710 764027
rect 672650 763987 672656 763999
rect 674704 763987 674710 763999
rect 674762 763987 674768 764039
rect 654448 763247 654454 763299
rect 654506 763287 654512 763299
rect 661072 763287 661078 763299
rect 654506 763259 661078 763287
rect 654506 763247 654512 763259
rect 661072 763247 661078 763259
rect 661130 763247 661136 763299
rect 670960 763173 670966 763225
rect 671018 763213 671024 763225
rect 672880 763213 672886 763225
rect 671018 763185 672886 763213
rect 671018 763173 671024 763185
rect 672880 763173 672886 763185
rect 672938 763213 672944 763225
rect 674704 763213 674710 763225
rect 672938 763185 674710 763213
rect 672938 763173 672944 763185
rect 674704 763173 674710 763185
rect 674762 763173 674768 763225
rect 672880 762507 672886 762559
rect 672938 762547 672944 762559
rect 674704 762547 674710 762559
rect 672938 762519 674710 762547
rect 672938 762507 672944 762519
rect 674704 762507 674710 762519
rect 674762 762507 674768 762559
rect 42928 758067 42934 758119
rect 42986 758107 42992 758119
rect 43216 758107 43222 758119
rect 42986 758079 43222 758107
rect 42986 758067 42992 758079
rect 43216 758067 43222 758079
rect 43274 758067 43280 758119
rect 42928 757919 42934 757971
rect 42986 757959 42992 757971
rect 44944 757959 44950 757971
rect 42986 757931 44950 757959
rect 42986 757919 42992 757931
rect 44944 757919 44950 757931
rect 45002 757919 45008 757971
rect 50416 757475 50422 757527
rect 50474 757515 50480 757527
rect 58192 757515 58198 757527
rect 50474 757487 58198 757515
rect 50474 757475 50480 757487
rect 58192 757475 58198 757487
rect 58250 757475 58256 757527
rect 42448 757253 42454 757305
rect 42506 757293 42512 757305
rect 43504 757293 43510 757305
rect 42506 757265 43510 757293
rect 42506 757253 42512 757265
rect 43504 757253 43510 757265
rect 43562 757253 43568 757305
rect 41968 757105 41974 757157
rect 42026 757145 42032 757157
rect 43696 757145 43702 757157
rect 42026 757117 43702 757145
rect 42026 757105 42032 757117
rect 43696 757105 43702 757117
rect 43754 757105 43760 757157
rect 41872 757031 41878 757083
rect 41930 757071 41936 757083
rect 43600 757071 43606 757083
rect 41930 757043 43606 757071
rect 41930 757031 41936 757043
rect 43600 757031 43606 757043
rect 43658 757031 43664 757083
rect 41776 756957 41782 757009
rect 41834 756957 41840 757009
rect 42064 756957 42070 757009
rect 42122 756997 42128 757009
rect 43312 756997 43318 757009
rect 42122 756969 43318 756997
rect 42122 756957 42128 756969
rect 43312 756957 43318 756969
rect 43370 756957 43376 757009
rect 41794 756787 41822 756957
rect 41776 756735 41782 756787
rect 41834 756735 41840 756787
rect 42160 754071 42166 754123
rect 42218 754111 42224 754123
rect 42928 754111 42934 754123
rect 42218 754083 42934 754111
rect 42218 754071 42224 754083
rect 42928 754071 42934 754083
rect 42986 754071 42992 754123
rect 42928 753923 42934 753975
rect 42986 753963 42992 753975
rect 43216 753963 43222 753975
rect 42986 753935 43222 753963
rect 42986 753923 42992 753935
rect 43216 753923 43222 753935
rect 43274 753923 43280 753975
rect 42064 753035 42070 753087
rect 42122 753075 42128 753087
rect 43120 753075 43126 753087
rect 42122 753047 43126 753075
rect 42122 753035 42128 753047
rect 43120 753035 43126 753047
rect 43178 753035 43184 753087
rect 42928 751891 42934 751903
rect 42850 751863 42934 751891
rect 42850 751829 42878 751863
rect 42928 751851 42934 751863
rect 42986 751851 42992 751903
rect 42064 751777 42070 751829
rect 42122 751817 42128 751829
rect 42736 751817 42742 751829
rect 42122 751789 42742 751817
rect 42122 751777 42128 751789
rect 42736 751777 42742 751789
rect 42794 751777 42800 751829
rect 42832 751777 42838 751829
rect 42890 751777 42896 751829
rect 42928 751703 42934 751755
rect 42986 751743 42992 751755
rect 43696 751743 43702 751755
rect 42986 751715 43702 751743
rect 42986 751703 42992 751715
rect 43696 751703 43702 751715
rect 43754 751703 43760 751755
rect 42064 751111 42070 751163
rect 42122 751151 42128 751163
rect 42832 751151 42838 751163
rect 42122 751123 42838 751151
rect 42122 751111 42128 751123
rect 42832 751111 42838 751123
rect 42890 751111 42896 751163
rect 42832 750963 42838 751015
rect 42890 751003 42896 751015
rect 43600 751003 43606 751015
rect 42890 750975 43606 751003
rect 42890 750963 42896 750975
rect 43600 750963 43606 750975
rect 43658 750963 43664 751015
rect 42160 750371 42166 750423
rect 42218 750411 42224 750423
rect 43120 750411 43126 750423
rect 42218 750383 43126 750411
rect 42218 750371 42224 750383
rect 43120 750371 43126 750383
rect 43178 750371 43184 750423
rect 43120 750223 43126 750275
rect 43178 750263 43184 750275
rect 43504 750263 43510 750275
rect 43178 750235 43510 750263
rect 43178 750223 43184 750235
rect 43504 750223 43510 750235
rect 43562 750223 43568 750275
rect 674032 750223 674038 750275
rect 674090 750263 674096 750275
rect 674416 750263 674422 750275
rect 674090 750235 674422 750263
rect 674090 750223 674096 750235
rect 674416 750223 674422 750235
rect 674474 750223 674480 750275
rect 42064 749927 42070 749979
rect 42122 749967 42128 749979
rect 42928 749967 42934 749979
rect 42122 749939 42934 749967
rect 42122 749927 42128 749939
rect 42928 749927 42934 749939
rect 42986 749927 42992 749979
rect 42256 748891 42262 748943
rect 42314 748931 42320 748943
rect 42832 748931 42838 748943
rect 42314 748903 42838 748931
rect 42314 748891 42320 748903
rect 42832 748891 42838 748903
rect 42890 748891 42896 748943
rect 649552 748817 649558 748869
rect 649610 748857 649616 748869
rect 679792 748857 679798 748869
rect 649610 748829 679798 748857
rect 649610 748817 649616 748829
rect 679792 748817 679798 748829
rect 679850 748817 679856 748869
rect 42160 747411 42166 747463
rect 42218 747451 42224 747463
rect 42448 747451 42454 747463
rect 42218 747423 42454 747451
rect 42218 747411 42224 747423
rect 42448 747411 42454 747423
rect 42506 747411 42512 747463
rect 42064 746079 42070 746131
rect 42122 746119 42128 746131
rect 43120 746119 43126 746131
rect 42122 746091 43126 746119
rect 42122 746079 42128 746091
rect 43120 746079 43126 746091
rect 43178 746079 43184 746131
rect 42160 745635 42166 745687
rect 42218 745675 42224 745687
rect 43024 745675 43030 745687
rect 42218 745647 43030 745675
rect 42218 745635 42224 745647
rect 43024 745635 43030 745647
rect 43082 745635 43088 745687
rect 42160 743785 42166 743837
rect 42218 743825 42224 743837
rect 42736 743825 42742 743837
rect 42218 743797 42742 743825
rect 42218 743785 42224 743797
rect 42736 743785 42742 743797
rect 42794 743785 42800 743837
rect 42064 743045 42070 743097
rect 42122 743085 42128 743097
rect 42832 743085 42838 743097
rect 42122 743057 42838 743085
rect 42122 743045 42128 743057
rect 42832 743045 42838 743057
rect 42890 743045 42896 743097
rect 47536 743045 47542 743097
rect 47594 743085 47600 743097
rect 58576 743085 58582 743097
rect 47594 743057 58582 743085
rect 47594 743045 47600 743057
rect 58576 743045 58582 743057
rect 58634 743045 58640 743097
rect 42160 742379 42166 742431
rect 42218 742419 42224 742431
rect 42928 742419 42934 742431
rect 42218 742391 42934 742419
rect 42218 742379 42224 742391
rect 42928 742379 42934 742391
rect 42986 742379 42992 742431
rect 674896 737865 674902 737917
rect 674954 737905 674960 737917
rect 675376 737905 675382 737917
rect 674954 737877 675382 737905
rect 674954 737865 674960 737877
rect 675376 737865 675382 737877
rect 675434 737865 675440 737917
rect 672496 737643 672502 737695
rect 672554 737683 672560 737695
rect 675472 737683 675478 737695
rect 672554 737655 675478 737683
rect 672554 737643 672560 737655
rect 675472 737643 675478 737655
rect 675530 737643 675536 737695
rect 660976 737347 660982 737399
rect 661034 737387 661040 737399
rect 675088 737387 675094 737399
rect 661034 737359 675094 737387
rect 661034 737347 661040 737359
rect 675088 737347 675094 737359
rect 675146 737347 675152 737399
rect 654448 737273 654454 737325
rect 654506 737313 654512 737325
rect 663952 737313 663958 737325
rect 654506 737285 663958 737313
rect 654506 737273 654512 737285
rect 663952 737273 663958 737285
rect 664010 737273 664016 737325
rect 42640 737199 42646 737251
rect 42698 737239 42704 737251
rect 53392 737239 53398 737251
rect 42698 737211 53398 737239
rect 42698 737199 42704 737211
rect 53392 737199 53398 737211
rect 53450 737199 53456 737251
rect 42352 736681 42358 736733
rect 42410 736721 42416 736733
rect 50416 736721 50422 736733
rect 42410 736693 50422 736721
rect 42410 736681 42416 736693
rect 50416 736681 50422 736693
rect 50474 736681 50480 736733
rect 674128 735645 674134 735697
rect 674186 735685 674192 735697
rect 675472 735685 675478 735697
rect 674186 735657 675478 735685
rect 674186 735645 674192 735657
rect 675472 735645 675478 735657
rect 675530 735645 675536 735697
rect 42352 735423 42358 735475
rect 42410 735463 42416 735475
rect 58960 735463 58966 735475
rect 42410 735435 58966 735463
rect 42410 735423 42416 735435
rect 58960 735423 58966 735435
rect 59018 735423 59024 735475
rect 675184 734905 675190 734957
rect 675242 734945 675248 734957
rect 675376 734945 675382 734957
rect 675242 734917 675382 734945
rect 675242 734905 675248 734917
rect 675376 734905 675382 734917
rect 675434 734905 675440 734957
rect 672304 733573 672310 733625
rect 672362 733613 672368 733625
rect 675472 733613 675478 733625
rect 672362 733585 675478 733613
rect 672362 733573 672368 733585
rect 675472 733573 675478 733585
rect 675530 733573 675536 733625
rect 675184 732315 675190 732367
rect 675242 732355 675248 732367
rect 675472 732355 675478 732367
rect 675242 732327 675478 732355
rect 675242 732315 675248 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 675088 732019 675094 732071
rect 675146 732059 675152 732071
rect 675376 732059 675382 732071
rect 675146 732031 675382 732059
rect 675146 732019 675152 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 674704 730465 674710 730517
rect 674762 730505 674768 730517
rect 675472 730505 675478 730517
rect 674762 730477 675478 730505
rect 674762 730465 674768 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 50416 728615 50422 728667
rect 50474 728655 50480 728667
rect 59536 728655 59542 728667
rect 50474 728627 59542 728655
rect 50474 728615 50480 728627
rect 59536 728615 59542 728627
rect 59594 728615 59600 728667
rect 674608 728615 674614 728667
rect 674666 728655 674672 728667
rect 675472 728655 675478 728667
rect 674666 728627 675478 728655
rect 674666 728615 674672 728627
rect 675472 728615 675478 728627
rect 675530 728615 675536 728667
rect 674800 726321 674806 726373
rect 674858 726361 674864 726373
rect 675088 726361 675094 726373
rect 674858 726333 675094 726361
rect 674858 726321 674864 726333
rect 675088 726321 675094 726333
rect 675146 726321 675152 726373
rect 663760 722473 663766 722525
rect 663818 722513 663824 722525
rect 674320 722513 674326 722525
rect 663818 722485 674326 722513
rect 663818 722473 663824 722485
rect 674320 722473 674326 722485
rect 674378 722473 674384 722525
rect 660880 721881 660886 721933
rect 660938 721921 660944 721933
rect 674800 721921 674806 721933
rect 660938 721893 674806 721921
rect 660938 721881 660944 721893
rect 674800 721881 674806 721893
rect 674858 721881 674864 721933
rect 661168 720845 661174 720897
rect 661226 720885 661232 720897
rect 674320 720885 674326 720897
rect 661226 720857 674326 720885
rect 661226 720845 661232 720857
rect 674320 720845 674326 720857
rect 674378 720845 674384 720897
rect 672592 720253 672598 720305
rect 672650 720293 672656 720305
rect 674800 720293 674806 720305
rect 672650 720265 674806 720293
rect 672650 720253 672656 720265
rect 674800 720253 674806 720265
rect 674858 720253 674864 720305
rect 674032 720031 674038 720083
rect 674090 720071 674096 720083
rect 674320 720071 674326 720083
rect 674090 720043 674326 720071
rect 674090 720031 674096 720043
rect 674320 720031 674326 720043
rect 674378 720031 674384 720083
rect 671920 718995 671926 719047
rect 671978 719035 671984 719047
rect 674800 719035 674806 719047
rect 671978 719007 674806 719035
rect 671978 718995 671984 719007
rect 674800 718995 674806 719007
rect 674858 718995 674864 719047
rect 42256 718699 42262 718751
rect 42314 718739 42320 718751
rect 44944 718739 44950 718751
rect 42314 718711 44950 718739
rect 42314 718699 42320 718711
rect 44944 718699 44950 718711
rect 45002 718699 45008 718751
rect 672880 717811 672886 717863
rect 672938 717851 672944 717863
rect 674512 717851 674518 717863
rect 672938 717823 674518 717851
rect 672938 717811 672944 717823
rect 674512 717811 674518 717823
rect 674570 717811 674576 717863
rect 672592 717145 672598 717197
rect 672650 717185 672656 717197
rect 672880 717185 672886 717197
rect 672650 717157 672886 717185
rect 672650 717145 672656 717157
rect 672880 717145 672886 717157
rect 672938 717145 672944 717197
rect 43120 717071 43126 717123
rect 43178 717111 43184 717123
rect 45040 717111 45046 717123
rect 43178 717083 45046 717111
rect 43178 717071 43184 717083
rect 45040 717071 45046 717083
rect 45098 717071 45104 717123
rect 670960 717071 670966 717123
rect 671018 717111 671024 717123
rect 679696 717111 679702 717123
rect 671018 717083 679702 717111
rect 671018 717071 671024 717083
rect 679696 717071 679702 717083
rect 679754 717071 679760 717123
rect 40240 714999 40246 715051
rect 40298 715039 40304 715051
rect 41872 715039 41878 715051
rect 40298 715011 41878 715039
rect 40298 714999 40304 715011
rect 41872 714999 41878 715011
rect 41930 714999 41936 715051
rect 53392 714259 53398 714311
rect 53450 714299 53456 714311
rect 59536 714299 59542 714311
rect 53450 714271 59542 714299
rect 53450 714259 53456 714271
rect 59536 714259 59542 714271
rect 59594 714259 59600 714311
rect 654448 714259 654454 714311
rect 654506 714299 654512 714311
rect 664144 714299 664150 714311
rect 654506 714271 664150 714299
rect 654506 714259 654512 714271
rect 664144 714259 664150 714271
rect 664202 714259 664208 714311
rect 41584 714111 41590 714163
rect 41642 714151 41648 714163
rect 43504 714151 43510 714163
rect 41642 714123 43510 714151
rect 41642 714111 41648 714123
rect 43504 714111 43510 714123
rect 43562 714111 43568 714163
rect 41488 714037 41494 714089
rect 41546 714037 41552 714089
rect 41680 714037 41686 714089
rect 41738 714077 41744 714089
rect 43600 714077 43606 714089
rect 41738 714049 43606 714077
rect 41738 714037 41744 714049
rect 43600 714037 43606 714049
rect 43658 714037 43664 714089
rect 41506 713559 41534 714037
rect 41968 713815 41974 713867
rect 42026 713855 42032 713867
rect 43312 713855 43318 713867
rect 42026 713827 43318 713855
rect 42026 713815 42032 713827
rect 43312 713815 43318 713827
rect 43370 713815 43376 713867
rect 41776 713559 41782 713571
rect 41506 713531 41782 713559
rect 41776 713519 41782 713531
rect 41834 713519 41840 713571
rect 43312 711561 43318 711573
rect 42946 711533 43318 711561
rect 42946 711499 42974 711533
rect 43312 711521 43318 711533
rect 43370 711521 43376 711573
rect 42928 711447 42934 711499
rect 42986 711447 42992 711499
rect 43120 711447 43126 711499
rect 43178 711487 43184 711499
rect 43178 711459 43454 711487
rect 43178 711447 43184 711459
rect 43426 711425 43454 711459
rect 43408 711373 43414 711425
rect 43466 711373 43472 711425
rect 42928 711299 42934 711351
rect 42986 711339 42992 711351
rect 42986 711311 43070 711339
rect 42986 711299 42992 711311
rect 43042 711265 43070 711311
rect 43696 711265 43702 711277
rect 43042 711237 43702 711265
rect 43696 711225 43702 711237
rect 43754 711225 43760 711277
rect 42160 710855 42166 710907
rect 42218 710895 42224 710907
rect 43408 710895 43414 710907
rect 42218 710867 43414 710895
rect 42218 710855 42224 710867
rect 43408 710855 43414 710867
rect 43466 710855 43472 710907
rect 672208 710485 672214 710537
rect 672266 710525 672272 710537
rect 674416 710525 674422 710537
rect 672266 710497 674422 710525
rect 672266 710485 672272 710497
rect 674416 710485 674422 710497
rect 674474 710485 674480 710537
rect 42160 709893 42166 709945
rect 42218 709933 42224 709945
rect 42352 709933 42358 709945
rect 42218 709905 42358 709933
rect 42218 709893 42224 709905
rect 42352 709893 42358 709905
rect 42410 709893 42416 709945
rect 672400 709893 672406 709945
rect 672458 709933 672464 709945
rect 674800 709933 674806 709945
rect 672458 709905 674806 709933
rect 672458 709893 672464 709905
rect 674800 709893 674806 709905
rect 674858 709893 674864 709945
rect 672016 709005 672022 709057
rect 672074 709045 672080 709057
rect 674416 709045 674422 709057
rect 672074 709017 674422 709045
rect 672074 709005 672080 709017
rect 674416 709005 674422 709017
rect 674474 709005 674480 709057
rect 42160 707895 42166 707947
rect 42218 707935 42224 707947
rect 43696 707935 43702 707947
rect 42218 707907 43702 707935
rect 42218 707895 42224 707907
rect 43696 707895 43702 707907
rect 43754 707895 43760 707947
rect 672688 707377 672694 707429
rect 672746 707417 672752 707429
rect 674416 707417 674422 707429
rect 672746 707389 674422 707417
rect 672746 707377 672752 707389
rect 674416 707377 674422 707389
rect 674474 707377 674480 707429
rect 42928 707229 42934 707281
rect 42986 707269 42992 707281
rect 43600 707269 43606 707281
rect 42986 707241 43606 707269
rect 42986 707229 42992 707241
rect 43600 707229 43606 707241
rect 43658 707229 43664 707281
rect 672112 706785 672118 706837
rect 672170 706825 672176 706837
rect 674800 706825 674806 706837
rect 672170 706797 674806 706825
rect 672170 706785 672176 706797
rect 674800 706785 674806 706797
rect 674858 706785 674864 706837
rect 42544 706415 42550 706467
rect 42602 706455 42608 706467
rect 43504 706455 43510 706467
rect 42602 706427 43510 706455
rect 42602 706415 42608 706427
rect 43504 706415 43510 706427
rect 43562 706415 43568 706467
rect 42256 705601 42262 705653
rect 42314 705641 42320 705653
rect 43120 705641 43126 705653
rect 42314 705613 43126 705641
rect 42314 705601 42320 705613
rect 43120 705601 43126 705613
rect 43178 705601 43184 705653
rect 42064 703677 42070 703729
rect 42122 703717 42128 703729
rect 42832 703717 42838 703729
rect 42122 703689 42838 703717
rect 42122 703677 42128 703689
rect 42832 703677 42838 703689
rect 42890 703677 42896 703729
rect 42160 702863 42166 702915
rect 42218 702903 42224 702915
rect 42928 702903 42934 702915
rect 42218 702875 42934 702903
rect 42218 702863 42224 702875
rect 42928 702863 42934 702875
rect 42986 702863 42992 702915
rect 649648 702715 649654 702767
rect 649706 702755 649712 702767
rect 679792 702755 679798 702767
rect 649706 702727 679798 702755
rect 649706 702715 649712 702727
rect 679792 702715 679798 702727
rect 679850 702715 679856 702767
rect 672496 702641 672502 702693
rect 672554 702681 672560 702693
rect 674800 702681 674806 702693
rect 672554 702653 674806 702681
rect 672554 702641 672560 702653
rect 674800 702641 674806 702653
rect 674858 702641 674864 702693
rect 42160 702271 42166 702323
rect 42218 702311 42224 702323
rect 42544 702311 42550 702323
rect 42218 702283 42550 702311
rect 42218 702271 42224 702283
rect 42544 702271 42550 702283
rect 42602 702271 42608 702323
rect 42064 700569 42070 700621
rect 42122 700609 42128 700621
rect 43024 700609 43030 700621
rect 42122 700581 43030 700609
rect 42122 700569 42128 700581
rect 43024 700569 43030 700581
rect 43082 700569 43088 700621
rect 42160 700051 42166 700103
rect 42218 700091 42224 700103
rect 42832 700091 42838 700103
rect 42218 700063 42838 700091
rect 42218 700051 42224 700063
rect 42832 700051 42838 700063
rect 42890 700051 42896 700103
rect 670960 699903 670966 699955
rect 671018 699943 671024 699955
rect 679696 699943 679702 699955
rect 671018 699915 679702 699943
rect 671018 699903 671024 699915
rect 679696 699903 679702 699915
rect 679754 699903 679760 699955
rect 42352 699829 42358 699881
rect 42410 699869 42416 699881
rect 59536 699869 59542 699881
rect 42410 699841 59542 699869
rect 42410 699829 42416 699841
rect 59536 699829 59542 699841
rect 59594 699829 59600 699881
rect 42640 693983 42646 694035
rect 42698 694023 42704 694035
rect 53392 694023 53398 694035
rect 42698 693995 53398 694023
rect 42698 693983 42704 693995
rect 53392 693983 53398 693995
rect 53450 693983 53456 694035
rect 672208 692873 672214 692925
rect 672266 692913 672272 692925
rect 675376 692913 675382 692925
rect 672266 692885 675382 692913
rect 672266 692873 672272 692885
rect 675376 692873 675382 692885
rect 675434 692873 675440 692925
rect 42640 692429 42646 692481
rect 42698 692469 42704 692481
rect 50416 692469 50422 692481
rect 42698 692441 50422 692469
rect 42698 692429 42704 692441
rect 50416 692429 50422 692441
rect 50474 692429 50480 692481
rect 672400 692429 672406 692481
rect 672458 692469 672464 692481
rect 674800 692469 674806 692481
rect 672458 692441 674806 692469
rect 672458 692429 672464 692441
rect 674800 692429 674806 692441
rect 674858 692469 674864 692481
rect 675472 692469 675478 692481
rect 674858 692441 675478 692469
rect 674858 692429 674864 692441
rect 675472 692429 675478 692441
rect 675530 692429 675536 692481
rect 654832 691245 654838 691297
rect 654890 691285 654896 691297
rect 666928 691285 666934 691297
rect 654890 691257 666934 691285
rect 654890 691245 654896 691257
rect 666928 691245 666934 691257
rect 666986 691245 666992 691297
rect 674320 690653 674326 690705
rect 674378 690693 674384 690705
rect 675472 690693 675478 690705
rect 674378 690665 675478 690693
rect 674378 690653 674384 690665
rect 675472 690653 675478 690665
rect 675530 690653 675536 690705
rect 675088 689765 675094 689817
rect 675146 689805 675152 689817
rect 675376 689805 675382 689817
rect 675146 689777 675382 689805
rect 675146 689765 675152 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 672112 688581 672118 688633
rect 672170 688621 672176 688633
rect 675472 688621 675478 688633
rect 672170 688593 675478 688621
rect 672170 688581 672176 688593
rect 675472 688581 675478 688593
rect 675530 688581 675536 688633
rect 674224 687323 674230 687375
rect 674282 687363 674288 687375
rect 675472 687363 675478 687375
rect 674282 687335 675478 687363
rect 674282 687323 674288 687335
rect 675472 687323 675478 687335
rect 675530 687323 675536 687375
rect 669616 686213 669622 686265
rect 669674 686253 669680 686265
rect 675376 686253 675382 686265
rect 669674 686225 675382 686253
rect 669674 686213 669680 686225
rect 675376 686213 675382 686225
rect 675434 686213 675440 686265
rect 50416 685473 50422 685525
rect 50474 685513 50480 685525
rect 58672 685513 58678 685525
rect 50474 685485 58678 685513
rect 50474 685473 50480 685485
rect 58672 685473 58678 685485
rect 58730 685473 58736 685525
rect 674512 685473 674518 685525
rect 674570 685513 674576 685525
rect 675472 685513 675478 685525
rect 674570 685485 675478 685513
rect 674570 685473 674576 685485
rect 675472 685473 675478 685485
rect 675530 685473 675536 685525
rect 674896 683623 674902 683675
rect 674954 683663 674960 683675
rect 675472 683663 675478 683675
rect 674954 683635 675478 683663
rect 674954 683623 674960 683635
rect 675472 683623 675478 683635
rect 675530 683623 675536 683675
rect 667024 677481 667030 677533
rect 667082 677521 667088 677533
rect 674800 677521 674806 677533
rect 667082 677493 674806 677521
rect 667082 677481 667088 677493
rect 674800 677481 674806 677493
rect 674858 677481 674864 677533
rect 649744 676815 649750 676867
rect 649802 676855 649808 676867
rect 653680 676855 653686 676867
rect 649802 676827 653686 676855
rect 649802 676815 649808 676827
rect 653680 676815 653686 676827
rect 653738 676815 653744 676867
rect 669712 676445 669718 676497
rect 669770 676485 669776 676497
rect 674416 676485 674422 676497
rect 669770 676457 674422 676485
rect 669770 676445 669776 676457
rect 674416 676445 674422 676457
rect 674474 676445 674480 676497
rect 664048 675853 664054 675905
rect 664106 675893 664112 675905
rect 674800 675893 674806 675905
rect 664106 675865 674806 675893
rect 664106 675853 664112 675865
rect 674800 675853 674806 675865
rect 674858 675853 674864 675905
rect 42352 675631 42358 675683
rect 42410 675671 42416 675683
rect 45040 675671 45046 675683
rect 42410 675643 45046 675671
rect 42410 675631 42416 675643
rect 45040 675631 45046 675643
rect 45098 675631 45104 675683
rect 671920 674817 671926 674869
rect 671978 674857 671984 674869
rect 674416 674857 674422 674869
rect 671978 674829 674422 674857
rect 671978 674817 671984 674829
rect 674416 674817 674422 674829
rect 674474 674817 674480 674869
rect 41584 674521 41590 674573
rect 41642 674561 41648 674573
rect 43120 674561 43126 674573
rect 41642 674533 43126 674561
rect 41642 674521 41648 674533
rect 43120 674521 43126 674533
rect 43178 674521 43184 674573
rect 672688 674003 672694 674055
rect 672746 674043 672752 674055
rect 674416 674043 674422 674055
rect 672746 674015 674422 674043
rect 672746 674003 672752 674015
rect 674416 674003 674422 674015
rect 674474 674003 674480 674055
rect 670960 673115 670966 673167
rect 671018 673155 671024 673167
rect 672496 673155 672502 673167
rect 671018 673127 672502 673155
rect 671018 673115 671024 673127
rect 672496 673115 672502 673127
rect 672554 673155 672560 673167
rect 674800 673155 674806 673167
rect 672554 673127 674806 673155
rect 672554 673115 672560 673127
rect 674800 673115 674806 673127
rect 674858 673115 674864 673167
rect 40240 672153 40246 672205
rect 40298 672193 40304 672205
rect 41008 672193 41014 672205
rect 40298 672165 41014 672193
rect 40298 672153 40304 672165
rect 41008 672153 41014 672165
rect 41066 672153 41072 672205
rect 41680 672005 41686 672057
rect 41738 672045 41744 672057
rect 42640 672045 42646 672057
rect 41738 672017 42646 672045
rect 41738 672005 41744 672017
rect 42640 672005 42646 672017
rect 42698 672005 42704 672057
rect 42256 671931 42262 671983
rect 42314 671971 42320 671983
rect 42448 671971 42454 671983
rect 42314 671943 42454 671971
rect 42314 671931 42320 671943
rect 42448 671931 42454 671943
rect 42506 671931 42512 671983
rect 43312 671339 43318 671391
rect 43370 671379 43376 671391
rect 45136 671379 45142 671391
rect 43370 671351 45142 671379
rect 43370 671339 43376 671351
rect 45136 671339 45142 671351
rect 45194 671339 45200 671391
rect 53392 671043 53398 671095
rect 53450 671083 53456 671095
rect 58384 671083 58390 671095
rect 53450 671055 58390 671083
rect 53450 671043 53456 671055
rect 58384 671043 58390 671055
rect 58442 671043 58448 671095
rect 672592 670969 672598 671021
rect 672650 671009 672656 671021
rect 675088 671009 675094 671021
rect 672650 670981 675094 671009
rect 672650 670969 672656 670981
rect 675088 670969 675094 670981
rect 675146 670969 675152 671021
rect 43120 670821 43126 670873
rect 43178 670861 43184 670873
rect 43504 670861 43510 670873
rect 43178 670833 43510 670861
rect 43178 670821 43184 670833
rect 43504 670821 43510 670833
rect 43562 670821 43568 670873
rect 41872 670747 41878 670799
rect 41930 670787 41936 670799
rect 43216 670787 43222 670799
rect 41930 670759 43222 670787
rect 41930 670747 41936 670759
rect 43216 670747 43222 670759
rect 43274 670747 43280 670799
rect 41776 670599 41782 670651
rect 41834 670599 41840 670651
rect 41968 670599 41974 670651
rect 42026 670639 42032 670651
rect 42928 670639 42934 670651
rect 42026 670611 42934 670639
rect 42026 670599 42032 670611
rect 42928 670599 42934 670611
rect 42986 670599 42992 670651
rect 41794 670355 41822 670599
rect 41776 670303 41782 670355
rect 41834 670303 41840 670355
rect 674416 669563 674422 669615
rect 674474 669603 674480 669615
rect 674896 669603 674902 669615
rect 674474 669575 674902 669603
rect 674474 669563 674480 669575
rect 674896 669563 674902 669575
rect 674954 669563 674960 669615
rect 42448 669193 42454 669245
rect 42506 669233 42512 669245
rect 42506 669205 42974 669233
rect 42506 669193 42512 669205
rect 42832 668897 42838 668949
rect 42890 668937 42896 668949
rect 42946 668937 42974 669205
rect 42890 668909 42974 668937
rect 42890 668897 42896 668909
rect 654448 668157 654454 668209
rect 654506 668197 654512 668209
rect 661264 668197 661270 668209
rect 654506 668169 661270 668197
rect 654506 668157 654512 668169
rect 661264 668157 661270 668169
rect 661322 668157 661328 668209
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 43312 667901 43318 667913
rect 42218 667873 43318 667901
rect 42218 667861 42224 667873
rect 43312 667861 43318 667873
rect 43370 667861 43376 667913
rect 42160 666677 42166 666729
rect 42218 666717 42224 666729
rect 42928 666717 42934 666729
rect 42218 666689 42934 666717
rect 42218 666677 42224 666689
rect 42928 666677 42934 666689
rect 42986 666677 42992 666729
rect 42160 664827 42166 664879
rect 42218 664867 42224 664879
rect 42832 664867 42838 664879
rect 42218 664839 42838 664867
rect 42218 664827 42224 664839
rect 42832 664827 42838 664839
rect 42890 664827 42896 664879
rect 42832 664679 42838 664731
rect 42890 664719 42896 664731
rect 43600 664719 43606 664731
rect 42890 664691 43606 664719
rect 42890 664679 42896 664691
rect 43600 664679 43606 664691
rect 43658 664679 43664 664731
rect 42160 664161 42166 664213
rect 42218 664201 42224 664213
rect 43120 664201 43126 664213
rect 42218 664173 43126 664201
rect 42218 664161 42224 664173
rect 43120 664161 43126 664173
rect 43178 664161 43184 664213
rect 43120 664013 43126 664065
rect 43178 664053 43184 664065
rect 43504 664053 43510 664065
rect 43178 664025 43510 664053
rect 43178 664013 43184 664025
rect 43504 664013 43510 664025
rect 43562 664013 43568 664065
rect 42544 663495 42550 663547
rect 42602 663495 42608 663547
rect 42160 663347 42166 663399
rect 42218 663387 42224 663399
rect 42562 663387 42590 663495
rect 42218 663359 42590 663387
rect 42218 663347 42224 663359
rect 42256 662385 42262 662437
rect 42314 662425 42320 662437
rect 43024 662425 43030 662437
rect 42314 662397 43030 662425
rect 42314 662385 42320 662397
rect 43024 662385 43030 662397
rect 43082 662385 43088 662437
rect 672304 661645 672310 661697
rect 672362 661685 672368 661697
rect 674704 661685 674710 661697
rect 672362 661657 674710 661685
rect 672362 661645 672368 661657
rect 674704 661645 674710 661657
rect 674762 661645 674768 661697
rect 42160 661053 42166 661105
rect 42218 661093 42224 661105
rect 42832 661093 42838 661105
rect 42218 661065 42838 661093
rect 42218 661053 42224 661065
rect 42832 661053 42838 661065
rect 42890 661053 42896 661105
rect 42160 659647 42166 659699
rect 42218 659687 42224 659699
rect 42928 659687 42934 659699
rect 42218 659659 42934 659687
rect 42218 659647 42224 659659
rect 42928 659647 42934 659659
rect 42986 659647 42992 659699
rect 42064 659055 42070 659107
rect 42122 659095 42128 659107
rect 42544 659095 42550 659107
rect 42122 659067 42550 659095
rect 42122 659055 42128 659067
rect 42544 659055 42550 659067
rect 42602 659055 42608 659107
rect 42160 656835 42166 656887
rect 42218 656875 42224 656887
rect 42832 656875 42838 656887
rect 42218 656847 42838 656875
rect 42218 656835 42224 656847
rect 42832 656835 42838 656847
rect 42890 656835 42896 656887
rect 42064 656761 42070 656813
rect 42122 656801 42128 656813
rect 43120 656801 43126 656813
rect 42122 656773 43126 656801
rect 42122 656761 42128 656773
rect 43120 656761 43126 656773
rect 43178 656761 43184 656813
rect 42832 656687 42838 656739
rect 42890 656727 42896 656739
rect 59536 656727 59542 656739
rect 42890 656699 59542 656727
rect 42890 656687 42896 656699
rect 59536 656687 59542 656699
rect 59594 656687 59600 656739
rect 649744 656687 649750 656739
rect 649802 656727 649808 656739
rect 679792 656727 679798 656739
rect 649802 656699 679798 656727
rect 649802 656687 649808 656699
rect 679792 656687 679798 656699
rect 679850 656687 679856 656739
rect 672400 650915 672406 650967
rect 672458 650955 672464 650967
rect 674800 650955 674806 650967
rect 672458 650927 674806 650955
rect 672458 650915 672464 650927
rect 674800 650915 674806 650927
rect 674858 650915 674864 650967
rect 674608 650841 674614 650893
rect 674666 650881 674672 650893
rect 674992 650881 674998 650893
rect 674666 650853 674998 650881
rect 674666 650841 674672 650853
rect 674992 650841 674998 650853
rect 675050 650841 675056 650893
rect 42448 649731 42454 649783
rect 42506 649771 42512 649783
rect 51856 649771 51862 649783
rect 42506 649743 51862 649771
rect 42506 649731 42512 649743
rect 51856 649731 51862 649743
rect 51914 649731 51920 649783
rect 42448 649509 42454 649561
rect 42506 649549 42512 649561
rect 53392 649549 53398 649561
rect 42506 649521 53398 649549
rect 42506 649509 42512 649521
rect 53392 649509 53398 649521
rect 53450 649509 53456 649561
rect 671920 648251 671926 648303
rect 671978 648291 671984 648303
rect 675280 648291 675286 648303
rect 671978 648263 675286 648291
rect 671978 648251 671984 648263
rect 675280 648251 675286 648263
rect 675338 648251 675344 648303
rect 672880 648029 672886 648081
rect 672938 648069 672944 648081
rect 675184 648069 675190 648081
rect 672938 648041 675190 648069
rect 672938 648029 672944 648041
rect 675184 648029 675190 648041
rect 675242 648029 675248 648081
rect 674800 647585 674806 647637
rect 674858 647625 674864 647637
rect 675088 647625 675094 647637
rect 674858 647597 675094 647625
rect 674858 647585 674864 647597
rect 675088 647585 675094 647597
rect 675146 647585 675152 647637
rect 674608 646401 674614 646453
rect 674666 646441 674672 646453
rect 675376 646441 675382 646453
rect 674666 646413 675382 646441
rect 674666 646401 674672 646413
rect 675376 646401 675382 646413
rect 675434 646401 675440 646453
rect 666736 645217 666742 645269
rect 666794 645257 666800 645269
rect 675184 645257 675190 645269
rect 666794 645229 675190 645257
rect 666794 645217 666800 645229
rect 675184 645217 675190 645229
rect 675242 645217 675248 645269
rect 654448 645143 654454 645195
rect 654506 645183 654512 645195
rect 669712 645183 669718 645195
rect 654506 645155 669718 645183
rect 654506 645143 654512 645155
rect 669712 645143 669718 645155
rect 669770 645143 669776 645195
rect 674800 645069 674806 645121
rect 674858 645109 674864 645121
rect 675088 645109 675094 645121
rect 674858 645081 675094 645109
rect 674858 645069 674864 645081
rect 675088 645069 675094 645081
rect 675146 645069 675152 645121
rect 671632 644551 671638 644603
rect 671690 644591 671696 644603
rect 675472 644591 675478 644603
rect 671690 644563 675478 644591
rect 671690 644551 671696 644563
rect 675472 644551 675478 644563
rect 675530 644551 675536 644603
rect 51856 644477 51862 644529
rect 51914 644517 51920 644529
rect 59536 644517 59542 644529
rect 51914 644489 59542 644517
rect 51914 644477 51920 644489
rect 59536 644477 59542 644489
rect 59594 644477 59600 644529
rect 672304 644033 672310 644085
rect 672362 644073 672368 644085
rect 675472 644073 675478 644085
rect 672362 644045 675478 644073
rect 672362 644033 672368 644045
rect 675472 644033 675478 644045
rect 675530 644033 675536 644085
rect 672592 643367 672598 643419
rect 672650 643407 672656 643419
rect 675376 643407 675382 643419
rect 672650 643379 675382 643407
rect 672650 643367 672656 643379
rect 675376 643367 675382 643379
rect 675434 643367 675440 643419
rect 671440 642257 671446 642309
rect 671498 642297 671504 642309
rect 675472 642297 675478 642309
rect 671498 642269 675478 642297
rect 671498 642257 671504 642269
rect 675472 642257 675478 642269
rect 675530 642257 675536 642309
rect 675184 641813 675190 641865
rect 675242 641853 675248 641865
rect 675376 641853 675382 641865
rect 675242 641825 675382 641853
rect 675242 641813 675248 641825
rect 675376 641813 675382 641825
rect 675434 641813 675440 641865
rect 670864 633599 670870 633651
rect 670922 633639 670928 633651
rect 674992 633639 674998 633651
rect 670922 633611 674998 633639
rect 670922 633599 670928 633611
rect 674992 633599 674998 633611
rect 675050 633599 675056 633651
rect 669808 632489 669814 632541
rect 669866 632529 669872 632541
rect 674704 632529 674710 632541
rect 669866 632501 674710 632529
rect 669866 632489 669872 632501
rect 674704 632489 674710 632501
rect 674762 632489 674768 632541
rect 42256 632415 42262 632467
rect 42314 632455 42320 632467
rect 45136 632455 45142 632467
rect 42314 632427 45142 632455
rect 42314 632415 42320 632427
rect 45136 632415 45142 632427
rect 45194 632415 45200 632467
rect 666832 631749 666838 631801
rect 666890 631789 666896 631801
rect 674704 631789 674710 631801
rect 666890 631761 674710 631789
rect 666890 631749 666896 631761
rect 674704 631749 674710 631761
rect 674762 631749 674768 631801
rect 670960 630713 670966 630765
rect 671018 630753 671024 630765
rect 672496 630753 672502 630765
rect 671018 630725 672502 630753
rect 671018 630713 671024 630725
rect 672496 630713 672502 630725
rect 672554 630713 672560 630765
rect 661072 630565 661078 630617
rect 661130 630605 661136 630617
rect 674128 630605 674134 630617
rect 661130 630577 674134 630605
rect 661130 630565 661136 630577
rect 674128 630565 674134 630577
rect 674186 630565 674192 630617
rect 672688 630491 672694 630543
rect 672746 630531 672752 630543
rect 673840 630531 673846 630543
rect 672746 630503 673846 630531
rect 672746 630491 672752 630503
rect 673840 630491 673846 630503
rect 673898 630491 673904 630543
rect 42928 628419 42934 628471
rect 42986 628459 42992 628471
rect 43600 628459 43606 628471
rect 42986 628431 43606 628459
rect 42986 628419 42992 628431
rect 43600 628419 43606 628431
rect 43658 628419 43664 628471
rect 42448 627901 42454 627953
rect 42506 627941 42512 627953
rect 47728 627941 47734 627953
rect 42506 627913 47734 627941
rect 42506 627901 42512 627913
rect 47728 627901 47734 627913
rect 47786 627901 47792 627953
rect 40048 627827 40054 627879
rect 40106 627867 40112 627879
rect 41200 627867 41206 627879
rect 40106 627839 41206 627867
rect 40106 627827 40112 627839
rect 41200 627827 41206 627839
rect 41258 627827 41264 627879
rect 43120 627827 43126 627879
rect 43178 627867 43184 627879
rect 43408 627867 43414 627879
rect 43178 627839 43414 627867
rect 43178 627827 43184 627839
rect 43408 627827 43414 627839
rect 43466 627827 43472 627879
rect 47632 627827 47638 627879
rect 47690 627867 47696 627879
rect 58384 627867 58390 627879
rect 47690 627839 58390 627867
rect 47690 627827 47696 627839
rect 58384 627827 58390 627839
rect 58442 627827 58448 627879
rect 671728 627827 671734 627879
rect 671786 627867 671792 627879
rect 673840 627867 673846 627879
rect 671786 627839 673846 627867
rect 671786 627827 671792 627839
rect 673840 627827 673846 627839
rect 673898 627827 673904 627879
rect 41680 627753 41686 627805
rect 41738 627793 41744 627805
rect 43504 627793 43510 627805
rect 41738 627765 43510 627793
rect 41738 627753 41744 627765
rect 43504 627753 43510 627765
rect 43562 627753 43568 627805
rect 41488 627679 41494 627731
rect 41546 627719 41552 627731
rect 43120 627719 43126 627731
rect 41546 627691 43126 627719
rect 41546 627679 41552 627691
rect 43120 627679 43126 627691
rect 43178 627679 43184 627731
rect 41776 627383 41782 627435
rect 41834 627383 41840 627435
rect 42064 627383 42070 627435
rect 42122 627423 42128 627435
rect 43024 627423 43030 627435
rect 42122 627395 43030 627423
rect 42122 627383 42128 627395
rect 43024 627383 43030 627395
rect 43082 627383 43088 627435
rect 41794 627213 41822 627383
rect 41776 627161 41782 627213
rect 41834 627161 41840 627213
rect 42928 625163 42934 625215
rect 42986 625203 42992 625215
rect 43408 625203 43414 625215
rect 42986 625175 43414 625203
rect 42986 625163 42992 625175
rect 43408 625163 43414 625175
rect 43466 625163 43472 625215
rect 42160 624645 42166 624697
rect 42218 624685 42224 624697
rect 42448 624685 42454 624697
rect 42218 624657 42454 624685
rect 42218 624645 42224 624657
rect 42448 624645 42454 624657
rect 42506 624645 42512 624697
rect 42160 623461 42166 623513
rect 42218 623501 42224 623513
rect 42928 623501 42934 623513
rect 42218 623473 42934 623501
rect 42218 623461 42224 623473
rect 42928 623461 42934 623473
rect 42986 623461 42992 623513
rect 42448 623313 42454 623365
rect 42506 623353 42512 623365
rect 42928 623353 42934 623365
rect 42506 623325 42934 623353
rect 42506 623313 42512 623325
rect 42928 623313 42934 623325
rect 42986 623313 42992 623365
rect 654448 622055 654454 622107
rect 654506 622095 654512 622107
rect 669904 622095 669910 622107
rect 654506 622067 669910 622095
rect 654506 622055 654512 622067
rect 669904 622055 669910 622067
rect 669962 622055 669968 622107
rect 42160 621611 42166 621663
rect 42218 621651 42224 621663
rect 43024 621651 43030 621663
rect 42218 621623 43030 621651
rect 42218 621611 42224 621623
rect 43024 621611 43030 621623
rect 43082 621611 43088 621663
rect 43024 621463 43030 621515
rect 43082 621503 43088 621515
rect 43504 621503 43510 621515
rect 43082 621475 43510 621503
rect 43082 621463 43088 621475
rect 43504 621463 43510 621475
rect 43562 621463 43568 621515
rect 42160 620353 42166 620405
rect 42218 620393 42224 620405
rect 43120 620393 43126 620405
rect 42218 620365 43126 620393
rect 42218 620353 42224 620365
rect 43120 620353 43126 620365
rect 43178 620353 43184 620405
rect 43120 620205 43126 620257
rect 43178 620245 43184 620257
rect 43600 620245 43606 620257
rect 43178 620217 43606 620245
rect 43178 620205 43184 620217
rect 43600 620205 43606 620217
rect 43658 620205 43664 620257
rect 672208 619169 672214 619221
rect 672266 619209 672272 619221
rect 673840 619209 673846 619221
rect 672266 619181 673846 619209
rect 672266 619169 672272 619181
rect 673840 619169 673846 619181
rect 673898 619169 673904 619221
rect 42064 617837 42070 617889
rect 42122 617877 42128 617889
rect 42448 617877 42454 617889
rect 42122 617849 42454 617877
rect 42122 617837 42128 617849
rect 42448 617837 42454 617849
rect 42506 617837 42512 617889
rect 672112 617837 672118 617889
rect 672170 617877 672176 617889
rect 673840 617877 673846 617889
rect 672170 617849 673846 617877
rect 672170 617837 672176 617849
rect 673840 617837 673846 617849
rect 673898 617837 673904 617889
rect 42160 617171 42166 617223
rect 42218 617211 42224 617223
rect 43120 617211 43126 617223
rect 42218 617183 43126 617211
rect 42218 617171 42224 617183
rect 43120 617171 43126 617183
rect 43178 617171 43184 617223
rect 42160 616653 42166 616705
rect 42218 616693 42224 616705
rect 42928 616693 42934 616705
rect 42218 616665 42934 616693
rect 42218 616653 42224 616665
rect 42928 616653 42934 616665
rect 42986 616653 42992 616705
rect 42160 615839 42166 615891
rect 42218 615879 42224 615891
rect 43024 615879 43030 615891
rect 42218 615851 43030 615879
rect 42218 615839 42224 615851
rect 43024 615839 43030 615851
rect 43082 615839 43088 615891
rect 42160 613989 42166 614041
rect 42218 614029 42224 614041
rect 42832 614029 42838 614041
rect 42218 614001 42838 614029
rect 42218 613989 42224 614001
rect 42832 613989 42838 614001
rect 42890 613989 42896 614041
rect 42160 613619 42166 613671
rect 42218 613659 42224 613671
rect 42448 613659 42454 613671
rect 42218 613631 42454 613659
rect 42218 613619 42224 613631
rect 42448 613619 42454 613631
rect 42506 613619 42512 613671
rect 42448 613471 42454 613523
rect 42506 613511 42512 613523
rect 58384 613511 58390 613523
rect 42506 613483 58390 613511
rect 42506 613471 42512 613483
rect 58384 613471 58390 613483
rect 58442 613471 58448 613523
rect 649840 613471 649846 613523
rect 649898 613511 649904 613523
rect 679696 613511 679702 613523
rect 649898 613483 679702 613511
rect 649898 613471 649904 613483
rect 679696 613471 679702 613483
rect 679754 613471 679760 613523
rect 654448 613397 654454 613449
rect 654506 613437 654512 613449
rect 669520 613437 669526 613449
rect 654506 613409 669526 613437
rect 654506 613397 654512 613409
rect 669520 613397 669526 613409
rect 669578 613397 669584 613449
rect 42064 612805 42070 612857
rect 42122 612845 42128 612857
rect 42736 612845 42742 612857
rect 42122 612817 42742 612845
rect 42122 612805 42128 612817
rect 42736 612805 42742 612817
rect 42794 612805 42800 612857
rect 42736 607699 42742 607751
rect 42794 607739 42800 607751
rect 51856 607739 51862 607751
rect 42794 607711 51862 607739
rect 42794 607699 42800 607711
rect 51856 607699 51862 607711
rect 51914 607699 51920 607751
rect 42736 606811 42742 606863
rect 42794 606851 42800 606863
rect 53392 606851 53398 606863
rect 42794 606823 53398 606851
rect 42794 606811 42800 606823
rect 53392 606811 53398 606823
rect 53450 606811 53456 606863
rect 672208 603629 672214 603681
rect 672266 603669 672272 603681
rect 674608 603669 674614 603681
rect 672266 603641 674614 603669
rect 672266 603629 672272 603641
rect 674608 603629 674614 603641
rect 674666 603669 674672 603681
rect 675280 603669 675286 603681
rect 674666 603641 675286 603669
rect 674666 603629 674672 603641
rect 675280 603629 675286 603641
rect 675338 603629 675344 603681
rect 673744 602815 673750 602867
rect 673802 602855 673808 602867
rect 674800 602855 674806 602867
rect 673802 602827 674806 602855
rect 673802 602815 673808 602827
rect 674800 602815 674806 602827
rect 674858 602855 674864 602867
rect 675472 602855 675478 602867
rect 674858 602827 675478 602855
rect 674858 602815 674864 602827
rect 675472 602815 675478 602827
rect 675530 602815 675536 602867
rect 672016 602667 672022 602719
rect 672074 602707 672080 602719
rect 675376 602707 675382 602719
rect 672074 602679 675382 602707
rect 672074 602667 672080 602679
rect 675376 602667 675382 602679
rect 675434 602667 675440 602719
rect 663760 602075 663766 602127
rect 663818 602115 663824 602127
rect 663818 602087 675326 602115
rect 663818 602075 663824 602087
rect 671824 602001 671830 602053
rect 671882 602041 671888 602053
rect 675184 602041 675190 602053
rect 671882 602013 675190 602041
rect 671882 602001 671888 602013
rect 675184 602001 675190 602013
rect 675242 602001 675248 602053
rect 672112 601927 672118 601979
rect 672170 601967 672176 601979
rect 675088 601967 675094 601979
rect 672170 601939 675094 601967
rect 672170 601927 672176 601939
rect 675088 601927 675094 601939
rect 675146 601927 675152 601979
rect 675298 601967 675326 602087
rect 675202 601939 675326 601967
rect 675202 601905 675230 601939
rect 51856 601853 51862 601905
rect 51914 601893 51920 601905
rect 59536 601893 59542 601905
rect 51914 601865 59542 601893
rect 51914 601853 51920 601865
rect 59536 601853 59542 601865
rect 59594 601853 59600 601905
rect 675184 601853 675190 601905
rect 675242 601853 675248 601905
rect 671344 599781 671350 599833
rect 671402 599821 671408 599833
rect 675376 599821 675382 599833
rect 671402 599793 675382 599821
rect 671402 599781 671408 599793
rect 675376 599781 675382 599793
rect 675434 599781 675440 599833
rect 671536 599263 671542 599315
rect 671594 599303 671600 599315
rect 675376 599303 675382 599315
rect 671594 599275 675382 599303
rect 671594 599263 671600 599275
rect 675376 599263 675382 599275
rect 675434 599263 675440 599315
rect 654448 599041 654454 599093
rect 654506 599081 654512 599093
rect 666832 599081 666838 599093
rect 654506 599053 666838 599081
rect 654506 599041 654512 599053
rect 666832 599041 666838 599053
rect 666890 599041 666896 599093
rect 672688 598375 672694 598427
rect 672746 598415 672752 598427
rect 675472 598415 675478 598427
rect 672746 598387 675478 598415
rect 672746 598375 672752 598387
rect 675472 598375 675478 598387
rect 675530 598375 675536 598427
rect 672496 597117 672502 597169
rect 672554 597157 672560 597169
rect 675472 597157 675478 597169
rect 672554 597129 675478 597157
rect 672554 597117 672560 597129
rect 675472 597117 675478 597129
rect 675530 597117 675536 597169
rect 675184 596821 675190 596873
rect 675242 596861 675248 596873
rect 675376 596861 675382 596873
rect 675242 596833 675382 596861
rect 675242 596821 675248 596833
rect 675376 596821 675382 596833
rect 675434 596821 675440 596873
rect 670864 590309 670870 590361
rect 670922 590349 670928 590361
rect 679696 590349 679702 590361
rect 670922 590321 679702 590349
rect 670922 590309 670928 590321
rect 679696 590309 679702 590321
rect 679754 590309 679760 590361
rect 42544 589199 42550 589251
rect 42602 589239 42608 589251
rect 45232 589239 45238 589251
rect 42602 589211 45238 589239
rect 42602 589199 42608 589211
rect 45232 589199 45238 589211
rect 45290 589199 45296 589251
rect 53392 587423 53398 587475
rect 53450 587463 53456 587475
rect 59536 587463 59542 587475
rect 53450 587435 59542 587463
rect 53450 587423 53456 587435
rect 59536 587423 59542 587435
rect 59594 587423 59600 587475
rect 42544 586535 42550 586587
rect 42602 586575 42608 586587
rect 43024 586575 43030 586587
rect 42602 586547 43030 586575
rect 42602 586535 42608 586547
rect 43024 586535 43030 586547
rect 43082 586535 43088 586587
rect 663952 586313 663958 586365
rect 664010 586353 664016 586365
rect 674416 586353 674422 586365
rect 664010 586325 674422 586353
rect 664010 586313 664016 586325
rect 674416 586313 674422 586325
rect 674474 586313 674480 586365
rect 42448 586091 42454 586143
rect 42506 586131 42512 586143
rect 43024 586131 43030 586143
rect 42506 586103 43030 586131
rect 42506 586091 42512 586103
rect 43024 586091 43030 586103
rect 43082 586091 43088 586143
rect 40048 585943 40054 585995
rect 40106 585983 40112 585995
rect 42448 585983 42454 585995
rect 40106 585955 42454 585983
rect 40106 585943 40112 585955
rect 42448 585943 42454 585955
rect 42506 585943 42512 585995
rect 664144 585425 664150 585477
rect 664202 585465 664208 585477
rect 674416 585465 674422 585477
rect 664202 585437 674422 585465
rect 664202 585425 664208 585437
rect 674416 585425 674422 585437
rect 674474 585425 674480 585477
rect 42832 585055 42838 585107
rect 42890 585095 42896 585107
rect 43120 585095 43126 585107
rect 42890 585067 43126 585095
rect 42890 585055 42896 585067
rect 43120 585055 43126 585067
rect 43178 585055 43184 585107
rect 654448 585055 654454 585107
rect 654506 585095 654512 585107
rect 661168 585095 661174 585107
rect 654506 585067 661174 585095
rect 654506 585055 654512 585067
rect 661168 585055 661174 585067
rect 661226 585055 661232 585107
rect 671728 584833 671734 584885
rect 671786 584873 671792 584885
rect 674608 584873 674614 584885
rect 671786 584845 674614 584873
rect 671786 584833 671792 584845
rect 674608 584833 674614 584845
rect 674666 584833 674672 584885
rect 42544 584759 42550 584811
rect 42602 584799 42608 584811
rect 43120 584799 43126 584811
rect 42602 584771 43126 584799
rect 42602 584759 42608 584771
rect 43120 584759 43126 584771
rect 43178 584759 43184 584811
rect 655120 584759 655126 584811
rect 655178 584799 655184 584811
rect 674704 584799 674710 584811
rect 655178 584771 674710 584799
rect 655178 584759 655184 584771
rect 674704 584759 674710 584771
rect 674762 584759 674768 584811
rect 42832 584685 42838 584737
rect 42890 584725 42896 584737
rect 50512 584725 50518 584737
rect 42890 584697 50518 584725
rect 42890 584685 42896 584697
rect 50512 584685 50518 584697
rect 50570 584685 50576 584737
rect 41776 584167 41782 584219
rect 41834 584167 41840 584219
rect 42160 584167 42166 584219
rect 42218 584207 42224 584219
rect 42928 584207 42934 584219
rect 42218 584179 42934 584207
rect 42218 584167 42224 584179
rect 42928 584167 42934 584179
rect 42986 584167 42992 584219
rect 41794 583997 41822 584167
rect 41776 583945 41782 583997
rect 41834 583945 41840 583997
rect 672400 583575 672406 583627
rect 672458 583615 672464 583627
rect 674704 583615 674710 583627
rect 672458 583587 674710 583615
rect 672458 583575 672464 583587
rect 674704 583575 674710 583587
rect 674762 583575 674768 583627
rect 670960 583353 670966 583405
rect 671018 583393 671024 583405
rect 674704 583393 674710 583405
rect 671018 583365 674710 583393
rect 671018 583353 671024 583365
rect 674704 583353 674710 583365
rect 674762 583393 674768 583405
rect 679984 583393 679990 583405
rect 674762 583365 679990 583393
rect 674762 583353 674768 583365
rect 679984 583353 679990 583365
rect 680042 583353 680048 583405
rect 42160 582095 42166 582147
rect 42218 582135 42224 582147
rect 42448 582135 42454 582147
rect 42218 582107 42454 582135
rect 42218 582095 42224 582107
rect 42448 582095 42454 582107
rect 42506 582095 42512 582147
rect 42064 581429 42070 581481
rect 42122 581469 42128 581481
rect 42832 581469 42838 581481
rect 42122 581441 42838 581469
rect 42122 581429 42128 581441
rect 42832 581429 42838 581441
rect 42890 581429 42896 581481
rect 42064 580245 42070 580297
rect 42122 580285 42128 580297
rect 43216 580285 43222 580297
rect 42122 580257 43222 580285
rect 42122 580245 42128 580257
rect 43216 580245 43222 580257
rect 43274 580245 43280 580297
rect 43312 580023 43318 580075
rect 43370 580063 43376 580075
rect 43600 580063 43606 580075
rect 43370 580035 43606 580063
rect 43370 580023 43376 580035
rect 43600 580023 43606 580035
rect 43658 580023 43664 580075
rect 42160 578987 42166 579039
rect 42218 579027 42224 579039
rect 43120 579027 43126 579039
rect 42218 578999 43126 579027
rect 42218 578987 42224 578999
rect 43120 578987 43126 578999
rect 43178 578987 43184 579039
rect 672400 578839 672406 578891
rect 672458 578879 672464 578891
rect 672784 578879 672790 578891
rect 672458 578851 672790 578879
rect 672458 578839 672464 578851
rect 672784 578839 672790 578851
rect 672842 578839 672848 578891
rect 42064 578395 42070 578447
rect 42122 578435 42128 578447
rect 42928 578435 42934 578447
rect 42122 578407 42934 578435
rect 42122 578395 42128 578407
rect 42928 578395 42934 578407
rect 42986 578395 42992 578447
rect 42160 577655 42166 577707
rect 42218 577695 42224 577707
rect 43024 577695 43030 577707
rect 42218 577667 43030 577695
rect 42218 577655 42224 577667
rect 43024 577655 43030 577667
rect 43082 577655 43088 577707
rect 42256 576027 42262 576079
rect 42314 576067 42320 576079
rect 42928 576067 42934 576079
rect 42314 576039 42934 576067
rect 42314 576027 42320 576039
rect 42928 576027 42934 576039
rect 42986 576027 42992 576079
rect 671920 575361 671926 575413
rect 671978 575401 671984 575413
rect 674704 575401 674710 575413
rect 671978 575373 674710 575401
rect 671978 575361 671984 575373
rect 674704 575361 674710 575373
rect 674762 575361 674768 575413
rect 671440 574473 671446 574525
rect 671498 574513 671504 574525
rect 674704 574513 674710 574525
rect 671498 574485 674710 574513
rect 671498 574473 671504 574485
rect 674704 574473 674710 574485
rect 674762 574473 674768 574525
rect 672304 573585 672310 573637
rect 672362 573625 672368 573637
rect 674416 573625 674422 573637
rect 672362 573597 674422 573625
rect 672362 573585 672368 573597
rect 674416 573585 674422 573597
rect 674474 573585 674480 573637
rect 42064 573437 42070 573489
rect 42122 573477 42128 573489
rect 42832 573477 42838 573489
rect 42122 573449 42838 573477
rect 42122 573437 42128 573449
rect 42832 573437 42838 573449
rect 42890 573437 42896 573489
rect 654448 573141 654454 573193
rect 654506 573181 654512 573193
rect 663952 573181 663958 573193
rect 654506 573153 663958 573181
rect 654506 573141 654512 573153
rect 663952 573141 663958 573153
rect 664010 573141 664016 573193
rect 672880 572993 672886 573045
rect 672938 573033 672944 573045
rect 674704 573033 674710 573045
rect 672938 573005 674710 573033
rect 672938 572993 672944 573005
rect 674704 572993 674710 573005
rect 674762 572993 674768 573045
rect 42160 572623 42166 572675
rect 42218 572663 42224 572675
rect 42448 572663 42454 572675
rect 42218 572635 42454 572663
rect 42218 572623 42224 572635
rect 42448 572623 42454 572635
rect 42506 572623 42512 572675
rect 42256 572475 42262 572527
rect 42314 572515 42320 572527
rect 42448 572515 42454 572527
rect 42314 572487 42454 572515
rect 42314 572475 42320 572487
rect 42448 572475 42454 572487
rect 42506 572475 42512 572527
rect 671632 571957 671638 572009
rect 671690 571997 671696 572009
rect 674416 571997 674422 572009
rect 671690 571969 674422 571997
rect 671690 571957 671696 571969
rect 674416 571957 674422 571969
rect 674474 571957 674480 572009
rect 672592 571365 672598 571417
rect 672650 571405 672656 571417
rect 674704 571405 674710 571417
rect 672650 571377 674710 571405
rect 672650 571365 672656 571377
rect 674704 571365 674710 571377
rect 674762 571365 674768 571417
rect 42160 570995 42166 571047
rect 42218 571035 42224 571047
rect 43024 571035 43030 571047
rect 42218 571007 43030 571035
rect 42218 570995 42224 571007
rect 43024 570995 43030 571007
rect 43082 570995 43088 571047
rect 42352 570255 42358 570307
rect 42410 570295 42416 570307
rect 59536 570295 59542 570307
rect 42410 570267 59542 570295
rect 42410 570255 42416 570267
rect 59536 570255 59542 570267
rect 59594 570255 59600 570307
rect 42064 570181 42070 570233
rect 42122 570221 42128 570233
rect 42448 570221 42454 570233
rect 42122 570193 42454 570221
rect 42122 570181 42128 570193
rect 42448 570181 42454 570193
rect 42506 570181 42512 570233
rect 42064 569663 42070 569715
rect 42122 569703 42128 569715
rect 42832 569703 42838 569715
rect 42122 569675 42838 569703
rect 42122 569663 42128 569675
rect 42832 569663 42838 569675
rect 42890 569663 42896 569715
rect 649936 567369 649942 567421
rect 649994 567409 650000 567421
rect 679792 567409 679798 567421
rect 649994 567381 679798 567409
rect 649994 567369 650000 567381
rect 679792 567369 679798 567381
rect 679850 567369 679856 567421
rect 34480 564483 34486 564535
rect 34538 564523 34544 564535
rect 53392 564523 53398 564535
rect 34538 564495 53398 564523
rect 34538 564483 34544 564495
rect 53392 564483 53398 564495
rect 53450 564483 53456 564535
rect 654448 564409 654454 564461
rect 654506 564449 654512 564461
rect 666640 564449 666646 564461
rect 654506 564421 666646 564449
rect 654506 564409 654512 564421
rect 666640 564409 666646 564421
rect 666698 564409 666704 564461
rect 672208 564409 672214 564461
rect 672266 564449 672272 564461
rect 674992 564449 674998 564461
rect 672266 564421 674998 564449
rect 672266 564409 672272 564421
rect 674992 564409 674998 564421
rect 675050 564409 675056 564461
rect 42448 563447 42454 563499
rect 42506 563487 42512 563499
rect 50512 563487 50518 563499
rect 42506 563459 50518 563487
rect 42506 563447 42512 563459
rect 50512 563447 50518 563459
rect 50570 563447 50576 563499
rect 673744 561597 673750 561649
rect 673802 561637 673808 561649
rect 675088 561637 675094 561649
rect 673802 561609 675094 561637
rect 673802 561597 673808 561609
rect 675088 561597 675094 561609
rect 675146 561597 675152 561649
rect 674224 559525 674230 559577
rect 674282 559565 674288 559577
rect 675376 559565 675382 559577
rect 674282 559537 675382 559565
rect 674282 559525 674288 559537
rect 675376 559525 675382 559537
rect 675434 559525 675440 559577
rect 672208 558711 672214 558763
rect 672266 558751 672272 558763
rect 672784 558751 672790 558763
rect 672266 558723 672790 558751
rect 672266 558711 672272 558723
rect 672784 558711 672790 558723
rect 672842 558711 672848 558763
rect 53392 558637 53398 558689
rect 53450 558677 53456 558689
rect 59536 558677 59542 558689
rect 53450 558649 59542 558677
rect 53450 558637 53456 558649
rect 59536 558637 59542 558649
rect 59594 558637 59600 558689
rect 674128 558045 674134 558097
rect 674186 558085 674192 558097
rect 675376 558085 675382 558097
rect 674186 558057 675382 558085
rect 674186 558045 674192 558057
rect 675376 558045 675382 558057
rect 675434 558045 675440 558097
rect 660880 555825 660886 555877
rect 660938 555865 660944 555877
rect 675184 555865 675190 555877
rect 660938 555837 675190 555865
rect 660938 555825 660944 555837
rect 675184 555825 675190 555837
rect 675242 555825 675248 555877
rect 674320 555011 674326 555063
rect 674378 555051 674384 555063
rect 675472 555051 675478 555063
rect 674378 555023 675478 555051
rect 674378 555011 674384 555023
rect 675472 555011 675478 555023
rect 675530 555011 675536 555063
rect 674032 554493 674038 554545
rect 674090 554533 674096 554545
rect 675376 554533 675382 554545
rect 674090 554505 675382 554533
rect 674090 554493 674096 554505
rect 675376 554493 675382 554505
rect 675434 554493 675440 554545
rect 674992 553901 674998 553953
rect 675050 553941 675056 553953
rect 675472 553941 675478 553953
rect 675050 553913 675478 553941
rect 675050 553901 675056 553913
rect 675472 553901 675478 553913
rect 675530 553901 675536 553953
rect 674896 553161 674902 553213
rect 674954 553201 674960 553213
rect 675376 553201 675382 553213
rect 674954 553173 675382 553201
rect 674954 553161 674960 553173
rect 675376 553161 675382 553173
rect 675434 553161 675440 553213
rect 674512 551903 674518 551955
rect 674570 551943 674576 551955
rect 675472 551943 675478 551955
rect 674570 551915 675478 551943
rect 674570 551903 674576 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 675184 551533 675190 551585
rect 675242 551573 675248 551585
rect 675376 551573 675382 551585
rect 675242 551545 675382 551573
rect 675242 551533 675248 551545
rect 675376 551533 675382 551545
rect 675434 551533 675440 551585
rect 654448 550127 654454 550179
rect 654506 550167 654512 550179
rect 661072 550167 661078 550179
rect 654506 550139 661078 550167
rect 654506 550127 654512 550139
rect 661072 550127 661078 550139
rect 661130 550127 661136 550179
rect 674608 550053 674614 550105
rect 674666 550093 674672 550105
rect 675472 550093 675478 550105
rect 674666 550065 675478 550093
rect 674666 550053 674672 550065
rect 675472 550053 675478 550065
rect 675530 550053 675536 550105
rect 674800 548203 674806 548255
rect 674858 548243 674864 548255
rect 675376 548243 675382 548255
rect 674858 548215 675382 548243
rect 674858 548203 674864 548215
rect 675376 548203 675382 548215
rect 675434 548203 675440 548255
rect 42640 546205 42646 546257
rect 42698 546245 42704 546257
rect 45328 546245 45334 546257
rect 42698 546217 45334 546245
rect 42698 546205 42704 546217
rect 45328 546205 45334 546217
rect 45386 546205 45392 546257
rect 42352 545539 42358 545591
rect 42410 545579 42416 545591
rect 42640 545579 42646 545591
rect 42410 545551 42646 545579
rect 42410 545539 42416 545551
rect 42640 545539 42646 545551
rect 42698 545539 42704 545591
rect 41968 544577 41974 544629
rect 42026 544617 42032 544629
rect 42928 544617 42934 544629
rect 42026 544589 42934 544617
rect 42026 544577 42032 544589
rect 42928 544577 42934 544589
rect 42986 544577 42992 544629
rect 50512 543689 50518 543741
rect 50570 543729 50576 543741
rect 59536 543729 59542 543741
rect 50570 543701 59542 543729
rect 50570 543689 50576 543701
rect 59536 543689 59542 543701
rect 59594 543689 59600 543741
rect 40144 542875 40150 542927
rect 40202 542915 40208 542927
rect 41968 542915 41974 542927
rect 40202 542887 41974 542915
rect 40202 542875 40208 542887
rect 41968 542875 41974 542887
rect 42026 542875 42032 542927
rect 43696 541469 43702 541521
rect 43754 541509 43760 541521
rect 53296 541509 53302 541521
rect 43754 541481 53302 541509
rect 43754 541469 43760 541481
rect 53296 541469 53302 541481
rect 53354 541469 53360 541521
rect 655312 541469 655318 541521
rect 655370 541509 655376 541521
rect 674704 541509 674710 541521
rect 655370 541481 674710 541509
rect 655370 541469 655376 541481
rect 674704 541469 674710 541481
rect 674762 541469 674768 541521
rect 666928 541321 666934 541373
rect 666986 541361 666992 541373
rect 674416 541361 674422 541373
rect 666986 541333 674422 541361
rect 666986 541321 666992 541333
rect 674416 541321 674422 541333
rect 674474 541321 674480 541373
rect 41680 541247 41686 541299
rect 41738 541287 41744 541299
rect 43408 541287 43414 541299
rect 41738 541259 43414 541287
rect 41738 541247 41744 541259
rect 43408 541247 43414 541259
rect 43466 541247 43472 541299
rect 674320 541025 674326 541077
rect 674378 541065 674384 541077
rect 674992 541065 674998 541077
rect 674378 541037 674998 541065
rect 674378 541025 674384 541037
rect 674992 541025 674998 541037
rect 675050 541025 675056 541077
rect 41776 540951 41782 541003
rect 41834 540951 41840 541003
rect 42160 540951 42166 541003
rect 42218 540991 42224 541003
rect 43312 540991 43318 541003
rect 42218 540963 43318 540991
rect 42218 540951 42224 540963
rect 43312 540951 43318 540963
rect 43370 540951 43376 541003
rect 41794 540781 41822 540951
rect 41776 540729 41782 540781
rect 41834 540729 41840 540781
rect 661264 540729 661270 540781
rect 661322 540769 661328 540781
rect 674704 540769 674710 540781
rect 661322 540741 674710 540769
rect 661322 540729 661328 540741
rect 674704 540729 674710 540741
rect 674762 540729 674768 540781
rect 672208 539841 672214 539893
rect 672266 539881 672272 539893
rect 674704 539881 674710 539893
rect 672266 539853 674710 539881
rect 672266 539841 672272 539853
rect 674704 539841 674710 539853
rect 674762 539841 674768 539893
rect 42928 538731 42934 538783
rect 42986 538771 42992 538783
rect 43504 538771 43510 538783
rect 42986 538743 43510 538771
rect 42986 538731 42992 538743
rect 43504 538731 43510 538743
rect 43562 538731 43568 538783
rect 42160 538139 42166 538191
rect 42218 538179 42224 538191
rect 43696 538179 43702 538191
rect 42218 538151 43702 538179
rect 42218 538139 42224 538151
rect 43696 538139 43702 538151
rect 43754 538139 43760 538191
rect 42064 537029 42070 537081
rect 42122 537069 42128 537081
rect 42832 537069 42838 537081
rect 42122 537041 42838 537069
rect 42122 537029 42128 537041
rect 42832 537029 42838 537041
rect 42890 537029 42896 537081
rect 42064 535771 42070 535823
rect 42122 535811 42128 535823
rect 43120 535811 43126 535823
rect 42122 535783 43126 535811
rect 42122 535771 42128 535783
rect 43120 535771 43126 535783
rect 43178 535771 43184 535823
rect 43216 535771 43222 535823
rect 43274 535771 43280 535823
rect 43234 535601 43262 535771
rect 676624 535697 676630 535749
rect 676682 535737 676688 535749
rect 679792 535737 679798 535749
rect 676682 535709 679798 535737
rect 676682 535697 676688 535709
rect 679792 535697 679798 535709
rect 679850 535697 679856 535749
rect 43216 535549 43222 535601
rect 43274 535549 43280 535601
rect 42160 535253 42166 535305
rect 42218 535293 42224 535305
rect 42736 535293 42742 535305
rect 42218 535265 42742 535293
rect 42218 535253 42224 535265
rect 42736 535253 42742 535265
rect 42794 535253 42800 535305
rect 42160 534439 42166 534491
rect 42218 534479 42224 534491
rect 43024 534479 43030 534491
rect 42218 534451 43030 534479
rect 42218 534439 42224 534451
rect 43024 534439 43030 534451
rect 43082 534439 43088 534491
rect 43024 534291 43030 534343
rect 43082 534331 43088 534343
rect 43408 534331 43414 534343
rect 43082 534303 43414 534331
rect 43082 534291 43088 534303
rect 43408 534291 43414 534303
rect 43466 534291 43472 534343
rect 42064 533699 42070 533751
rect 42122 533739 42128 533751
rect 42928 533739 42934 533751
rect 42122 533711 42934 533739
rect 42122 533699 42128 533711
rect 42928 533699 42934 533711
rect 42986 533699 42992 533751
rect 42928 533551 42934 533603
rect 42986 533591 42992 533603
rect 43504 533591 43510 533603
rect 42986 533563 43510 533591
rect 42986 533551 42992 533563
rect 43504 533551 43510 533563
rect 43562 533551 43568 533603
rect 42256 532811 42262 532863
rect 42314 532851 42320 532863
rect 42640 532851 42646 532863
rect 42314 532823 42646 532851
rect 42314 532811 42320 532823
rect 42640 532811 42646 532823
rect 42698 532811 42704 532863
rect 672112 532737 672118 532789
rect 672170 532777 672176 532789
rect 673840 532777 673846 532789
rect 672170 532749 673846 532777
rect 672170 532737 672176 532749
rect 673840 532737 673846 532749
rect 673898 532737 673904 532789
rect 42160 531331 42166 531383
rect 42218 531371 42224 531383
rect 43120 531371 43126 531383
rect 42218 531343 43126 531371
rect 42218 531331 42224 531343
rect 43120 531331 43126 531343
rect 43178 531331 43184 531383
rect 671824 530813 671830 530865
rect 671882 530853 671888 530865
rect 673840 530853 673846 530865
rect 671882 530825 673846 530853
rect 671882 530813 671888 530825
rect 673840 530813 673846 530825
rect 673898 530813 673904 530865
rect 42256 530295 42262 530347
rect 42314 530335 42320 530347
rect 42832 530335 42838 530347
rect 42314 530307 42838 530335
rect 42314 530295 42320 530307
rect 42832 530295 42838 530307
rect 42890 530295 42896 530347
rect 672496 529851 672502 529903
rect 672554 529891 672560 529903
rect 673840 529891 673846 529903
rect 672554 529863 673846 529891
rect 672554 529851 672560 529863
rect 673840 529851 673846 529863
rect 673898 529851 673904 529903
rect 671536 529777 671542 529829
rect 671594 529817 671600 529829
rect 673744 529817 673750 529829
rect 671594 529789 673750 529817
rect 671594 529777 671600 529789
rect 673744 529777 673750 529789
rect 673802 529777 673808 529829
rect 42256 529629 42262 529681
rect 42314 529669 42320 529681
rect 43024 529669 43030 529681
rect 42314 529641 43030 529669
rect 42314 529629 42320 529641
rect 43024 529629 43030 529641
rect 43082 529629 43088 529681
rect 672016 529185 672022 529237
rect 672074 529225 672080 529237
rect 673840 529225 673846 529237
rect 672074 529197 673846 529225
rect 672074 529185 672080 529197
rect 673840 529185 673846 529197
rect 673898 529185 673904 529237
rect 42160 527631 42166 527683
rect 42218 527671 42224 527683
rect 42928 527671 42934 527683
rect 42218 527643 42934 527671
rect 42218 527631 42224 527643
rect 42928 527631 42934 527643
rect 42986 527631 42992 527683
rect 42064 527187 42070 527239
rect 42122 527227 42128 527239
rect 42640 527227 42646 527239
rect 42122 527199 42646 527227
rect 42122 527187 42128 527199
rect 42640 527187 42646 527199
rect 42698 527187 42704 527239
rect 42352 527039 42358 527091
rect 42410 527079 42416 527091
rect 59440 527079 59446 527091
rect 42410 527051 59446 527079
rect 42410 527039 42416 527051
rect 59440 527039 59446 527051
rect 59498 527039 59504 527091
rect 654448 527039 654454 527091
rect 654506 527079 654512 527091
rect 669808 527079 669814 527091
rect 654506 527051 669814 527079
rect 654506 527039 654512 527051
rect 669808 527039 669814 527051
rect 669866 527039 669872 527091
rect 672688 526891 672694 526943
rect 672746 526931 672752 526943
rect 673840 526931 673846 526943
rect 672746 526903 673846 526931
rect 672746 526891 672752 526903
rect 673840 526891 673846 526903
rect 673898 526891 673904 526943
rect 671344 526817 671350 526869
rect 671402 526857 671408 526869
rect 673744 526857 673750 526869
rect 671402 526829 673750 526857
rect 671402 526817 671408 526829
rect 673744 526817 673750 526829
rect 673802 526817 673808 526869
rect 42160 526447 42166 526499
rect 42218 526487 42224 526499
rect 42736 526487 42742 526499
rect 42218 526459 42742 526487
rect 42218 526447 42224 526459
rect 42736 526447 42742 526459
rect 42794 526447 42800 526499
rect 650032 521267 650038 521319
rect 650090 521307 650096 521319
rect 679792 521307 679798 521319
rect 650090 521279 679798 521307
rect 650090 521267 650096 521279
rect 679792 521267 679798 521279
rect 679850 521267 679856 521319
rect 654448 517937 654454 517989
rect 654506 517977 654512 517989
rect 663856 517977 663862 517989
rect 654506 517949 663862 517977
rect 654506 517937 654512 517949
rect 663856 517937 663862 517949
rect 663914 517937 663920 517989
rect 50608 512683 50614 512735
rect 50666 512723 50672 512735
rect 59536 512723 59542 512735
rect 50666 512695 59542 512723
rect 50666 512683 50672 512695
rect 59536 512683 59542 512695
rect 59594 512683 59600 512735
rect 654448 504025 654454 504077
rect 654506 504065 654512 504077
rect 666640 504065 666646 504077
rect 654506 504037 666646 504065
rect 654506 504025 654512 504037
rect 666640 504025 666646 504037
rect 666698 504025 666704 504077
rect 53392 498253 53398 498305
rect 53450 498293 53456 498305
rect 58096 498293 58102 498305
rect 53450 498265 58102 498293
rect 53450 498253 53456 498265
rect 58096 498253 58102 498265
rect 58154 498253 58160 498305
rect 674032 498031 674038 498083
rect 674090 498071 674096 498083
rect 674992 498071 674998 498083
rect 674090 498043 674998 498071
rect 674090 498031 674096 498043
rect 674992 498031 674998 498043
rect 675050 498031 675056 498083
rect 674224 497883 674230 497935
rect 674282 497883 674288 497935
rect 674704 497883 674710 497935
rect 674762 497923 674768 497935
rect 674896 497923 674902 497935
rect 674762 497895 674902 497923
rect 674762 497883 674768 497895
rect 674896 497883 674902 497895
rect 674954 497883 674960 497935
rect 674242 497713 674270 497883
rect 674224 497661 674230 497713
rect 674282 497661 674288 497713
rect 674320 497587 674326 497639
rect 674378 497627 674384 497639
rect 674512 497627 674518 497639
rect 674378 497599 674518 497627
rect 674378 497587 674384 497599
rect 674512 497587 674518 497599
rect 674570 497587 674576 497639
rect 669712 497291 669718 497343
rect 669770 497331 669776 497343
rect 674416 497331 674422 497343
rect 669770 497303 674422 497331
rect 669770 497291 669776 497303
rect 674416 497291 674422 497303
rect 674474 497291 674480 497343
rect 669904 496477 669910 496529
rect 669962 496517 669968 496529
rect 674416 496517 674422 496529
rect 669962 496489 674422 496517
rect 669962 496477 669968 496489
rect 674416 496477 674422 496489
rect 674474 496477 674480 496529
rect 655216 495515 655222 495567
rect 655274 495555 655280 495567
rect 674704 495555 674710 495567
rect 655274 495527 674710 495555
rect 655274 495515 655280 495527
rect 674704 495515 674710 495527
rect 674762 495515 674768 495567
rect 674800 494257 674806 494309
rect 674858 494297 674864 494309
rect 679696 494297 679702 494309
rect 674858 494269 679702 494297
rect 674858 494257 674864 494269
rect 679696 494257 679702 494269
rect 679754 494257 679760 494309
rect 654448 492481 654454 492533
rect 654506 492521 654512 492533
rect 663856 492521 663862 492533
rect 654506 492493 663862 492521
rect 654506 492481 654512 492493
rect 663856 492481 663862 492493
rect 663914 492481 663920 492533
rect 53296 483823 53302 483875
rect 53354 483863 53360 483875
rect 59536 483863 59542 483875
rect 53354 483835 59542 483863
rect 53354 483823 53360 483835
rect 59536 483823 59542 483835
rect 59594 483823 59600 483875
rect 654448 480937 654454 480989
rect 654506 480977 654512 480989
rect 666928 480977 666934 480989
rect 654506 480949 666934 480977
rect 654506 480937 654512 480949
rect 666928 480937 666934 480949
rect 666986 480937 666992 480989
rect 650128 478125 650134 478177
rect 650186 478165 650192 478177
rect 679792 478165 679798 478177
rect 650186 478137 679798 478165
rect 650186 478125 650192 478137
rect 679792 478125 679798 478137
rect 679850 478125 679856 478177
rect 654448 469985 654454 470037
rect 654506 470025 654512 470037
rect 660976 470025 660982 470037
rect 654506 469997 660982 470025
rect 654506 469985 654512 469997
rect 660976 469985 660982 469997
rect 661034 469985 661040 470037
rect 50512 469467 50518 469519
rect 50570 469507 50576 469519
rect 59536 469507 59542 469519
rect 50570 469479 59542 469507
rect 50570 469467 50576 469479
rect 59536 469467 59542 469479
rect 59594 469467 59600 469519
rect 654352 457923 654358 457975
rect 654410 457963 654416 457975
rect 660976 457963 660982 457975
rect 654410 457935 660982 457963
rect 654410 457923 654416 457935
rect 660976 457923 660982 457935
rect 661034 457923 661040 457975
rect 45424 455037 45430 455089
rect 45482 455077 45488 455089
rect 59536 455077 59542 455089
rect 45482 455049 59542 455077
rect 45482 455037 45488 455049
rect 59536 455037 59542 455049
rect 59594 455037 59600 455089
rect 654448 446379 654454 446431
rect 654506 446419 654512 446431
rect 669712 446419 669718 446431
rect 654506 446391 669718 446419
rect 654506 446379 654512 446391
rect 669712 446379 669718 446391
rect 669770 446379 669776 446431
rect 45520 440681 45526 440733
rect 45578 440721 45584 440733
rect 59536 440721 59542 440733
rect 45578 440693 59542 440721
rect 45578 440681 45584 440693
rect 59536 440681 59542 440693
rect 59594 440681 59600 440733
rect 42640 436907 42646 436959
rect 42698 436947 42704 436959
rect 50608 436947 50614 436959
rect 42698 436919 50614 436947
rect 42698 436907 42704 436919
rect 50608 436907 50614 436919
rect 50666 436907 50672 436959
rect 42640 436093 42646 436145
rect 42698 436133 42704 436145
rect 53392 436133 53398 436145
rect 42698 436105 53398 436133
rect 42698 436093 42704 436105
rect 53392 436093 53398 436105
rect 53450 436093 53456 436145
rect 654352 432023 654358 432075
rect 654410 432063 654416 432075
rect 664048 432063 664054 432075
rect 654410 432035 664054 432063
rect 654410 432023 654416 432035
rect 664048 432023 664054 432035
rect 664106 432023 664112 432075
rect 53392 426251 53398 426303
rect 53450 426291 53456 426303
rect 59344 426291 59350 426303
rect 53450 426263 59350 426291
rect 53450 426251 53456 426263
rect 59344 426251 59350 426263
rect 59402 426251 59408 426303
rect 654448 423291 654454 423343
rect 654506 423331 654512 423343
rect 669616 423331 669622 423343
rect 654506 423303 669622 423331
rect 654506 423291 654512 423303
rect 669616 423291 669622 423303
rect 669674 423291 669680 423343
rect 41872 419961 41878 420013
rect 41930 420001 41936 420013
rect 42352 420001 42358 420013
rect 41930 419973 42358 420001
rect 41930 419961 41936 419973
rect 42352 419961 42358 419973
rect 42410 419961 42416 420013
rect 42640 418555 42646 418607
rect 42698 418595 42704 418607
rect 44656 418595 44662 418607
rect 42698 418567 44662 418595
rect 42698 418555 42704 418567
rect 44656 418555 44662 418567
rect 44714 418555 44720 418607
rect 42160 413523 42166 413575
rect 42218 413563 42224 413575
rect 43216 413563 43222 413575
rect 42218 413535 43222 413563
rect 42218 413523 42224 413535
rect 43216 413523 43222 413535
rect 43274 413523 43280 413575
rect 41776 413375 41782 413427
rect 41834 413375 41840 413427
rect 41794 413205 41822 413375
rect 41776 413153 41782 413205
rect 41834 413153 41840 413205
rect 53488 411821 53494 411873
rect 53546 411861 53552 411873
rect 57808 411861 57814 411873
rect 53546 411833 57814 411861
rect 53546 411821 53552 411833
rect 57808 411821 57814 411833
rect 57866 411821 57872 411873
rect 42160 411303 42166 411355
rect 42218 411343 42224 411355
rect 42352 411343 42358 411355
rect 42218 411315 42358 411343
rect 42218 411303 42224 411315
rect 42352 411303 42358 411315
rect 42410 411303 42416 411355
rect 42352 411155 42358 411207
rect 42410 411195 42416 411207
rect 43120 411195 43126 411207
rect 42410 411167 43126 411195
rect 42410 411155 42416 411167
rect 43120 411155 43126 411167
rect 43178 411155 43184 411207
rect 42064 410489 42070 410541
rect 42122 410529 42128 410541
rect 47440 410529 47446 410541
rect 42122 410501 47446 410529
rect 42122 410489 42128 410501
rect 47440 410489 47446 410501
rect 47498 410489 47504 410541
rect 661168 409897 661174 409949
rect 661226 409937 661232 409949
rect 674416 409937 674422 409949
rect 661226 409909 674422 409937
rect 661226 409897 661232 409909
rect 674416 409897 674422 409909
rect 674474 409897 674480 409949
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42736 409493 42742 409505
rect 42218 409465 42742 409493
rect 42218 409453 42224 409465
rect 42736 409453 42742 409465
rect 42794 409453 42800 409505
rect 666832 409305 666838 409357
rect 666890 409345 666896 409357
rect 674704 409345 674710 409357
rect 666890 409317 674710 409345
rect 666890 409305 666896 409317
rect 674704 409305 674710 409317
rect 674762 409305 674768 409357
rect 655024 408935 655030 408987
rect 655082 408975 655088 408987
rect 669520 408975 669526 408987
rect 655082 408947 669526 408975
rect 655082 408935 655088 408947
rect 669520 408935 669526 408947
rect 669578 408935 669584 408987
rect 663952 408417 663958 408469
rect 664010 408457 664016 408469
rect 674704 408457 674710 408469
rect 664010 408429 674710 408457
rect 664010 408417 664016 408429
rect 674704 408417 674710 408429
rect 674762 408417 674768 408469
rect 42160 408195 42166 408247
rect 42218 408235 42224 408247
rect 42832 408235 42838 408247
rect 42218 408207 42838 408235
rect 42218 408195 42224 408207
rect 42832 408195 42838 408207
rect 42890 408195 42896 408247
rect 42064 407455 42070 407507
rect 42122 407495 42128 407507
rect 43120 407495 43126 407507
rect 42122 407467 43126 407495
rect 42122 407455 42128 407467
rect 43120 407455 43126 407467
rect 43178 407455 43184 407507
rect 42160 406863 42166 406915
rect 42218 406903 42224 406915
rect 43024 406903 43030 406915
rect 42218 406875 43030 406903
rect 42218 406863 42224 406875
rect 43024 406863 43030 406875
rect 43082 406863 43088 406915
rect 42160 403829 42166 403881
rect 42218 403869 42224 403881
rect 42928 403869 42934 403881
rect 42218 403841 42934 403869
rect 42218 403829 42224 403841
rect 42928 403829 42934 403841
rect 42986 403829 42992 403881
rect 42064 402941 42070 402993
rect 42122 402981 42128 402993
rect 42352 402981 42358 402993
rect 42122 402953 42358 402981
rect 42122 402941 42128 402953
rect 42352 402941 42358 402953
rect 42410 402941 42416 402993
rect 654448 397465 654454 397517
rect 654506 397505 654512 397517
rect 663952 397505 663958 397517
rect 654506 397477 663958 397505
rect 654506 397465 654512 397477
rect 663952 397465 663958 397477
rect 664010 397465 664016 397517
rect 42352 393913 42358 393965
rect 42410 393953 42416 393965
rect 50512 393953 50518 393965
rect 42410 393925 50518 393953
rect 42410 393913 42416 393925
rect 50512 393913 50518 393925
rect 50570 393913 50576 393965
rect 42352 393173 42358 393225
rect 42410 393213 42416 393225
rect 45424 393213 45430 393225
rect 42410 393185 45430 393213
rect 42410 393173 42416 393185
rect 45424 393173 45430 393185
rect 45482 393173 45488 393225
rect 42352 392285 42358 392337
rect 42410 392325 42416 392337
rect 53296 392325 53302 392337
rect 42410 392297 53302 392325
rect 42410 392285 42416 392297
rect 53296 392285 53302 392297
rect 53354 392285 53360 392337
rect 650224 391693 650230 391745
rect 650282 391733 650288 391745
rect 679792 391733 679798 391745
rect 650282 391705 679798 391733
rect 650282 391693 650288 391705
rect 679792 391693 679798 391705
rect 679850 391693 679856 391745
rect 653872 385921 653878 385973
rect 653930 385961 653936 385973
rect 669616 385961 669622 385973
rect 653930 385933 669622 385961
rect 653930 385921 653936 385933
rect 669616 385921 669622 385933
rect 669674 385921 669680 385973
rect 674320 384293 674326 384345
rect 674378 384333 674384 384345
rect 675088 384333 675094 384345
rect 674378 384305 675094 384333
rect 674378 384293 674384 384305
rect 675088 384293 675094 384305
rect 675146 384293 675152 384345
rect 674128 383109 674134 383161
rect 674186 383149 674192 383161
rect 675376 383149 675382 383161
rect 674186 383121 675382 383149
rect 674186 383109 674192 383121
rect 675376 383109 675382 383121
rect 675434 383109 675440 383161
rect 45712 383035 45718 383087
rect 45770 383075 45776 383087
rect 59536 383075 59542 383087
rect 45770 383047 59542 383075
rect 45770 383035 45776 383047
rect 59536 383035 59542 383047
rect 59594 383035 59600 383087
rect 674608 382443 674614 382495
rect 674666 382483 674672 382495
rect 675472 382483 675478 382495
rect 674666 382455 675478 382483
rect 674666 382443 674672 382455
rect 675472 382443 675478 382455
rect 675530 382443 675536 382495
rect 674704 378151 674710 378203
rect 674762 378191 674768 378203
rect 675376 378191 675382 378203
rect 674762 378163 675382 378191
rect 674762 378151 674768 378163
rect 675376 378151 675382 378163
rect 675434 378151 675440 378203
rect 674416 377559 674422 377611
rect 674474 377599 674480 377611
rect 675376 377599 675382 377611
rect 674474 377571 675382 377599
rect 674474 377559 674480 377571
rect 675376 377559 675382 377571
rect 675434 377559 675440 377611
rect 654160 377189 654166 377241
rect 654218 377229 654224 377241
rect 666736 377229 666742 377241
rect 654218 377201 666742 377229
rect 654218 377189 654224 377201
rect 666736 377189 666742 377201
rect 666794 377189 666800 377241
rect 674512 376819 674518 376871
rect 674570 376859 674576 376871
rect 675472 376859 675478 376871
rect 674570 376831 675478 376859
rect 674570 376819 674576 376831
rect 675472 376819 675478 376831
rect 675530 376819 675536 376871
rect 674032 375709 674038 375761
rect 674090 375749 674096 375761
rect 675472 375749 675478 375761
rect 674090 375721 675478 375749
rect 674090 375709 674096 375721
rect 675472 375709 675478 375721
rect 675530 375709 675536 375761
rect 42160 375191 42166 375243
rect 42218 375231 42224 375243
rect 45424 375231 45430 375243
rect 42218 375203 45430 375231
rect 42218 375191 42224 375203
rect 45424 375191 45430 375203
rect 45482 375191 45488 375243
rect 37360 372527 37366 372579
rect 37418 372567 37424 372579
rect 42928 372567 42934 372579
rect 37418 372539 42934 372567
rect 37418 372527 37424 372539
rect 42928 372527 42934 372539
rect 42986 372527 42992 372579
rect 42064 370159 42070 370211
rect 42122 370159 42128 370211
rect 42256 370159 42262 370211
rect 42314 370199 42320 370211
rect 43312 370199 43318 370211
rect 42314 370171 43318 370199
rect 42314 370159 42320 370171
rect 43312 370159 43318 370171
rect 43370 370159 43376 370211
rect 42082 369829 42110 370159
rect 42160 369937 42166 369989
rect 42218 369977 42224 369989
rect 42352 369977 42358 369989
rect 42218 369949 42358 369977
rect 42218 369937 42224 369949
rect 42352 369937 42358 369949
rect 42410 369937 42416 369989
rect 42352 369829 42358 369841
rect 42082 369801 42358 369829
rect 42352 369789 42358 369801
rect 42410 369789 42416 369841
rect 50512 368679 50518 368731
rect 50570 368719 50576 368731
rect 59536 368719 59542 368731
rect 50570 368691 59542 368719
rect 50570 368679 50576 368691
rect 59536 368679 59542 368691
rect 59594 368679 59600 368731
rect 42064 368087 42070 368139
rect 42122 368127 42128 368139
rect 42352 368127 42358 368139
rect 42122 368099 42358 368127
rect 42122 368087 42128 368099
rect 42352 368087 42358 368099
rect 42410 368087 42416 368139
rect 42064 367347 42070 367399
rect 42122 367387 42128 367399
rect 50320 367387 50326 367399
rect 42122 367359 50326 367387
rect 42122 367347 42128 367359
rect 50320 367347 50326 367359
rect 50378 367347 50384 367399
rect 42064 366237 42070 366289
rect 42122 366277 42128 366289
rect 43024 366277 43030 366289
rect 42122 366249 43030 366277
rect 42122 366237 42128 366249
rect 43024 366237 43030 366249
rect 43082 366237 43088 366289
rect 43024 366089 43030 366141
rect 43082 366129 43088 366141
rect 43312 366129 43318 366141
rect 43082 366101 43318 366129
rect 43082 366089 43088 366101
rect 43312 366089 43318 366101
rect 43370 366089 43376 366141
rect 42160 364979 42166 365031
rect 42218 365019 42224 365031
rect 42736 365019 42742 365031
rect 42218 364991 42742 365019
rect 42218 364979 42224 364991
rect 42736 364979 42742 364991
rect 42794 364979 42800 365031
rect 42064 364239 42070 364291
rect 42122 364279 42128 364291
rect 42928 364279 42934 364291
rect 42122 364251 42934 364279
rect 42122 364239 42128 364251
rect 42928 364239 42934 364251
rect 42986 364239 42992 364291
rect 42352 364091 42358 364143
rect 42410 364131 42416 364143
rect 42832 364131 42838 364143
rect 42410 364103 42838 364131
rect 42410 364091 42416 364103
rect 42832 364091 42838 364103
rect 42890 364091 42896 364143
rect 661072 363869 661078 363921
rect 661130 363909 661136 363921
rect 674416 363909 674422 363921
rect 661130 363881 674422 363909
rect 661130 363869 661136 363881
rect 674416 363869 674422 363881
rect 674474 363869 674480 363921
rect 42160 363647 42166 363699
rect 42218 363687 42224 363699
rect 43120 363687 43126 363699
rect 42218 363659 43126 363687
rect 42218 363647 42224 363659
rect 43120 363647 43126 363659
rect 43178 363647 43184 363699
rect 654448 363351 654454 363403
rect 654506 363391 654512 363403
rect 661168 363391 661174 363403
rect 654506 363363 661174 363391
rect 654506 363351 654512 363363
rect 661168 363351 661174 363363
rect 661226 363351 661232 363403
rect 669808 363277 669814 363329
rect 669866 363317 669872 363329
rect 674608 363317 674614 363329
rect 669866 363289 674614 363317
rect 669866 363277 669872 363289
rect 674608 363277 674614 363289
rect 674666 363277 674672 363329
rect 655120 363055 655126 363107
rect 655178 363095 655184 363107
rect 674704 363095 674710 363107
rect 655178 363067 674710 363095
rect 655178 363055 655184 363067
rect 674704 363055 674710 363067
rect 674762 363055 674768 363107
rect 42256 362093 42262 362145
rect 42314 362133 42320 362145
rect 43024 362133 43030 362145
rect 42314 362105 43030 362133
rect 42314 362093 42320 362105
rect 43024 362093 43030 362105
rect 43082 362093 43088 362145
rect 42352 350697 42358 350749
rect 42410 350737 42416 350749
rect 53392 350737 53398 350749
rect 42410 350709 53398 350737
rect 42410 350697 42416 350709
rect 53392 350697 53398 350709
rect 53450 350697 53456 350749
rect 42640 349661 42646 349713
rect 42698 349701 42704 349713
rect 53488 349701 53494 349713
rect 42698 349673 53494 349701
rect 42698 349661 42704 349673
rect 53488 349661 53494 349673
rect 53546 349661 53552 349713
rect 42352 349069 42358 349121
rect 42410 349109 42416 349121
rect 45520 349109 45526 349121
rect 42410 349081 45526 349109
rect 42410 349069 42416 349081
rect 45520 349069 45526 349081
rect 45578 349069 45584 349121
rect 650320 345591 650326 345643
rect 650378 345631 650384 345643
rect 679792 345631 679798 345643
rect 650378 345603 679798 345631
rect 650378 345591 650384 345603
rect 679792 345591 679798 345603
rect 679850 345591 679856 345643
rect 674512 340929 674518 340981
rect 674570 340969 674576 340981
rect 675472 340969 675478 340981
rect 674570 340941 675478 340969
rect 674570 340929 674576 340941
rect 675472 340929 675478 340941
rect 675530 340929 675536 340981
rect 53296 339819 53302 339871
rect 53354 339859 53360 339871
rect 59536 339859 59542 339871
rect 53354 339831 59542 339859
rect 53354 339819 53360 339831
rect 59536 339819 59542 339831
rect 59594 339819 59600 339871
rect 654160 339819 654166 339871
rect 654218 339859 654224 339871
rect 666736 339859 666742 339871
rect 654218 339831 666742 339859
rect 654218 339819 654224 339831
rect 666736 339819 666742 339831
rect 666794 339819 666800 339871
rect 674032 339523 674038 339575
rect 674090 339563 674096 339575
rect 675376 339563 675382 339575
rect 674090 339535 675382 339563
rect 674090 339523 674096 339535
rect 675376 339523 675382 339535
rect 675434 339523 675440 339575
rect 674320 336563 674326 336615
rect 674378 336603 674384 336615
rect 675376 336603 675382 336615
rect 674378 336575 675382 336603
rect 674378 336563 674384 336575
rect 675376 336563 675382 336575
rect 675434 336563 675440 336615
rect 674896 336267 674902 336319
rect 674954 336307 674960 336319
rect 675088 336307 675094 336319
rect 674954 336279 675094 336307
rect 674954 336267 674960 336279
rect 675088 336267 675094 336279
rect 675146 336267 675152 336319
rect 674704 332715 674710 332767
rect 674762 332755 674768 332767
rect 675376 332755 675382 332767
rect 674762 332727 675382 332755
rect 674762 332715 674768 332727
rect 675376 332715 675382 332727
rect 675434 332715 675440 332767
rect 674224 332197 674230 332249
rect 674282 332237 674288 332249
rect 675472 332237 675478 332249
rect 674282 332209 675478 332237
rect 674282 332197 674288 332209
rect 675472 332197 675478 332209
rect 675530 332197 675536 332249
rect 42352 331975 42358 332027
rect 42410 332015 42416 332027
rect 45616 332015 45622 332027
rect 42410 331987 45622 332015
rect 42410 331975 42416 331987
rect 45616 331975 45622 331987
rect 45674 331975 45680 332027
rect 674992 331753 674998 331805
rect 675050 331793 675056 331805
rect 675376 331793 675382 331805
rect 675050 331765 675382 331793
rect 675050 331753 675056 331765
rect 675376 331753 675382 331765
rect 675434 331753 675440 331805
rect 653968 329755 653974 329807
rect 654026 329795 654032 329807
rect 663760 329795 663766 329807
rect 654026 329767 663766 329795
rect 654026 329755 654032 329767
rect 663760 329755 663766 329767
rect 663818 329755 663824 329807
rect 37264 329311 37270 329363
rect 37322 329351 37328 329363
rect 41776 329351 41782 329363
rect 37322 329323 41782 329351
rect 37322 329311 37328 329323
rect 41776 329311 41782 329323
rect 41834 329311 41840 329363
rect 37360 329163 37366 329215
rect 37418 329203 37424 329215
rect 41680 329203 41686 329215
rect 37418 329175 41686 329203
rect 37418 329163 37424 329175
rect 41680 329163 41686 329175
rect 41738 329163 41744 329215
rect 37168 328349 37174 328401
rect 37226 328389 37232 328401
rect 37226 328361 42494 328389
rect 37226 328349 37232 328361
rect 42466 328241 42494 328361
rect 43120 328275 43126 328327
rect 43178 328315 43184 328327
rect 43312 328315 43318 328327
rect 43178 328287 43318 328315
rect 43178 328275 43184 328287
rect 43312 328275 43318 328287
rect 43370 328275 43376 328327
rect 42466 328213 42974 328241
rect 42946 328093 42974 328213
rect 43024 328093 43030 328105
rect 42946 328065 43030 328093
rect 43024 328053 43030 328065
rect 43082 328053 43088 328105
rect 41680 327239 41686 327291
rect 41738 327279 41744 327291
rect 42352 327279 42358 327291
rect 41738 327251 42358 327279
rect 41738 327239 41744 327251
rect 42352 327239 42358 327251
rect 42410 327239 42416 327291
rect 41776 327017 41782 327069
rect 41834 327017 41840 327069
rect 41794 326773 41822 327017
rect 41776 326721 41782 326773
rect 41834 326721 41840 326773
rect 53392 325463 53398 325515
rect 53450 325503 53456 325515
rect 59536 325503 59542 325515
rect 53450 325475 59542 325503
rect 53450 325463 53456 325475
rect 59536 325463 59542 325475
rect 59594 325463 59600 325515
rect 42064 324871 42070 324923
rect 42122 324911 42128 324923
rect 42736 324911 42742 324923
rect 42122 324883 42742 324911
rect 42122 324871 42128 324883
rect 42736 324871 42742 324883
rect 42794 324871 42800 324923
rect 42160 324131 42166 324183
rect 42218 324171 42224 324183
rect 53200 324171 53206 324183
rect 42218 324143 53206 324171
rect 42218 324131 42224 324143
rect 53200 324131 53206 324143
rect 53258 324131 53264 324183
rect 42160 323095 42166 323147
rect 42218 323135 42224 323147
rect 43024 323135 43030 323147
rect 42218 323107 43030 323135
rect 42218 323095 42224 323107
rect 43024 323095 43030 323107
rect 43082 323095 43088 323147
rect 43024 322947 43030 322999
rect 43082 322987 43088 322999
rect 43312 322987 43318 322999
rect 43082 322959 43318 322987
rect 43082 322947 43088 322959
rect 43312 322947 43318 322959
rect 43370 322947 43376 322999
rect 42064 321763 42070 321815
rect 42122 321803 42128 321815
rect 43120 321803 43126 321815
rect 42122 321775 43126 321803
rect 42122 321763 42128 321775
rect 43120 321763 43126 321775
rect 43178 321763 43184 321815
rect 42160 321245 42166 321297
rect 42218 321285 42224 321297
rect 42352 321285 42358 321297
rect 42218 321257 42358 321285
rect 42218 321245 42224 321257
rect 42352 321245 42358 321257
rect 42410 321245 42416 321297
rect 42160 320579 42166 320631
rect 42218 320619 42224 320631
rect 43024 320619 43030 320631
rect 42218 320591 43030 320619
rect 42218 320579 42224 320591
rect 43024 320579 43030 320591
rect 43082 320579 43088 320631
rect 663856 319913 663862 319965
rect 663914 319953 663920 319965
rect 674704 319953 674710 319965
rect 663914 319925 674710 319953
rect 663914 319913 663920 319925
rect 674704 319913 674710 319925
rect 674762 319913 674768 319965
rect 666640 318877 666646 318929
rect 666698 318917 666704 318929
rect 674416 318917 674422 318929
rect 666698 318889 674422 318917
rect 666698 318877 666704 318889
rect 674416 318877 674422 318889
rect 674474 318877 674480 318929
rect 666928 318285 666934 318337
rect 666986 318325 666992 318337
rect 674704 318325 674710 318337
rect 666986 318297 674710 318325
rect 666986 318285 666992 318297
rect 674704 318285 674710 318297
rect 674762 318285 674768 318337
rect 42064 316879 42070 316931
rect 42122 316919 42128 316931
rect 43408 316919 43414 316931
rect 42122 316891 43414 316919
rect 42122 316879 42128 316891
rect 43408 316879 43414 316891
rect 43466 316879 43472 316931
rect 45520 311033 45526 311085
rect 45578 311073 45584 311085
rect 59536 311073 59542 311085
rect 45578 311045 59542 311073
rect 45578 311033 45584 311045
rect 59536 311033 59542 311045
rect 59594 311033 59600 311085
rect 42256 307481 42262 307533
rect 42314 307521 42320 307533
rect 45712 307521 45718 307533
rect 42314 307493 45718 307521
rect 42314 307481 42320 307493
rect 45712 307481 45718 307493
rect 45770 307481 45776 307533
rect 42256 306741 42262 306793
rect 42314 306781 42320 306793
rect 50512 306781 50518 306793
rect 42314 306753 50518 306781
rect 42314 306741 42320 306753
rect 50512 306741 50518 306753
rect 50570 306741 50576 306793
rect 42832 305483 42838 305535
rect 42890 305523 42896 305535
rect 59056 305523 59062 305535
rect 42890 305495 59062 305523
rect 42890 305483 42896 305495
rect 59056 305483 59062 305495
rect 59114 305483 59120 305535
rect 650416 299563 650422 299615
rect 650474 299603 650480 299615
rect 679792 299603 679798 299615
rect 650474 299575 679798 299603
rect 650474 299563 650480 299575
rect 679792 299563 679798 299575
rect 679850 299563 679856 299615
rect 674896 299489 674902 299541
rect 674954 299529 674960 299541
rect 676816 299529 676822 299541
rect 674954 299501 676822 299529
rect 674954 299489 674960 299501
rect 676816 299489 676822 299501
rect 676874 299489 676880 299541
rect 675184 299415 675190 299467
rect 675242 299455 675248 299467
rect 676912 299455 676918 299467
rect 675242 299427 676918 299455
rect 675242 299415 675248 299427
rect 676912 299415 676918 299427
rect 676970 299415 676976 299467
rect 675280 299341 675286 299393
rect 675338 299381 675344 299393
rect 677008 299381 677014 299393
rect 675338 299353 677014 299381
rect 675338 299341 675344 299353
rect 677008 299341 677014 299353
rect 677066 299341 677072 299393
rect 45712 296677 45718 296729
rect 45770 296717 45776 296729
rect 59536 296717 59542 296729
rect 45770 296689 59542 296717
rect 45770 296677 45776 296689
rect 59536 296677 59542 296689
rect 59594 296677 59600 296729
rect 674320 295937 674326 295989
rect 674378 295977 674384 295989
rect 675376 295977 675382 295989
rect 674378 295949 675382 295977
rect 674378 295937 674384 295949
rect 675376 295937 675382 295949
rect 675434 295937 675440 295989
rect 674608 295345 674614 295397
rect 674666 295385 674672 295397
rect 675472 295385 675478 295397
rect 674666 295357 675478 295385
rect 674666 295345 674672 295357
rect 675472 295345 675478 295357
rect 675530 295345 675536 295397
rect 674416 292681 674422 292733
rect 674474 292721 674480 292733
rect 675184 292721 675190 292733
rect 674474 292693 675190 292721
rect 674474 292681 674480 292693
rect 675184 292681 675190 292693
rect 675242 292681 675248 292733
rect 42640 289055 42646 289107
rect 42698 289095 42704 289107
rect 43216 289095 43222 289107
rect 42698 289067 43222 289095
rect 42698 289055 42704 289067
rect 43216 289055 43222 289067
rect 43274 289095 43280 289107
rect 45904 289095 45910 289107
rect 43274 289067 45910 289095
rect 43274 289055 43280 289067
rect 45904 289055 45910 289067
rect 45962 289055 45968 289107
rect 674896 288537 674902 288589
rect 674954 288577 674960 288589
rect 675472 288577 675478 288589
rect 674954 288549 675478 288577
rect 674954 288537 674960 288549
rect 675472 288537 675478 288549
rect 675530 288537 675536 288589
rect 39952 287945 39958 287997
rect 40010 287985 40016 287997
rect 42640 287985 42646 287997
rect 40010 287957 42646 287985
rect 40010 287945 40016 287957
rect 42640 287945 42646 287957
rect 42698 287945 42704 287997
rect 674032 287723 674038 287775
rect 674090 287763 674096 287775
rect 675376 287763 675382 287775
rect 674090 287735 675382 287763
rect 674090 287723 674096 287735
rect 675376 287723 675382 287735
rect 675434 287723 675440 287775
rect 673936 287205 673942 287257
rect 673994 287245 674000 287257
rect 675472 287245 675478 287257
rect 673994 287217 675478 287245
rect 673994 287205 674000 287217
rect 675472 287205 675478 287217
rect 675530 287205 675536 287257
rect 37360 286835 37366 286887
rect 37418 286875 37424 286887
rect 42736 286875 42742 286887
rect 37418 286847 42742 286875
rect 37418 286835 37424 286847
rect 42736 286835 42742 286847
rect 42794 286835 42800 286887
rect 674224 286761 674230 286813
rect 674282 286801 674288 286813
rect 675376 286801 675382 286813
rect 674282 286773 675382 286801
rect 674282 286761 674288 286773
rect 675376 286761 675382 286773
rect 675434 286761 675440 286813
rect 41776 283801 41782 283853
rect 41834 283801 41840 283853
rect 42160 283801 42166 283853
rect 42218 283841 42224 283853
rect 43312 283841 43318 283853
rect 42218 283813 43318 283841
rect 42218 283801 42224 283813
rect 43312 283801 43318 283813
rect 43370 283801 43376 283853
rect 41794 283409 41822 283801
rect 41776 283357 41782 283409
rect 41834 283357 41840 283409
rect 653776 282395 653782 282447
rect 653834 282435 653840 282447
rect 660880 282435 660886 282447
rect 653834 282407 660886 282435
rect 653834 282395 653840 282407
rect 660880 282395 660886 282407
rect 660938 282395 660944 282447
rect 45808 282247 45814 282299
rect 45866 282287 45872 282299
rect 57616 282287 57622 282299
rect 45866 282259 57622 282287
rect 45866 282247 45872 282259
rect 57616 282247 57622 282259
rect 57674 282247 57680 282299
rect 42160 281729 42166 281781
rect 42218 281769 42224 281781
rect 42640 281769 42646 281781
rect 42218 281741 42646 281769
rect 42218 281729 42224 281741
rect 42640 281729 42646 281741
rect 42698 281729 42704 281781
rect 42160 281063 42166 281115
rect 42218 281103 42224 281115
rect 47536 281103 47542 281115
rect 42218 281075 47542 281103
rect 42218 281063 42224 281075
rect 47536 281063 47542 281075
rect 47594 281063 47600 281115
rect 42160 279879 42166 279931
rect 42218 279919 42224 279931
rect 42736 279919 42742 279931
rect 42218 279891 42742 279919
rect 42218 279879 42224 279891
rect 42736 279879 42742 279891
rect 42794 279879 42800 279931
rect 42160 278547 42166 278599
rect 42218 278587 42224 278599
rect 42544 278587 42550 278599
rect 42218 278559 42550 278587
rect 42218 278547 42224 278559
rect 42544 278547 42550 278559
rect 42602 278547 42608 278599
rect 42160 277807 42166 277859
rect 42218 277847 42224 277859
rect 43120 277847 43126 277859
rect 42218 277819 43126 277847
rect 42218 277807 42224 277819
rect 43120 277807 43126 277819
rect 43178 277807 43184 277859
rect 43216 277807 43222 277859
rect 43274 277807 43280 277859
rect 43234 277637 43262 277807
rect 43216 277585 43222 277637
rect 43274 277585 43280 277637
rect 42064 277363 42070 277415
rect 42122 277403 42128 277415
rect 42832 277403 42838 277415
rect 42122 277375 42838 277403
rect 42122 277363 42128 277375
rect 42832 277363 42838 277375
rect 42890 277363 42896 277415
rect 64624 275143 64630 275195
rect 64682 275183 64688 275195
rect 67216 275183 67222 275195
rect 64682 275155 67222 275183
rect 64682 275143 64688 275155
rect 67216 275143 67222 275155
rect 67274 275143 67280 275195
rect 64720 275069 64726 275121
rect 64778 275109 64784 275121
rect 66832 275109 66838 275121
rect 64778 275081 66838 275109
rect 64778 275069 64784 275081
rect 66832 275069 66838 275081
rect 66890 275069 66896 275121
rect 512752 274995 512758 275047
rect 512810 275035 512816 275047
rect 649360 275035 649366 275047
rect 512810 275007 649366 275035
rect 512810 274995 512816 275007
rect 649360 274995 649366 275007
rect 649418 274995 649424 275047
rect 669712 274921 669718 274973
rect 669770 274961 669776 274973
rect 674704 274961 674710 274973
rect 669770 274933 674710 274961
rect 669770 274921 669776 274933
rect 674704 274921 674710 274933
rect 674762 274921 674768 274973
rect 522256 274551 522262 274603
rect 522314 274591 522320 274603
rect 522544 274591 522550 274603
rect 522314 274563 522550 274591
rect 522314 274551 522320 274563
rect 522544 274551 522550 274563
rect 522602 274551 522608 274603
rect 42256 274477 42262 274529
rect 42314 274517 42320 274529
rect 42736 274517 42742 274529
rect 42314 274489 42742 274517
rect 42314 274477 42320 274489
rect 42736 274477 42742 274489
rect 42794 274477 42800 274529
rect 660976 274033 660982 274085
rect 661034 274073 661040 274085
rect 674704 274073 674710 274085
rect 661034 274045 674710 274073
rect 661034 274033 661040 274045
rect 674704 274033 674710 274045
rect 674762 274033 674768 274085
rect 42256 273737 42262 273789
rect 42314 273777 42320 273789
rect 43120 273777 43126 273789
rect 42314 273749 43126 273777
rect 42314 273737 42320 273749
rect 43120 273737 43126 273749
rect 43178 273737 43184 273789
rect 282160 273737 282166 273789
rect 282218 273777 282224 273789
rect 299440 273777 299446 273789
rect 282218 273749 299446 273777
rect 282218 273737 282224 273749
rect 299440 273737 299446 273749
rect 299498 273737 299504 273789
rect 319696 273737 319702 273789
rect 319754 273777 319760 273789
rect 339760 273777 339766 273789
rect 319754 273749 339766 273777
rect 319754 273737 319760 273749
rect 339760 273737 339766 273749
rect 339818 273737 339824 273789
rect 403120 273515 403126 273567
rect 403178 273555 403184 273567
rect 410416 273555 410422 273567
rect 403178 273527 410422 273555
rect 403178 273515 403184 273527
rect 410416 273515 410422 273527
rect 410474 273515 410480 273567
rect 64816 273441 64822 273493
rect 64874 273481 64880 273493
rect 72592 273481 72598 273493
rect 64874 273453 72598 273481
rect 64874 273441 64880 273453
rect 72592 273441 72598 273453
rect 72650 273441 72656 273493
rect 437776 273441 437782 273493
rect 437834 273481 437840 273493
rect 443536 273481 443542 273493
rect 437834 273453 443542 273481
rect 437834 273441 437840 273453
rect 443536 273441 443542 273453
rect 443594 273441 443600 273493
rect 100912 273367 100918 273419
rect 100970 273407 100976 273419
rect 120784 273407 120790 273419
rect 100970 273379 120790 273407
rect 100970 273367 100976 273379
rect 120784 273367 120790 273379
rect 120842 273367 120848 273419
rect 207280 273367 207286 273419
rect 207338 273407 207344 273419
rect 208432 273407 208438 273419
rect 207338 273379 208438 273407
rect 207338 273367 207344 273379
rect 208432 273367 208438 273379
rect 208490 273367 208496 273419
rect 645136 273367 645142 273419
rect 645194 273407 645200 273419
rect 665200 273407 665206 273419
rect 645194 273379 665206 273407
rect 645194 273367 645200 273379
rect 665200 273367 665206 273379
rect 665258 273367 665264 273419
rect 256336 273293 256342 273345
rect 256394 273333 256400 273345
rect 276400 273333 276406 273345
rect 256394 273305 276406 273333
rect 256394 273293 256400 273305
rect 276400 273293 276406 273305
rect 276458 273293 276464 273345
rect 664048 273293 664054 273345
rect 664106 273333 664112 273345
rect 674704 273333 674710 273345
rect 664106 273305 674710 273333
rect 664106 273293 664112 273305
rect 674704 273293 674710 273305
rect 674762 273293 674768 273345
rect 66160 273219 66166 273271
rect 66218 273259 66224 273271
rect 80560 273259 80566 273271
rect 66218 273231 80566 273259
rect 66218 273219 66224 273231
rect 80560 273219 80566 273231
rect 80618 273219 80624 273271
rect 308464 272257 308470 272309
rect 308522 272297 308528 272309
rect 392656 272297 392662 272309
rect 308522 272269 392662 272297
rect 308522 272257 308528 272269
rect 392656 272257 392662 272269
rect 392714 272257 392720 272309
rect 297808 272183 297814 272235
rect 297866 272223 297872 272235
rect 391120 272223 391126 272235
rect 297866 272195 391126 272223
rect 297866 272183 297872 272195
rect 391120 272183 391126 272195
rect 391178 272183 391184 272235
rect 283504 272109 283510 272161
rect 283562 272149 283568 272161
rect 411952 272149 411958 272161
rect 283562 272121 411958 272149
rect 283562 272109 283568 272121
rect 411952 272109 411958 272121
rect 412010 272109 412016 272161
rect 64912 270925 64918 270977
rect 64970 270965 64976 270977
rect 67600 270965 67606 270977
rect 64970 270937 67606 270965
rect 64970 270925 64976 270937
rect 67600 270925 67606 270937
rect 67658 270925 67664 270977
rect 378448 270703 378454 270755
rect 378506 270743 378512 270755
rect 379504 270743 379510 270755
rect 378506 270715 379510 270743
rect 378506 270703 378512 270715
rect 379504 270703 379510 270715
rect 379562 270703 379568 270755
rect 67216 270629 67222 270681
rect 67274 270669 67280 270681
rect 72112 270669 72118 270681
rect 67274 270641 72118 270669
rect 67274 270629 67280 270641
rect 72112 270629 72118 270641
rect 72170 270629 72176 270681
rect 112240 270629 112246 270681
rect 112298 270669 112304 270681
rect 132976 270669 132982 270681
rect 112298 270641 132982 270669
rect 112298 270629 112304 270641
rect 132976 270629 132982 270641
rect 133034 270629 133040 270681
rect 137104 270629 137110 270681
rect 137162 270669 137168 270681
rect 140464 270669 140470 270681
rect 137162 270641 140470 270669
rect 137162 270629 137168 270641
rect 140464 270629 140470 270641
rect 140522 270629 140528 270681
rect 158608 270629 158614 270681
rect 158666 270669 158672 270681
rect 161200 270669 161206 270681
rect 158666 270641 161206 270669
rect 158666 270629 158672 270641
rect 161200 270629 161206 270641
rect 161258 270629 161264 270681
rect 162160 270629 162166 270681
rect 162218 270669 162224 270681
rect 164080 270669 164086 270681
rect 162218 270641 164086 270669
rect 162218 270629 162224 270641
rect 164080 270629 164086 270641
rect 164138 270629 164144 270681
rect 165808 270629 165814 270681
rect 165866 270669 165872 270681
rect 166960 270669 166966 270681
rect 165866 270641 166966 270669
rect 165866 270629 165872 270641
rect 166960 270629 166966 270641
rect 167018 270629 167024 270681
rect 172816 270629 172822 270681
rect 172874 270669 172880 270681
rect 175600 270669 175606 270681
rect 172874 270641 175606 270669
rect 172874 270629 172880 270641
rect 175600 270629 175606 270641
rect 175658 270629 175664 270681
rect 176464 270629 176470 270681
rect 176522 270669 176528 270681
rect 178480 270669 178486 270681
rect 176522 270641 178486 270669
rect 176522 270629 176528 270641
rect 178480 270629 178486 270641
rect 178538 270629 178544 270681
rect 180016 270629 180022 270681
rect 180074 270669 180080 270681
rect 181360 270669 181366 270681
rect 180074 270641 181366 270669
rect 180074 270629 180080 270641
rect 181360 270629 181366 270641
rect 181418 270629 181424 270681
rect 183472 270629 183478 270681
rect 183530 270669 183536 270681
rect 184240 270669 184246 270681
rect 183530 270641 184246 270669
rect 183530 270629 183536 270641
rect 184240 270629 184246 270641
rect 184298 270629 184304 270681
rect 184336 270629 184342 270681
rect 184394 270669 184400 270681
rect 426928 270669 426934 270681
rect 184394 270641 426934 270669
rect 184394 270629 184400 270641
rect 426928 270629 426934 270641
rect 426986 270629 426992 270681
rect 427888 270629 427894 270681
rect 427946 270669 427952 270681
rect 540400 270669 540406 270681
rect 427946 270641 540406 270669
rect 427946 270629 427952 270641
rect 540400 270629 540406 270641
rect 540458 270629 540464 270681
rect 72592 270555 72598 270607
rect 72650 270595 72656 270607
rect 80656 270595 80662 270607
rect 72650 270567 80662 270595
rect 72650 270555 72656 270567
rect 80656 270555 80662 270567
rect 80714 270555 80720 270607
rect 108592 270555 108598 270607
rect 108650 270595 108656 270607
rect 130000 270595 130006 270607
rect 108650 270567 130006 270595
rect 108650 270555 108656 270567
rect 130000 270555 130006 270567
rect 130058 270555 130064 270607
rect 130096 270555 130102 270607
rect 130154 270595 130160 270607
rect 139888 270595 139894 270607
rect 130154 270567 139894 270595
rect 130154 270555 130160 270567
rect 139888 270555 139894 270567
rect 139946 270555 139952 270607
rect 433072 270595 433078 270607
rect 178882 270567 433078 270595
rect 105040 270481 105046 270533
rect 105098 270521 105104 270533
rect 139312 270521 139318 270533
rect 105098 270493 139318 270521
rect 105098 270481 105104 270493
rect 139312 270481 139318 270493
rect 139370 270481 139376 270533
rect 174064 270481 174070 270533
rect 174122 270521 174128 270533
rect 178882 270521 178910 270567
rect 433072 270555 433078 270567
rect 433130 270555 433136 270607
rect 521968 270555 521974 270607
rect 522026 270595 522032 270607
rect 551056 270595 551062 270607
rect 522026 270567 551062 270595
rect 522026 270555 522032 270567
rect 551056 270555 551062 270567
rect 551114 270555 551120 270607
rect 174122 270493 178910 270521
rect 174122 270481 174128 270493
rect 179152 270481 179158 270533
rect 179210 270521 179216 270533
rect 440560 270521 440566 270533
rect 179210 270493 440566 270521
rect 179210 270481 179216 270493
rect 440560 270481 440566 270493
rect 440618 270481 440624 270533
rect 508336 270481 508342 270533
rect 508394 270521 508400 270533
rect 566512 270521 566518 270533
rect 508394 270493 566518 270521
rect 508394 270481 508400 270493
rect 566512 270481 566518 270493
rect 566570 270481 566576 270533
rect 101488 270407 101494 270459
rect 101546 270447 101552 270459
rect 139696 270447 139702 270459
rect 101546 270419 139702 270447
rect 101546 270407 101552 270419
rect 139696 270407 139702 270419
rect 139754 270407 139760 270459
rect 164560 270407 164566 270459
rect 164618 270447 164624 270459
rect 427984 270447 427990 270459
rect 164618 270419 427990 270447
rect 164618 270407 164624 270419
rect 427984 270407 427990 270419
rect 428042 270407 428048 270459
rect 429328 270407 429334 270459
rect 429386 270447 429392 270459
rect 429386 270419 432638 270447
rect 429386 270407 429392 270419
rect 97936 270333 97942 270385
rect 97994 270373 98000 270385
rect 132880 270373 132886 270385
rect 97994 270345 132886 270373
rect 97994 270333 98000 270345
rect 132880 270333 132886 270345
rect 132938 270333 132944 270385
rect 132976 270333 132982 270385
rect 133034 270373 133040 270385
rect 139120 270373 139126 270385
rect 133034 270345 139126 270373
rect 133034 270333 133040 270345
rect 139120 270333 139126 270345
rect 139178 270333 139184 270385
rect 159760 270333 159766 270385
rect 159818 270373 159824 270385
rect 424432 270373 424438 270385
rect 159818 270345 424438 270373
rect 159818 270333 159824 270345
rect 424432 270333 424438 270345
rect 424490 270333 424496 270385
rect 432304 270333 432310 270385
rect 432362 270373 432368 270385
rect 432610 270373 432638 270419
rect 432688 270407 432694 270459
rect 432746 270447 432752 270459
rect 564208 270447 564214 270459
rect 432746 270419 564214 270447
rect 432746 270407 432752 270419
rect 564208 270407 564214 270419
rect 564266 270407 564272 270459
rect 567664 270373 567670 270385
rect 432362 270345 432542 270373
rect 432610 270345 567670 270373
rect 432362 270333 432368 270345
rect 94384 270259 94390 270311
rect 94442 270299 94448 270311
rect 140176 270299 140182 270311
rect 94442 270271 140182 270299
rect 94442 270259 94448 270271
rect 140176 270259 140182 270271
rect 140234 270259 140240 270311
rect 163408 270259 163414 270311
rect 163466 270299 163472 270311
rect 432400 270299 432406 270311
rect 163466 270271 432406 270299
rect 163466 270259 163472 270271
rect 432400 270259 432406 270271
rect 432458 270259 432464 270311
rect 432514 270299 432542 270345
rect 567664 270333 567670 270345
rect 567722 270333 567728 270385
rect 577264 270299 577270 270311
rect 432514 270271 577270 270299
rect 577264 270259 577270 270271
rect 577322 270259 577328 270311
rect 89584 270185 89590 270237
rect 89642 270225 89648 270237
rect 139792 270225 139798 270237
rect 89642 270197 139798 270225
rect 89642 270185 89648 270197
rect 139792 270185 139798 270197
rect 139850 270185 139856 270237
rect 157360 270185 157366 270237
rect 157418 270225 157424 270237
rect 429232 270225 429238 270237
rect 157418 270197 429238 270225
rect 157418 270185 157424 270197
rect 429232 270185 429238 270197
rect 429290 270185 429296 270237
rect 432112 270185 432118 270237
rect 432170 270225 432176 270237
rect 580816 270225 580822 270237
rect 432170 270197 580822 270225
rect 432170 270185 432176 270197
rect 580816 270185 580822 270197
rect 580874 270185 580880 270237
rect 84784 270111 84790 270163
rect 84842 270151 84848 270163
rect 140368 270151 140374 270163
rect 84842 270123 140374 270151
rect 84842 270111 84848 270123
rect 140368 270111 140374 270123
rect 140426 270111 140432 270163
rect 152560 270111 152566 270163
rect 152618 270151 152624 270163
rect 424240 270151 424246 270163
rect 152618 270123 424246 270151
rect 152618 270111 152624 270123
rect 424240 270111 424246 270123
rect 424298 270111 424304 270163
rect 424816 270111 424822 270163
rect 424874 270151 424880 270163
rect 578416 270151 578422 270163
rect 424874 270123 578422 270151
rect 424874 270111 424880 270123
rect 578416 270111 578422 270123
rect 578474 270111 578480 270163
rect 80080 270037 80086 270089
rect 80138 270077 80144 270089
rect 139408 270077 139414 270089
rect 80138 270049 139414 270077
rect 80138 270037 80144 270049
rect 139408 270037 139414 270049
rect 139466 270037 139472 270089
rect 150256 270037 150262 270089
rect 150314 270077 150320 270089
rect 427312 270077 427318 270089
rect 150314 270049 427318 270077
rect 150314 270037 150320 270049
rect 427312 270037 427318 270049
rect 427370 270037 427376 270089
rect 427792 270037 427798 270089
rect 427850 270077 427856 270089
rect 582064 270077 582070 270089
rect 427850 270049 582070 270077
rect 427850 270037 427856 270049
rect 582064 270037 582070 270049
rect 582122 270037 582128 270089
rect 75280 269963 75286 270015
rect 75338 270003 75344 270015
rect 75338 269975 133406 270003
rect 75338 269963 75344 269975
rect 68176 269815 68182 269867
rect 68234 269855 68240 269867
rect 133264 269855 133270 269867
rect 68234 269827 133270 269855
rect 68234 269815 68240 269827
rect 133264 269815 133270 269827
rect 133322 269815 133328 269867
rect 133378 269855 133406 269975
rect 133552 269963 133558 270015
rect 133610 270003 133616 270015
rect 140272 270003 140278 270015
rect 133610 269975 140278 270003
rect 133610 269963 133616 269975
rect 140272 269963 140278 269975
rect 140330 269963 140336 270015
rect 146704 269963 146710 270015
rect 146762 270003 146768 270015
rect 426256 270003 426262 270015
rect 146762 269975 426262 270003
rect 146762 269963 146768 269975
rect 426256 269963 426262 269975
rect 426314 269963 426320 270015
rect 427120 269963 427126 270015
rect 427178 270003 427184 270015
rect 585520 270003 585526 270015
rect 427178 269975 585526 270003
rect 427178 269963 427184 269975
rect 585520 269963 585526 269975
rect 585578 269963 585584 270015
rect 139504 269889 139510 269941
rect 139562 269929 139568 269941
rect 425776 269929 425782 269941
rect 139562 269901 425782 269929
rect 139562 269889 139568 269901
rect 425776 269889 425782 269901
rect 425834 269889 425840 269941
rect 427216 269889 427222 269941
rect 427274 269929 427280 269941
rect 589168 269929 589174 269941
rect 427274 269901 589174 269929
rect 427274 269889 427280 269901
rect 589168 269889 589174 269901
rect 589226 269889 589232 269941
rect 140080 269855 140086 269867
rect 133378 269827 140086 269855
rect 140080 269815 140086 269827
rect 140138 269815 140144 269867
rect 141904 269815 141910 269867
rect 141962 269855 141968 269867
rect 429904 269855 429910 269867
rect 141962 269827 429910 269855
rect 141962 269815 141968 269827
rect 429904 269815 429910 269827
rect 429962 269815 429968 269867
rect 431152 269815 431158 269867
rect 431210 269855 431216 269867
rect 432688 269855 432694 269867
rect 431210 269827 432694 269855
rect 431210 269815 431216 269827
rect 432688 269815 432694 269827
rect 432746 269815 432752 269867
rect 434896 269815 434902 269867
rect 434954 269855 434960 269867
rect 598672 269855 598678 269867
rect 434954 269827 598678 269855
rect 434954 269815 434960 269827
rect 598672 269815 598678 269827
rect 598730 269815 598736 269867
rect 132496 269741 132502 269793
rect 132554 269781 132560 269793
rect 423184 269781 423190 269793
rect 132554 269753 423190 269781
rect 132554 269741 132560 269753
rect 423184 269741 423190 269753
rect 423242 269741 423248 269793
rect 429616 269741 429622 269793
rect 429674 269781 429680 269793
rect 596272 269781 596278 269793
rect 429674 269753 596278 269781
rect 429674 269741 429680 269753
rect 596272 269741 596278 269753
rect 596330 269741 596336 269793
rect 134800 269667 134806 269719
rect 134858 269707 134864 269719
rect 423472 269707 423478 269719
rect 134858 269679 423478 269707
rect 134858 269667 134864 269679
rect 423472 269667 423478 269679
rect 423530 269667 423536 269719
rect 429520 269667 429526 269719
rect 429578 269707 429584 269719
rect 599824 269707 599830 269719
rect 429578 269679 599830 269707
rect 429578 269667 429584 269679
rect 599824 269667 599830 269679
rect 599882 269667 599888 269719
rect 127696 269593 127702 269645
rect 127754 269633 127760 269645
rect 423376 269633 423382 269645
rect 127754 269605 423382 269633
rect 127754 269593 127760 269605
rect 423376 269593 423382 269605
rect 423434 269593 423440 269645
rect 426256 269593 426262 269645
rect 426314 269633 426320 269645
rect 428944 269633 428950 269645
rect 426314 269605 428950 269633
rect 426314 269593 426320 269605
rect 428944 269593 428950 269605
rect 429002 269593 429008 269645
rect 429712 269593 429718 269645
rect 429770 269633 429776 269645
rect 603376 269633 603382 269645
rect 429770 269605 603382 269633
rect 429770 269593 429776 269605
rect 603376 269593 603382 269605
rect 603434 269593 603440 269645
rect 121648 269519 121654 269571
rect 121706 269559 121712 269571
rect 425968 269559 425974 269571
rect 121706 269531 425974 269559
rect 121706 269519 121712 269531
rect 425968 269519 425974 269531
rect 426026 269519 426032 269571
rect 426832 269519 426838 269571
rect 426890 269559 426896 269571
rect 621232 269559 621238 269571
rect 426890 269531 621238 269559
rect 426890 269519 426896 269531
rect 621232 269519 621238 269531
rect 621290 269519 621296 269571
rect 128848 269445 128854 269497
rect 128906 269485 128912 269497
rect 440080 269485 440086 269497
rect 128906 269457 440086 269485
rect 128906 269445 128912 269457
rect 440080 269445 440086 269457
rect 440138 269445 440144 269497
rect 459088 269445 459094 269497
rect 459146 269485 459152 269497
rect 620080 269485 620086 269497
rect 459146 269457 620086 269485
rect 459146 269445 459152 269457
rect 620080 269445 620086 269457
rect 620138 269445 620144 269497
rect 114640 269371 114646 269423
rect 114698 269411 114704 269423
rect 427504 269411 427510 269423
rect 114698 269383 427510 269411
rect 114698 269371 114704 269383
rect 427504 269371 427510 269383
rect 427562 269371 427568 269423
rect 429424 269371 429430 269423
rect 429482 269411 429488 269423
rect 431152 269411 431158 269423
rect 429482 269383 431158 269411
rect 429482 269371 429488 269383
rect 431152 269371 431158 269383
rect 431210 269371 431216 269423
rect 432016 269371 432022 269423
rect 432074 269411 432080 269423
rect 605776 269411 605782 269423
rect 432074 269383 605782 269411
rect 432074 269371 432080 269383
rect 605776 269371 605782 269383
rect 605834 269371 605840 269423
rect 109840 269297 109846 269349
rect 109898 269337 109904 269349
rect 426448 269337 426454 269349
rect 109898 269309 426454 269337
rect 109898 269297 109904 269309
rect 426448 269297 426454 269309
rect 426506 269297 426512 269349
rect 429136 269297 429142 269349
rect 429194 269337 429200 269349
rect 616432 269337 616438 269349
rect 429194 269309 616438 269337
rect 429194 269297 429200 269309
rect 616432 269297 616438 269309
rect 616490 269297 616496 269349
rect 102640 269223 102646 269275
rect 102698 269263 102704 269275
rect 436816 269263 436822 269275
rect 102698 269235 436822 269263
rect 102698 269223 102704 269235
rect 436816 269223 436822 269235
rect 436874 269223 436880 269275
rect 452656 269223 452662 269275
rect 452714 269263 452720 269275
rect 648688 269263 648694 269275
rect 452714 269235 648694 269263
rect 452714 269223 452720 269235
rect 648688 269223 648694 269235
rect 648746 269223 648752 269275
rect 115792 269149 115798 269201
rect 115850 269189 115856 269201
rect 140560 269189 140566 269201
rect 115850 269161 140566 269189
rect 115850 269149 115856 269161
rect 140560 269149 140566 269161
rect 140618 269149 140624 269201
rect 166864 269149 166870 269201
rect 166922 269189 166928 269201
rect 421648 269189 421654 269201
rect 166922 269161 421654 269189
rect 166922 269149 166928 269161
rect 421648 269149 421654 269161
rect 421706 269149 421712 269201
rect 427696 269149 427702 269201
rect 427754 269189 427760 269201
rect 526096 269189 526102 269201
rect 427754 269161 526102 269189
rect 427754 269149 427760 269161
rect 526096 269149 526102 269161
rect 526154 269149 526160 269201
rect 119344 269075 119350 269127
rect 119402 269115 119408 269127
rect 140752 269115 140758 269127
rect 119402 269087 140758 269115
rect 119402 269075 119408 269087
rect 140752 269075 140758 269087
rect 140810 269075 140816 269127
rect 171664 269075 171670 269127
rect 171722 269115 171728 269127
rect 184336 269115 184342 269127
rect 171722 269087 184342 269115
rect 171722 269075 171728 269087
rect 184336 269075 184342 269087
rect 184394 269075 184400 269127
rect 184720 269075 184726 269127
rect 184778 269115 184784 269127
rect 184778 269087 419006 269115
rect 184778 269075 184784 269087
rect 133264 269001 133270 269053
rect 133322 269041 133328 269053
rect 140848 269041 140854 269053
rect 133322 269013 140854 269041
rect 133322 269001 133328 269013
rect 140848 269001 140854 269013
rect 140906 269001 140912 269053
rect 202576 269001 202582 269053
rect 202634 269041 202640 269053
rect 204304 269041 204310 269053
rect 202634 269013 204310 269041
rect 202634 269001 202640 269013
rect 204304 269001 204310 269013
rect 204362 269001 204368 269053
rect 418864 269041 418870 269053
rect 204418 269013 418870 269041
rect 126448 268927 126454 268979
rect 126506 268967 126512 268979
rect 140656 268967 140662 268979
rect 126506 268939 140662 268967
rect 126506 268927 126512 268939
rect 140656 268927 140662 268939
rect 140714 268927 140720 268979
rect 189520 268927 189526 268979
rect 189578 268967 189584 268979
rect 204418 268967 204446 269013
rect 418864 269001 418870 269013
rect 418922 269001 418928 269053
rect 418978 269041 419006 269087
rect 429040 269075 429046 269127
rect 429098 269115 429104 269127
rect 469360 269115 469366 269127
rect 429098 269087 469366 269115
rect 429098 269075 429104 269087
rect 469360 269075 469366 269087
rect 469418 269075 469424 269127
rect 480880 269075 480886 269127
rect 480938 269115 480944 269127
rect 489712 269115 489718 269127
rect 480938 269087 489718 269115
rect 480938 269075 480944 269087
rect 489712 269075 489718 269087
rect 489770 269075 489776 269127
rect 552208 269115 552214 269127
rect 532258 269087 552214 269115
rect 434608 269041 434614 269053
rect 418978 269013 434614 269041
rect 434608 269001 434614 269013
rect 434666 269001 434672 269053
rect 470800 269001 470806 269053
rect 470858 269041 470864 269053
rect 499696 269041 499702 269053
rect 470858 269013 499702 269041
rect 470858 269001 470864 269013
rect 499696 269001 499702 269013
rect 499754 269001 499760 269053
rect 509776 269001 509782 269053
rect 509834 269041 509840 269053
rect 532258 269041 532286 269087
rect 552208 269075 552214 269087
rect 552266 269075 552272 269127
rect 509834 269013 532286 269041
rect 509834 269001 509840 269013
rect 417616 268967 417622 268979
rect 189578 268939 204446 268967
rect 204514 268939 417622 268967
rect 189578 268927 189584 268939
rect 130000 268853 130006 268905
rect 130058 268893 130064 268905
rect 139600 268893 139606 268905
rect 130058 268865 139606 268893
rect 130058 268853 130064 268865
rect 139600 268853 139606 268865
rect 139658 268853 139664 268905
rect 132880 268779 132886 268831
rect 132938 268819 132944 268831
rect 140944 268819 140950 268831
rect 132938 268791 140950 268819
rect 132938 268779 132944 268791
rect 140944 268779 140950 268791
rect 141002 268779 141008 268831
rect 188272 268779 188278 268831
rect 188330 268819 188336 268831
rect 204514 268819 204542 268939
rect 417616 268927 417622 268939
rect 417674 268927 417680 268979
rect 418960 268927 418966 268979
rect 419018 268967 419024 268979
rect 429040 268967 429046 268979
rect 419018 268939 429046 268967
rect 419018 268927 419024 268939
rect 429040 268927 429046 268939
rect 429098 268927 429104 268979
rect 430000 268927 430006 268979
rect 430058 268967 430064 268979
rect 446416 268967 446422 268979
rect 430058 268939 446422 268967
rect 430058 268927 430064 268939
rect 446416 268927 446422 268939
rect 446474 268927 446480 268979
rect 446530 268939 459230 268967
rect 212176 268853 212182 268905
rect 212234 268893 212240 268905
rect 212944 268893 212950 268905
rect 212234 268865 212950 268893
rect 212234 268853 212240 268865
rect 212944 268853 212950 268865
rect 213002 268853 213008 268905
rect 219184 268853 219190 268905
rect 219242 268893 219248 268905
rect 221488 268893 221494 268905
rect 219242 268865 221494 268893
rect 219242 268853 219248 268865
rect 221488 268853 221494 268865
rect 221546 268853 221552 268905
rect 225232 268853 225238 268905
rect 225290 268893 225296 268905
rect 227344 268893 227350 268905
rect 225290 268865 227350 268893
rect 225290 268853 225296 268865
rect 227344 268853 227350 268865
rect 227402 268853 227408 268905
rect 389872 268893 389878 268905
rect 227458 268865 389878 268893
rect 188330 268791 204542 268819
rect 188330 268779 188336 268791
rect 210928 268779 210934 268831
rect 210986 268819 210992 268831
rect 213040 268819 213046 268831
rect 210986 268791 213046 268819
rect 210986 268779 210992 268791
rect 213040 268779 213046 268791
rect 213098 268779 213104 268831
rect 222832 268779 222838 268831
rect 222890 268819 222896 268831
rect 227458 268819 227486 268865
rect 389872 268853 389878 268865
rect 389930 268853 389936 268905
rect 389968 268853 389974 268905
rect 390026 268893 390032 268905
rect 391696 268893 391702 268905
rect 390026 268865 391702 268893
rect 390026 268853 390032 268865
rect 391696 268853 391702 268865
rect 391754 268853 391760 268905
rect 397648 268853 397654 268905
rect 397706 268893 397712 268905
rect 400720 268893 400726 268905
rect 397706 268865 400726 268893
rect 397706 268853 397712 268865
rect 400720 268853 400726 268865
rect 400778 268853 400784 268905
rect 401488 268853 401494 268905
rect 401546 268893 401552 268905
rect 408304 268893 408310 268905
rect 401546 268865 408310 268893
rect 401546 268853 401552 268865
rect 408304 268853 408310 268865
rect 408362 268853 408368 268905
rect 426544 268853 426550 268905
rect 426602 268893 426608 268905
rect 430192 268893 430198 268905
rect 426602 268865 430198 268893
rect 426602 268853 426608 268865
rect 430192 268853 430198 268865
rect 430250 268853 430256 268905
rect 446530 268893 446558 268939
rect 439138 268865 446558 268893
rect 222890 268791 227486 268819
rect 222890 268779 222896 268791
rect 227632 268779 227638 268831
rect 227690 268819 227696 268831
rect 230128 268819 230134 268831
rect 227690 268791 230134 268819
rect 227690 268779 227696 268791
rect 230128 268779 230134 268791
rect 230186 268779 230192 268831
rect 234640 268779 234646 268831
rect 234698 268819 234704 268831
rect 235888 268819 235894 268831
rect 234698 268791 235894 268819
rect 234698 268779 234704 268791
rect 235888 268779 235894 268791
rect 235946 268779 235952 268831
rect 252496 268779 252502 268831
rect 252554 268819 252560 268831
rect 253360 268819 253366 268831
rect 252554 268791 253366 268819
rect 252554 268779 252560 268791
rect 253360 268779 253366 268791
rect 253418 268779 253424 268831
rect 259696 268779 259702 268831
rect 259754 268819 259760 268831
rect 262000 268819 262006 268831
rect 259754 268791 262006 268819
rect 259754 268779 259760 268791
rect 262000 268779 262006 268791
rect 262058 268779 262064 268831
rect 266800 268779 266806 268831
rect 266858 268819 266864 268831
rect 267760 268819 267766 268831
rect 266858 268791 267766 268819
rect 266858 268779 266864 268791
rect 267760 268779 267766 268791
rect 267818 268779 267824 268831
rect 274000 268779 274006 268831
rect 274058 268819 274064 268831
rect 276400 268819 276406 268831
rect 274058 268791 276406 268819
rect 274058 268779 274064 268791
rect 276400 268779 276406 268791
rect 276458 268779 276464 268831
rect 298960 268779 298966 268831
rect 299018 268819 299024 268831
rect 300304 268819 300310 268831
rect 299018 268791 300310 268819
rect 299018 268779 299024 268791
rect 300304 268779 300310 268791
rect 300362 268779 300368 268831
rect 300400 268779 300406 268831
rect 300458 268819 300464 268831
rect 358480 268819 358486 268831
rect 300458 268791 358486 268819
rect 300458 268779 300464 268791
rect 358480 268779 358486 268791
rect 358538 268779 358544 268831
rect 364432 268779 364438 268831
rect 364490 268819 364496 268831
rect 366640 268819 366646 268831
rect 364490 268791 366646 268819
rect 364490 268779 364496 268791
rect 366640 268779 366646 268791
rect 366698 268779 366704 268831
rect 377488 268779 377494 268831
rect 377546 268819 377552 268831
rect 439138 268819 439166 268865
rect 377546 268791 439166 268819
rect 459202 268819 459230 268939
rect 460816 268927 460822 268979
rect 460874 268967 460880 268979
rect 509680 268967 509686 268979
rect 460874 268939 470942 268967
rect 460874 268927 460880 268939
rect 459280 268853 459286 268905
rect 459338 268893 459344 268905
rect 470800 268893 470806 268905
rect 459338 268865 470806 268893
rect 459338 268853 459344 268865
rect 470800 268853 470806 268865
rect 470858 268853 470864 268905
rect 470914 268893 470942 268939
rect 479554 268939 509686 268967
rect 479554 268893 479582 268939
rect 509680 268927 509686 268939
rect 509738 268927 509744 268979
rect 470914 268865 479582 268893
rect 489712 268853 489718 268905
rect 489770 268893 489776 268905
rect 533200 268893 533206 268905
rect 489770 268865 533206 268893
rect 489770 268853 489776 268865
rect 533200 268853 533206 268865
rect 533258 268853 533264 268905
rect 460816 268819 460822 268831
rect 459202 268791 460822 268819
rect 377546 268779 377552 268791
rect 460816 268779 460822 268791
rect 460874 268779 460880 268831
rect 122896 268705 122902 268757
rect 122954 268745 122960 268757
rect 139984 268745 139990 268757
rect 122954 268717 139990 268745
rect 122954 268705 122960 268717
rect 139984 268705 139990 268717
rect 140042 268705 140048 268757
rect 295408 268705 295414 268757
rect 295466 268745 295472 268757
rect 299536 268745 299542 268757
rect 295466 268717 299542 268745
rect 295466 268705 295472 268717
rect 299536 268705 299542 268717
rect 299594 268705 299600 268757
rect 300976 268705 300982 268757
rect 301034 268745 301040 268757
rect 306064 268745 306070 268757
rect 301034 268717 306070 268745
rect 301034 268705 301040 268717
rect 306064 268705 306070 268717
rect 306122 268705 306128 268757
rect 342064 268705 342070 268757
rect 342122 268745 342128 268757
rect 348784 268745 348790 268757
rect 342122 268717 348790 268745
rect 342122 268705 342128 268717
rect 348784 268705 348790 268717
rect 348842 268705 348848 268757
rect 364240 268705 364246 268757
rect 364298 268745 364304 268757
rect 370288 268745 370294 268757
rect 364298 268717 370294 268745
rect 364298 268705 364304 268717
rect 370288 268705 370294 268717
rect 370346 268705 370352 268757
rect 376240 268705 376246 268757
rect 376298 268745 376304 268757
rect 377200 268745 377206 268757
rect 376298 268717 377206 268745
rect 376298 268705 376304 268717
rect 377200 268705 377206 268717
rect 377258 268705 377264 268757
rect 378160 268705 378166 268757
rect 378218 268745 378224 268757
rect 393904 268745 393910 268757
rect 378218 268717 393910 268745
rect 378218 268705 378224 268717
rect 393904 268705 393910 268717
rect 393962 268705 393968 268757
rect 439120 268745 439126 268757
rect 394402 268717 439126 268745
rect 147952 268631 147958 268683
rect 148010 268671 148016 268683
rect 149680 268671 149686 268683
rect 148010 268643 149686 268671
rect 148010 268631 148016 268643
rect 149680 268631 149686 268643
rect 149738 268631 149744 268683
rect 226384 268631 226390 268683
rect 226442 268671 226448 268683
rect 227440 268671 227446 268683
rect 226442 268643 227446 268671
rect 226442 268631 226448 268643
rect 227440 268631 227446 268643
rect 227498 268631 227504 268683
rect 276304 268631 276310 268683
rect 276362 268671 276368 268683
rect 388720 268671 388726 268683
rect 276362 268643 388726 268671
rect 276362 268631 276368 268643
rect 388720 268631 388726 268643
rect 388778 268631 388784 268683
rect 190672 268557 190678 268609
rect 190730 268597 190736 268609
rect 192880 268597 192886 268609
rect 190730 268569 192886 268597
rect 190730 268557 190736 268569
rect 192880 268557 192886 268569
rect 192938 268557 192944 268609
rect 310672 268557 310678 268609
rect 310730 268597 310736 268609
rect 310730 268569 378782 268597
rect 310730 268557 310736 268569
rect 288208 268483 288214 268535
rect 288266 268523 288272 268535
rect 299152 268523 299158 268535
rect 288266 268495 299158 268523
rect 288266 268483 288272 268495
rect 299152 268483 299158 268495
rect 299210 268483 299216 268535
rect 307984 268523 307990 268535
rect 299362 268495 307990 268523
rect 283408 268409 283414 268461
rect 283466 268449 283472 268461
rect 288016 268449 288022 268461
rect 283466 268421 288022 268449
rect 283466 268409 283472 268421
rect 288016 268409 288022 268421
rect 288074 268409 288080 268461
rect 290608 268409 290614 268461
rect 290666 268449 290672 268461
rect 299362 268449 299390 268495
rect 307984 268483 307990 268495
rect 308042 268483 308048 268535
rect 308176 268483 308182 268535
rect 308234 268523 308240 268535
rect 378754 268523 378782 268569
rect 387280 268557 387286 268609
rect 387338 268597 387344 268609
rect 394402 268597 394430 268717
rect 439120 268705 439126 268717
rect 439178 268705 439184 268757
rect 439312 268705 439318 268757
rect 439370 268745 439376 268757
rect 548752 268745 548758 268757
rect 439370 268717 548758 268745
rect 439370 268705 439376 268717
rect 548752 268705 548758 268717
rect 548810 268705 548816 268757
rect 407728 268631 407734 268683
rect 407786 268671 407792 268683
rect 408976 268671 408982 268683
rect 407786 268643 408982 268671
rect 407786 268631 407792 268643
rect 408976 268631 408982 268643
rect 409034 268631 409040 268683
rect 417616 268631 417622 268683
rect 417674 268671 417680 268683
rect 426256 268671 426262 268683
rect 417674 268643 426262 268671
rect 417674 268631 417680 268643
rect 426256 268631 426262 268643
rect 426314 268631 426320 268683
rect 429040 268631 429046 268683
rect 429098 268671 429104 268683
rect 459280 268671 459286 268683
rect 429098 268643 459286 268671
rect 429098 268631 429104 268643
rect 459280 268631 459286 268643
rect 459338 268631 459344 268683
rect 387338 268569 394430 268597
rect 387338 268557 387344 268569
rect 408688 268557 408694 268609
rect 408746 268597 408752 268609
rect 508240 268597 508246 268609
rect 408746 268569 508246 268597
rect 408746 268557 408752 268569
rect 508240 268557 508246 268569
rect 508298 268557 508304 268609
rect 389680 268523 389686 268535
rect 308234 268495 378686 268523
rect 378754 268495 389686 268523
rect 308234 268483 308240 268495
rect 310672 268449 310678 268461
rect 290666 268421 299390 268449
rect 300514 268421 310678 268449
rect 290666 268409 290672 268421
rect 286192 268335 286198 268387
rect 286250 268375 286256 268387
rect 300400 268375 300406 268387
rect 286250 268347 300406 268375
rect 286250 268335 286256 268347
rect 300400 268335 300406 268347
rect 300458 268335 300464 268387
rect 281104 268261 281110 268313
rect 281162 268301 281168 268313
rect 298768 268301 298774 268313
rect 281162 268273 298774 268301
rect 281162 268261 281168 268273
rect 298768 268261 298774 268273
rect 298826 268261 298832 268313
rect 144304 268187 144310 268239
rect 144362 268227 144368 268239
rect 146512 268227 146518 268239
rect 144362 268199 146518 268227
rect 144362 268187 144368 268199
rect 146512 268187 146518 268199
rect 146570 268187 146576 268239
rect 288016 268187 288022 268239
rect 288074 268227 288080 268239
rect 300514 268227 300542 268421
rect 310672 268409 310678 268421
rect 310730 268409 310736 268461
rect 378658 268449 378686 268495
rect 389680 268483 389686 268495
rect 389738 268483 389744 268535
rect 390544 268483 390550 268535
rect 390602 268523 390608 268535
rect 400336 268523 400342 268535
rect 390602 268495 400342 268523
rect 390602 268483 390608 268495
rect 400336 268483 400342 268495
rect 400394 268483 400400 268535
rect 406576 268483 406582 268535
rect 406634 268523 406640 268535
rect 501136 268523 501142 268535
rect 406634 268495 501142 268523
rect 406634 268483 406640 268495
rect 501136 268483 501142 268495
rect 501194 268483 501200 268535
rect 390352 268449 390358 268461
rect 310786 268421 378590 268449
rect 378658 268421 390358 268449
rect 300592 268335 300598 268387
rect 300650 268375 300656 268387
rect 302416 268375 302422 268387
rect 300650 268347 302422 268375
rect 300650 268335 300656 268347
rect 302416 268335 302422 268347
rect 302474 268335 302480 268387
rect 304912 268261 304918 268313
rect 304970 268301 304976 268313
rect 310786 268301 310814 268421
rect 315664 268335 315670 268387
rect 315722 268375 315728 268387
rect 378562 268375 378590 268421
rect 390352 268409 390358 268421
rect 390410 268409 390416 268461
rect 391792 268409 391798 268461
rect 391850 268449 391856 268461
rect 403600 268449 403606 268461
rect 391850 268421 403606 268449
rect 391850 268409 391856 268421
rect 403600 268409 403606 268421
rect 403658 268409 403664 268461
rect 425680 268409 425686 268461
rect 425738 268449 425744 268461
rect 494032 268449 494038 268461
rect 425738 268421 494038 268449
rect 425738 268409 425744 268421
rect 494032 268409 494038 268421
rect 494090 268409 494096 268461
rect 499696 268409 499702 268461
rect 499754 268449 499760 268461
rect 518896 268449 518902 268461
rect 499754 268421 518902 268449
rect 499754 268409 499760 268421
rect 518896 268409 518902 268421
rect 518954 268409 518960 268461
rect 389008 268375 389014 268387
rect 315722 268347 378302 268375
rect 378562 268347 389014 268375
rect 315722 268335 315728 268347
rect 304970 268273 310814 268301
rect 304970 268261 304976 268273
rect 348400 268261 348406 268313
rect 348458 268301 348464 268313
rect 378160 268301 378166 268313
rect 348458 268273 378166 268301
rect 348458 268261 348464 268273
rect 378160 268261 378166 268273
rect 378218 268261 378224 268313
rect 378274 268301 378302 268347
rect 389008 268335 389014 268347
rect 389066 268335 389072 268387
rect 389872 268335 389878 268387
rect 389930 268375 389936 268387
rect 398800 268375 398806 268387
rect 389930 268347 398806 268375
rect 389930 268335 389936 268347
rect 398800 268335 398806 268347
rect 398858 268335 398864 268387
rect 408592 268335 408598 268387
rect 408650 268375 408656 268387
rect 418960 268375 418966 268387
rect 408650 268347 418966 268375
rect 408650 268335 408656 268347
rect 418960 268335 418966 268347
rect 419018 268335 419024 268387
rect 423280 268335 423286 268387
rect 423338 268375 423344 268387
rect 486832 268375 486838 268387
rect 423338 268347 486838 268375
rect 423338 268335 423344 268347
rect 486832 268335 486838 268347
rect 486890 268335 486896 268387
rect 393328 268301 393334 268313
rect 378274 268273 393334 268301
rect 393328 268261 393334 268273
rect 393386 268261 393392 268313
rect 424912 268261 424918 268313
rect 424970 268301 424976 268313
rect 479728 268301 479734 268313
rect 424970 268273 479734 268301
rect 424970 268261 424976 268273
rect 479728 268261 479734 268273
rect 479786 268261 479792 268313
rect 288074 268199 300542 268227
rect 288074 268187 288080 268199
rect 335824 268187 335830 268239
rect 335882 268227 335888 268239
rect 342064 268227 342070 268239
rect 335882 268199 342070 268227
rect 335882 268187 335888 268199
rect 342064 268187 342070 268199
rect 342122 268187 342128 268239
rect 378928 268227 378934 268239
rect 342178 268199 378934 268227
rect 301840 268113 301846 268165
rect 301898 268153 301904 268165
rect 316720 268153 316726 268165
rect 301898 268125 316726 268153
rect 301898 268113 301904 268125
rect 316720 268113 316726 268125
rect 316778 268113 316784 268165
rect 333424 268113 333430 268165
rect 333482 268153 333488 268165
rect 342178 268153 342206 268199
rect 378928 268187 378934 268199
rect 378986 268187 378992 268239
rect 388912 268187 388918 268239
rect 388970 268227 388976 268239
rect 396496 268227 396502 268239
rect 388970 268199 396502 268227
rect 388970 268187 388976 268199
rect 396496 268187 396502 268199
rect 396554 268187 396560 268239
rect 408976 268187 408982 268239
rect 409034 268227 409040 268239
rect 429040 268227 429046 268239
rect 409034 268199 429046 268227
rect 409034 268187 409040 268199
rect 429040 268187 429046 268199
rect 429098 268187 429104 268239
rect 476176 268227 476182 268239
rect 463522 268199 476182 268227
rect 333482 268125 342206 268153
rect 333482 268113 333488 268125
rect 368560 268113 368566 268165
rect 368618 268153 368624 268165
rect 376720 268153 376726 268165
rect 368618 268125 376726 268153
rect 368618 268113 368624 268125
rect 376720 268113 376726 268125
rect 376778 268113 376784 268165
rect 380176 268153 380182 268165
rect 376834 268125 380182 268153
rect 301744 268039 301750 268091
rect 301802 268079 301808 268091
rect 313264 268079 313270 268091
rect 301802 268051 313270 268079
rect 301802 268039 301808 268051
rect 313264 268039 313270 268051
rect 313322 268039 313328 268091
rect 332272 268039 332278 268091
rect 332330 268079 332336 268091
rect 348112 268079 348118 268091
rect 332330 268051 348118 268079
rect 332330 268039 332336 268051
rect 348112 268039 348118 268051
rect 348170 268039 348176 268091
rect 348208 268039 348214 268091
rect 348266 268079 348272 268091
rect 348266 268051 348542 268079
rect 348266 268039 348272 268051
rect 301360 267965 301366 268017
rect 301418 268005 301424 268017
rect 309616 268005 309622 268017
rect 301418 267977 309622 268005
rect 301418 267965 301424 267977
rect 309616 267965 309622 267977
rect 309674 267965 309680 268017
rect 328720 267965 328726 268017
rect 328778 268005 328784 268017
rect 328778 267977 339710 268005
rect 328778 267965 328784 267977
rect 151408 267891 151414 267943
rect 151466 267931 151472 267943
rect 152560 267931 152566 267943
rect 151466 267903 152566 267931
rect 151466 267891 151472 267903
rect 152560 267891 152566 267903
rect 152618 267891 152624 267943
rect 339682 267931 339710 267977
rect 339760 267965 339766 268017
rect 339818 268005 339824 268017
rect 348400 268005 348406 268017
rect 339818 267977 348406 268005
rect 339818 267965 339824 267977
rect 348400 267965 348406 267977
rect 348458 267965 348464 268017
rect 347536 267931 347542 267943
rect 339682 267903 347542 267931
rect 347536 267891 347542 267903
rect 347594 267891 347600 267943
rect 348514 267931 348542 268051
rect 358384 268039 358390 268091
rect 358442 268079 358448 268091
rect 376834 268079 376862 268125
rect 380176 268113 380182 268125
rect 380234 268113 380240 268165
rect 399568 268153 399574 268165
rect 383266 268125 399574 268153
rect 378448 268079 378454 268091
rect 358442 268051 376862 268079
rect 376930 268051 378454 268079
rect 358442 268039 358448 268051
rect 358480 267965 358486 268017
rect 358538 268005 358544 268017
rect 376930 268005 376958 268051
rect 378448 268039 378454 268051
rect 378506 268039 378512 268091
rect 383266 268079 383294 268125
rect 399568 268113 399574 268125
rect 399626 268113 399632 268165
rect 418864 268113 418870 268165
rect 418922 268153 418928 268165
rect 426544 268153 426550 268165
rect 418922 268125 426550 268153
rect 418922 268113 418928 268125
rect 426544 268113 426550 268125
rect 426602 268113 426608 268165
rect 440656 268113 440662 268165
rect 440714 268113 440720 268165
rect 463522 268153 463550 268199
rect 476176 268187 476182 268199
rect 476234 268187 476240 268239
rect 460738 268125 463550 268153
rect 378658 268051 383294 268079
rect 358538 267977 376958 268005
rect 358538 267965 358544 267977
rect 377200 267965 377206 268017
rect 377258 268005 377264 268017
rect 378658 268005 378686 268051
rect 383344 268039 383350 268091
rect 383402 268079 383408 268091
rect 399856 268079 399862 268091
rect 383402 268051 399862 268079
rect 383402 268039 383408 268051
rect 399856 268039 399862 268051
rect 399914 268039 399920 268091
rect 430480 268039 430486 268091
rect 430538 268079 430544 268091
rect 440674 268079 440702 268113
rect 430538 268051 440702 268079
rect 430538 268039 430544 268051
rect 377258 267977 378686 268005
rect 377258 267965 377264 267977
rect 378928 267965 378934 268017
rect 378986 268005 378992 268017
rect 395056 268005 395062 268017
rect 378986 267977 395062 268005
rect 378986 267965 378992 267977
rect 395056 267965 395062 267977
rect 395114 267965 395120 268017
rect 440656 267965 440662 268017
rect 440714 268005 440720 268017
rect 460738 268005 460766 268125
rect 440714 267977 460766 268005
rect 440714 267965 440720 267977
rect 368560 267931 368566 267943
rect 348514 267903 368566 267931
rect 368560 267891 368566 267903
rect 368618 267891 368624 267943
rect 394576 267931 394582 267943
rect 374530 267903 394582 267931
rect 326320 267817 326326 267869
rect 326378 267857 326384 267869
rect 328048 267857 328054 267869
rect 326378 267829 328054 267857
rect 326378 267817 326384 267829
rect 328048 267817 328054 267829
rect 328106 267817 328112 267869
rect 339568 267817 339574 267869
rect 339626 267857 339632 267869
rect 349264 267857 349270 267869
rect 339626 267829 349270 267857
rect 339626 267817 339632 267829
rect 349264 267817 349270 267829
rect 349322 267817 349328 267869
rect 365584 267817 365590 267869
rect 365642 267857 365648 267869
rect 374530 267857 374558 267903
rect 394576 267891 394582 267903
rect 394634 267891 394640 267943
rect 401872 267891 401878 267943
rect 401930 267931 401936 267943
rect 415504 267931 415510 267943
rect 401930 267903 415510 267931
rect 401930 267891 401936 267903
rect 415504 267891 415510 267903
rect 415562 267891 415568 267943
rect 521392 267891 521398 267943
rect 521450 267931 521456 267943
rect 522256 267931 522262 267943
rect 521450 267903 522262 267931
rect 521450 267891 521456 267903
rect 522256 267891 522262 267903
rect 522314 267891 522320 267943
rect 365642 267829 374558 267857
rect 365642 267817 365648 267829
rect 376720 267817 376726 267869
rect 376778 267857 376784 267869
rect 386992 267857 386998 267869
rect 376778 267829 386998 267857
rect 376778 267817 376784 267829
rect 386992 267817 386998 267829
rect 387050 267817 387056 267869
rect 508432 267817 508438 267869
rect 508490 267857 508496 267869
rect 512752 267857 512758 267869
rect 508490 267829 512758 267857
rect 508490 267817 508496 267829
rect 512752 267817 512758 267829
rect 512810 267817 512816 267869
rect 139216 267743 139222 267795
rect 139274 267783 139280 267795
rect 139696 267783 139702 267795
rect 139274 267755 139702 267783
rect 139274 267743 139280 267755
rect 139696 267743 139702 267755
rect 139754 267743 139760 267795
rect 247792 267743 247798 267795
rect 247850 267783 247856 267795
rect 372496 267783 372502 267795
rect 247850 267755 372502 267783
rect 247850 267743 247856 267755
rect 372496 267743 372502 267755
rect 372554 267743 372560 267795
rect 372592 267743 372598 267795
rect 372650 267783 372656 267795
rect 397744 267783 397750 267795
rect 372650 267755 397750 267783
rect 372650 267743 372656 267755
rect 397744 267743 397750 267755
rect 397802 267743 397808 267795
rect 402544 267743 402550 267795
rect 402602 267783 402608 267795
rect 429808 267783 429814 267795
rect 402602 267755 429814 267783
rect 402602 267743 402608 267755
rect 429808 267743 429814 267755
rect 429866 267743 429872 267795
rect 622096 267743 622102 267795
rect 622154 267783 622160 267795
rect 633136 267783 633142 267795
rect 622154 267755 633142 267783
rect 622154 267743 622160 267755
rect 633136 267743 633142 267755
rect 633194 267743 633200 267795
rect 244240 267669 244246 267721
rect 244298 267709 244304 267721
rect 378544 267709 378550 267721
rect 244298 267681 378550 267709
rect 244298 267669 244304 267681
rect 378544 267669 378550 267681
rect 378602 267669 378608 267721
rect 379984 267669 379990 267721
rect 380042 267709 380048 267721
rect 399376 267709 399382 267721
rect 380042 267681 399382 267709
rect 380042 267669 380048 267681
rect 399376 267669 399382 267681
rect 399434 267669 399440 267721
rect 402928 267669 402934 267721
rect 402986 267709 402992 267721
rect 436912 267709 436918 267721
rect 402986 267681 436918 267709
rect 402986 267669 402992 267681
rect 436912 267669 436918 267681
rect 436970 267669 436976 267721
rect 240688 267595 240694 267647
rect 240746 267635 240752 267647
rect 378352 267635 378358 267647
rect 240746 267607 378358 267635
rect 240746 267595 240752 267607
rect 378352 267595 378358 267607
rect 378410 267595 378416 267647
rect 378466 267607 378686 267635
rect 215728 267521 215734 267573
rect 215786 267561 215792 267573
rect 378466 267561 378494 267607
rect 215786 267533 378494 267561
rect 378658 267561 378686 267607
rect 378736 267595 378742 267647
rect 378794 267635 378800 267647
rect 397552 267635 397558 267647
rect 378794 267607 397558 267635
rect 378794 267595 378800 267607
rect 397552 267595 397558 267607
rect 397610 267595 397616 267647
rect 404080 267595 404086 267647
rect 404138 267635 404144 267647
rect 454672 267635 454678 267647
rect 404138 267607 454678 267635
rect 404138 267595 404144 267607
rect 454672 267595 454678 267607
rect 454730 267595 454736 267647
rect 403312 267561 403318 267573
rect 378658 267533 403318 267561
rect 215786 267521 215792 267533
rect 403312 267521 403318 267533
rect 403370 267521 403376 267573
rect 404368 267521 404374 267573
rect 404426 267561 404432 267573
rect 461872 267561 461878 267573
rect 404426 267533 461878 267561
rect 404426 267521 404432 267533
rect 461872 267521 461878 267533
rect 461930 267521 461936 267573
rect 208528 267447 208534 267499
rect 208586 267487 208592 267499
rect 379984 267487 379990 267499
rect 208586 267459 379990 267487
rect 208586 267447 208592 267459
rect 379984 267447 379990 267459
rect 380042 267447 380048 267499
rect 380080 267447 380086 267499
rect 380138 267487 380144 267499
rect 398992 267487 398998 267499
rect 380138 267459 398998 267487
rect 380138 267447 380144 267459
rect 398992 267447 398998 267459
rect 399050 267447 399056 267499
rect 404848 267447 404854 267499
rect 404906 267487 404912 267499
rect 468976 267487 468982 267499
rect 404906 267459 468982 267487
rect 404906 267447 404912 267459
rect 468976 267447 468982 267459
rect 469034 267447 469040 267499
rect 204976 267373 204982 267425
rect 205034 267413 205040 267425
rect 395536 267413 395542 267425
rect 205034 267385 395542 267413
rect 205034 267373 205040 267385
rect 395536 267373 395542 267385
rect 395594 267373 395600 267425
rect 399088 267413 399094 267425
rect 395650 267385 399094 267413
rect 354832 267299 354838 267351
rect 354890 267339 354896 267351
rect 372592 267339 372598 267351
rect 354890 267311 372598 267339
rect 354890 267299 354896 267311
rect 372592 267299 372598 267311
rect 372650 267299 372656 267351
rect 378832 267299 378838 267351
rect 378890 267339 378896 267351
rect 378890 267311 390782 267339
rect 378890 267299 378896 267311
rect 351280 267225 351286 267277
rect 351338 267265 351344 267277
rect 378736 267265 378742 267277
rect 351338 267237 378742 267265
rect 351338 267225 351344 267237
rect 378736 267225 378742 267237
rect 378794 267225 378800 267277
rect 379792 267225 379798 267277
rect 379850 267265 379856 267277
rect 379850 267237 382334 267265
rect 379850 267225 379856 267237
rect 336976 267151 336982 267203
rect 337034 267191 337040 267203
rect 339760 267191 339766 267203
rect 337034 267163 339766 267191
rect 337034 267151 337040 267163
rect 339760 267151 339766 267163
rect 339818 267151 339824 267203
rect 352912 267151 352918 267203
rect 352970 267191 352976 267203
rect 382192 267191 382198 267203
rect 352970 267163 382198 267191
rect 352970 267151 352976 267163
rect 382192 267151 382198 267163
rect 382250 267151 382256 267203
rect 382306 267191 382334 267237
rect 383152 267225 383158 267277
rect 383210 267265 383216 267277
rect 390640 267265 390646 267277
rect 383210 267237 390646 267265
rect 383210 267225 383216 267237
rect 390640 267225 390646 267237
rect 390698 267225 390704 267277
rect 390754 267265 390782 267311
rect 390832 267299 390838 267351
rect 390890 267339 390896 267351
rect 395650 267339 395678 267385
rect 399088 267373 399094 267385
rect 399146 267373 399152 267425
rect 402160 267373 402166 267425
rect 402218 267413 402224 267425
rect 422608 267413 422614 267425
rect 402218 267385 422614 267413
rect 402218 267373 402224 267385
rect 422608 267373 422614 267385
rect 422666 267373 422672 267425
rect 424432 267373 424438 267425
rect 424490 267413 424496 267425
rect 431632 267413 431638 267425
rect 424490 267385 431638 267413
rect 424490 267373 424496 267385
rect 431632 267373 431638 267385
rect 431690 267373 431696 267425
rect 547504 267413 547510 267425
rect 437410 267385 547510 267413
rect 390890 267311 395678 267339
rect 390890 267299 390896 267311
rect 397456 267299 397462 267351
rect 397514 267339 397520 267351
rect 399952 267339 399958 267351
rect 397514 267311 399958 267339
rect 397514 267299 397520 267311
rect 399952 267299 399958 267311
rect 400010 267299 400016 267351
rect 423664 267299 423670 267351
rect 423722 267339 423728 267351
rect 437410 267339 437438 267385
rect 547504 267373 547510 267385
rect 547562 267373 547568 267425
rect 423722 267311 437438 267339
rect 423722 267299 423728 267311
rect 480688 267299 480694 267351
rect 480746 267339 480752 267351
rect 489808 267339 489814 267351
rect 480746 267311 489814 267339
rect 480746 267299 480752 267311
rect 489808 267299 489814 267311
rect 489866 267299 489872 267351
rect 398416 267265 398422 267277
rect 390754 267237 398422 267265
rect 398416 267225 398422 267237
rect 398474 267225 398480 267277
rect 398800 267225 398806 267277
rect 398858 267265 398864 267277
rect 407344 267265 407350 267277
rect 398858 267237 407350 267265
rect 398858 267225 398864 267237
rect 407344 267225 407350 267237
rect 407402 267225 407408 267277
rect 535696 267225 535702 267277
rect 535754 267265 535760 267277
rect 536176 267265 536182 267277
rect 535754 267237 536182 267265
rect 535754 267225 535760 267237
rect 536176 267225 536182 267237
rect 536234 267225 536240 267277
rect 382306 267163 398942 267191
rect 256912 267077 256918 267129
rect 256970 267117 256976 267129
rect 277840 267117 277846 267129
rect 256970 267089 277846 267117
rect 256970 267077 256976 267089
rect 277840 267077 277846 267089
rect 277898 267077 277904 267129
rect 285616 267077 285622 267129
rect 285674 267117 285680 267129
rect 367888 267117 367894 267129
rect 285674 267089 367894 267117
rect 285674 267077 285680 267089
rect 367888 267077 367894 267089
rect 367946 267077 367952 267129
rect 372496 267077 372502 267129
rect 372554 267117 372560 267129
rect 372554 267089 381950 267117
rect 372554 267077 372560 267089
rect 182416 267003 182422 267055
rect 182474 267043 182480 267055
rect 277936 267043 277942 267055
rect 182474 267015 277942 267043
rect 182474 267003 182480 267015
rect 277936 267003 277942 267015
rect 277994 267003 278000 267055
rect 282832 267003 282838 267055
rect 282890 267043 282896 267055
rect 372688 267043 372694 267055
rect 282890 267015 372694 267043
rect 282890 267003 282896 267015
rect 372688 267003 372694 267015
rect 372746 267003 372752 267055
rect 381922 267043 381950 267089
rect 382000 267077 382006 267129
rect 382058 267117 382064 267129
rect 398800 267117 398806 267129
rect 382058 267089 398806 267117
rect 382058 267077 382064 267089
rect 398800 267077 398806 267089
rect 398858 267077 398864 267129
rect 382192 267043 382198 267055
rect 381922 267015 382198 267043
rect 382192 267003 382198 267015
rect 382250 267003 382256 267055
rect 382288 267003 382294 267055
rect 382346 267043 382352 267055
rect 393040 267043 393046 267055
rect 382346 267015 393046 267043
rect 382346 267003 382352 267015
rect 393040 267003 393046 267015
rect 393098 267003 393104 267055
rect 398914 267043 398942 267163
rect 399088 267151 399094 267203
rect 399146 267191 399152 267203
rect 600976 267191 600982 267203
rect 399146 267163 600982 267191
rect 399146 267151 399152 267163
rect 600976 267151 600982 267163
rect 601034 267151 601040 267203
rect 399184 267077 399190 267129
rect 399242 267117 399248 267129
rect 604624 267117 604630 267129
rect 399242 267089 604630 267117
rect 399242 267077 399248 267089
rect 604624 267077 604630 267089
rect 604682 267077 604688 267129
rect 610480 267077 610486 267129
rect 610538 267117 610544 267129
rect 621904 267117 621910 267129
rect 610538 267089 621910 267117
rect 610538 267077 610544 267089
rect 621904 267077 621910 267089
rect 621962 267077 621968 267129
rect 608176 267043 608182 267055
rect 398914 267015 608182 267043
rect 608176 267003 608182 267015
rect 608234 267003 608240 267055
rect 610288 267003 610294 267055
rect 610346 267043 610352 267055
rect 612016 267043 612022 267055
rect 610346 267015 612022 267043
rect 610346 267003 610352 267015
rect 612016 267003 612022 267015
rect 612074 267003 612080 267055
rect 235984 266929 235990 266981
rect 236042 266969 236048 266981
rect 337360 266969 337366 266981
rect 236042 266941 337366 266969
rect 236042 266929 236048 266941
rect 337360 266929 337366 266941
rect 337418 266929 337424 266981
rect 348496 266929 348502 266981
rect 348554 266969 348560 266981
rect 368560 266969 368566 266981
rect 348554 266941 368566 266969
rect 348554 266929 348560 266941
rect 368560 266929 368566 266941
rect 368618 266929 368624 266981
rect 378544 266929 378550 266981
rect 378602 266969 378608 266981
rect 382576 266969 382582 266981
rect 378602 266941 382582 266969
rect 378602 266929 378608 266941
rect 382576 266929 382582 266941
rect 382634 266929 382640 266981
rect 382672 266929 382678 266981
rect 382730 266969 382736 266981
rect 382730 266941 393086 266969
rect 382730 266929 382736 266941
rect 221584 266855 221590 266907
rect 221642 266895 221648 266907
rect 360208 266895 360214 266907
rect 221642 266867 360214 266895
rect 221642 266855 221648 266867
rect 360208 266855 360214 266867
rect 360266 266855 360272 266907
rect 362032 266855 362038 266907
rect 362090 266895 362096 266907
rect 378832 266895 378838 266907
rect 362090 266867 378838 266895
rect 362090 266855 362096 266867
rect 378832 266855 378838 266867
rect 378890 266855 378896 266907
rect 387856 266895 387862 266907
rect 379138 266867 387862 266895
rect 72112 266781 72118 266833
rect 72170 266821 72176 266833
rect 83632 266821 83638 266833
rect 72170 266793 83638 266821
rect 72170 266781 72176 266793
rect 83632 266781 83638 266793
rect 83690 266781 83696 266833
rect 233488 266781 233494 266833
rect 233546 266821 233552 266833
rect 256912 266821 256918 266833
rect 233546 266793 256918 266821
rect 233546 266781 233552 266793
rect 256912 266781 256918 266793
rect 256970 266781 256976 266833
rect 277840 266781 277846 266833
rect 277898 266821 277904 266833
rect 277898 266793 378686 266821
rect 277898 266781 277904 266793
rect 229936 266707 229942 266759
rect 229994 266747 230000 266759
rect 377200 266747 377206 266759
rect 229994 266719 377206 266747
rect 229994 266707 230000 266719
rect 377200 266707 377206 266719
rect 377258 266707 377264 266759
rect 378658 266747 378686 266793
rect 378736 266781 378742 266833
rect 378794 266821 378800 266833
rect 379138 266821 379166 266867
rect 387856 266855 387862 266867
rect 387914 266855 387920 266907
rect 393058 266895 393086 266941
rect 398992 266929 398998 266981
rect 399050 266969 399056 266981
rect 498256 266969 498262 266981
rect 399050 266941 498262 266969
rect 399050 266929 399056 266941
rect 498256 266929 498262 266941
rect 498314 266929 498320 266981
rect 498352 266929 498358 266981
rect 498410 266929 498416 266981
rect 498544 266929 498550 266981
rect 498602 266969 498608 266981
rect 611728 266969 611734 266981
rect 498602 266941 611734 266969
rect 498602 266929 498608 266941
rect 611728 266929 611734 266941
rect 611786 266929 611792 266981
rect 418960 266895 418966 266907
rect 393058 266867 418966 266895
rect 418960 266855 418966 266867
rect 419018 266855 419024 266907
rect 460816 266855 460822 266907
rect 460874 266895 460880 266907
rect 485200 266895 485206 266907
rect 460874 266867 485206 266895
rect 460874 266855 460880 266867
rect 485200 266855 485206 266867
rect 485258 266855 485264 266907
rect 495280 266855 495286 266907
rect 495338 266895 495344 266907
rect 498370 266895 498398 266929
rect 495338 266867 498398 266895
rect 495338 266855 495344 266867
rect 570256 266855 570262 266907
rect 570314 266895 570320 266907
rect 610480 266895 610486 266907
rect 570314 266867 610486 266895
rect 570314 266855 570320 266867
rect 610480 266855 610486 266867
rect 610538 266855 610544 266907
rect 378794 266793 379166 266821
rect 378794 266781 378800 266793
rect 379216 266781 379222 266833
rect 379274 266821 379280 266833
rect 398512 266821 398518 266833
rect 379274 266793 398518 266821
rect 379274 266781 379280 266793
rect 398512 266781 398518 266793
rect 398570 266781 398576 266833
rect 398800 266781 398806 266833
rect 398858 266821 398864 266833
rect 480688 266821 480694 266833
rect 398858 266793 480694 266821
rect 398858 266781 398864 266793
rect 480688 266781 480694 266793
rect 480746 266781 480752 266833
rect 489808 266781 489814 266833
rect 489866 266821 489872 266833
rect 535504 266821 535510 266833
rect 489866 266793 535510 266821
rect 489866 266781 489872 266793
rect 535504 266781 535510 266793
rect 535562 266781 535568 266833
rect 535600 266781 535606 266833
rect 535658 266821 535664 266833
rect 590224 266821 590230 266833
rect 535658 266793 590230 266821
rect 535658 266781 535664 266793
rect 590224 266781 590230 266793
rect 590282 266781 590288 266833
rect 590512 266781 590518 266833
rect 590570 266821 590576 266833
rect 610384 266821 610390 266833
rect 590570 266793 610390 266821
rect 590570 266781 590576 266793
rect 610384 266781 610390 266793
rect 610442 266781 610448 266833
rect 610672 266781 610678 266833
rect 610730 266821 610736 266833
rect 626032 266821 626038 266833
rect 610730 266793 626038 266821
rect 610730 266781 610736 266793
rect 626032 266781 626038 266793
rect 626090 266781 626096 266833
rect 381232 266747 381238 266759
rect 378658 266719 381238 266747
rect 381232 266707 381238 266719
rect 381290 266707 381296 266759
rect 382576 266707 382582 266759
rect 382634 266747 382640 266759
rect 383632 266747 383638 266759
rect 382634 266719 383638 266747
rect 382634 266707 382640 266719
rect 383632 266707 383638 266719
rect 383690 266707 383696 266759
rect 383728 266707 383734 266759
rect 383786 266747 383792 266759
rect 386320 266747 386326 266759
rect 383786 266719 386326 266747
rect 383786 266707 383792 266719
rect 386320 266707 386326 266719
rect 386378 266707 386384 266759
rect 393040 266707 393046 266759
rect 393098 266747 393104 266759
rect 480784 266747 480790 266759
rect 393098 266719 480790 266747
rect 393098 266707 393104 266719
rect 480784 266707 480790 266719
rect 480842 266707 480848 266759
rect 489712 266707 489718 266759
rect 489770 266747 489776 266759
rect 590128 266747 590134 266759
rect 489770 266719 590134 266747
rect 489770 266707 489776 266719
rect 590128 266707 590134 266719
rect 590186 266707 590192 266759
rect 590608 266707 590614 266759
rect 590666 266747 590672 266759
rect 610288 266747 610294 266759
rect 590666 266719 610294 266747
rect 590666 266707 590672 266719
rect 610288 266707 610294 266719
rect 610346 266707 610352 266759
rect 612016 266707 612022 266759
rect 612074 266747 612080 266759
rect 629584 266747 629590 266759
rect 612074 266719 629590 266747
rect 612074 266707 612080 266719
rect 629584 266707 629590 266719
rect 629642 266707 629648 266759
rect 66832 266633 66838 266685
rect 66890 266673 66896 266685
rect 80560 266673 80566 266685
rect 66890 266645 80566 266673
rect 66890 266633 66896 266645
rect 80560 266633 80566 266645
rect 80618 266633 80624 266685
rect 135952 266633 135958 266685
rect 136010 266673 136016 266685
rect 282256 266673 282262 266685
rect 136010 266645 282262 266673
rect 136010 266633 136016 266645
rect 282256 266633 282262 266645
rect 282314 266633 282320 266685
rect 289264 266633 289270 266685
rect 289322 266673 289328 266685
rect 377488 266673 377494 266685
rect 289322 266645 377494 266673
rect 289322 266633 289328 266645
rect 377488 266633 377494 266645
rect 377546 266633 377552 266685
rect 378544 266633 378550 266685
rect 378602 266673 378608 266685
rect 386704 266673 386710 266685
rect 378602 266645 386710 266673
rect 378602 266633 378608 266645
rect 386704 266633 386710 266645
rect 386762 266633 386768 266685
rect 418960 266633 418966 266685
rect 419018 266673 419024 266685
rect 460816 266673 460822 266685
rect 419018 266645 460822 266673
rect 419018 266633 419024 266645
rect 460816 266633 460822 266645
rect 460874 266633 460880 266685
rect 535504 266633 535510 266685
rect 535562 266673 535568 266685
rect 538480 266673 538486 266685
rect 535562 266645 538486 266673
rect 535562 266633 535568 266645
rect 538480 266633 538486 266645
rect 538538 266633 538544 266685
rect 561520 266633 561526 266685
rect 561578 266673 561584 266685
rect 570256 266673 570262 266685
rect 561578 266645 570262 266673
rect 561578 266633 561584 266645
rect 570256 266633 570262 266645
rect 570314 266633 570320 266685
rect 125296 266559 125302 266611
rect 125354 266599 125360 266611
rect 277840 266599 277846 266611
rect 125354 266571 277846 266599
rect 125354 266559 125360 266571
rect 277840 266559 277846 266571
rect 277898 266559 277904 266611
rect 286576 266559 286582 266611
rect 286634 266599 286640 266611
rect 378640 266599 378646 266611
rect 286634 266571 378646 266599
rect 286634 266559 286640 266571
rect 378640 266559 378646 266571
rect 378698 266559 378704 266611
rect 378832 266559 378838 266611
rect 378890 266599 378896 266611
rect 397456 266599 397462 266611
rect 378890 266571 397462 266599
rect 378890 266559 378896 266571
rect 397456 266559 397462 266571
rect 397514 266559 397520 266611
rect 397648 266559 397654 266611
rect 397706 266599 397712 266611
rect 535792 266599 535798 266611
rect 397706 266571 535798 266599
rect 397706 266559 397712 266571
rect 535792 266559 535798 266571
rect 535850 266559 535856 266611
rect 535984 266559 535990 266611
rect 536042 266599 536048 266611
rect 636688 266599 636694 266611
rect 536042 266571 636694 266599
rect 536042 266559 536048 266571
rect 636688 266559 636694 266571
rect 636746 266559 636752 266611
rect 194320 266485 194326 266537
rect 194378 266525 194384 266537
rect 373072 266525 373078 266537
rect 194378 266497 373078 266525
rect 194378 266485 194384 266497
rect 373072 266485 373078 266497
rect 373130 266485 373136 266537
rect 374800 266485 374806 266537
rect 374858 266525 374864 266537
rect 383440 266525 383446 266537
rect 374858 266497 383446 266525
rect 374858 266485 374864 266497
rect 383440 266485 383446 266497
rect 383498 266485 383504 266537
rect 385744 266525 385750 266537
rect 383554 266497 385750 266525
rect 201328 266411 201334 266463
rect 201386 266451 201392 266463
rect 378064 266451 378070 266463
rect 201386 266423 378070 266451
rect 201386 266411 201392 266423
rect 378064 266411 378070 266423
rect 378122 266411 378128 266463
rect 378160 266411 378166 266463
rect 378218 266451 378224 266463
rect 383344 266451 383350 266463
rect 378218 266423 383350 266451
rect 378218 266411 378224 266423
rect 383344 266411 383350 266423
rect 383402 266411 383408 266463
rect 383554 266451 383582 266497
rect 385744 266485 385750 266497
rect 385802 266485 385808 266537
rect 393424 266485 393430 266537
rect 393482 266525 393488 266537
rect 535696 266525 535702 266537
rect 393482 266497 535702 266525
rect 393482 266485 393488 266497
rect 535696 266485 535702 266497
rect 535754 266485 535760 266537
rect 545680 266485 545686 266537
rect 545738 266525 545744 266537
rect 640240 266525 640246 266537
rect 545738 266497 640246 266525
rect 545738 266485 545744 266497
rect 640240 266485 640246 266497
rect 640298 266485 640304 266537
rect 383458 266423 383582 266451
rect 82480 266337 82486 266389
rect 82538 266377 82544 266389
rect 282544 266377 282550 266389
rect 82538 266349 282550 266377
rect 82538 266337 82544 266349
rect 282544 266337 282550 266349
rect 282602 266337 282608 266389
rect 282640 266337 282646 266389
rect 282698 266377 282704 266389
rect 383458 266377 383486 266423
rect 383824 266411 383830 266463
rect 383882 266451 383888 266463
rect 643888 266451 643894 266463
rect 383882 266423 643894 266451
rect 383882 266411 383888 266423
rect 643888 266411 643894 266423
rect 643946 266411 643952 266463
rect 282698 266349 383486 266377
rect 282698 266337 282704 266349
rect 383536 266337 383542 266389
rect 383594 266377 383600 266389
rect 393424 266377 393430 266389
rect 383594 266349 393430 266377
rect 383594 266337 383600 266349
rect 393424 266337 393430 266349
rect 393482 266337 393488 266389
rect 398800 266337 398806 266389
rect 398858 266377 398864 266389
rect 647440 266377 647446 266389
rect 398858 266349 647446 266377
rect 398858 266337 398864 266349
rect 647440 266337 647446 266349
rect 647498 266337 647504 266389
rect 254896 266263 254902 266315
rect 254954 266303 254960 266315
rect 374800 266303 374806 266315
rect 254954 266275 374806 266303
rect 254954 266263 254960 266275
rect 374800 266263 374806 266275
rect 374858 266263 374864 266315
rect 374896 266263 374902 266315
rect 374954 266303 374960 266315
rect 394864 266303 394870 266315
rect 374954 266275 394870 266303
rect 374954 266263 374960 266275
rect 394864 266263 394870 266275
rect 394922 266263 394928 266315
rect 408112 266263 408118 266315
rect 408170 266303 408176 266315
rect 427696 266303 427702 266315
rect 408170 266275 427702 266303
rect 408170 266263 408176 266275
rect 427696 266263 427702 266275
rect 427754 266263 427760 266315
rect 480784 266263 480790 266315
rect 480842 266303 480848 266315
rect 489712 266303 489718 266315
rect 480842 266275 489718 266303
rect 480842 266263 480848 266275
rect 489712 266263 489718 266275
rect 489770 266263 489776 266315
rect 498448 266263 498454 266315
rect 498506 266303 498512 266315
rect 535408 266303 535414 266315
rect 498506 266275 535414 266303
rect 498506 266263 498512 266275
rect 535408 266263 535414 266275
rect 535466 266263 535472 266315
rect 541744 266263 541750 266315
rect 541802 266303 541808 266315
rect 542800 266303 542806 266315
rect 541802 266275 542806 266303
rect 541802 266263 541808 266275
rect 542800 266263 542806 266275
rect 542858 266263 542864 266315
rect 258544 266189 258550 266241
rect 258602 266229 258608 266241
rect 378544 266229 378550 266241
rect 258602 266201 378550 266229
rect 258602 266189 258608 266201
rect 378544 266189 378550 266201
rect 378602 266189 378608 266241
rect 378754 266201 378974 266229
rect 262096 266115 262102 266167
rect 262154 266155 262160 266167
rect 378754 266155 378782 266201
rect 262154 266127 378782 266155
rect 262154 266115 262160 266127
rect 287920 266041 287926 266093
rect 287978 266081 287984 266093
rect 378736 266081 378742 266093
rect 287978 266053 378742 266081
rect 287978 266041 287984 266053
rect 378736 266041 378742 266053
rect 378794 266041 378800 266093
rect 272752 265967 272758 266019
rect 272810 266007 272816 266019
rect 348496 266007 348502 266019
rect 272810 265979 348502 266007
rect 272810 265967 272816 265979
rect 348496 265967 348502 265979
rect 348554 265967 348560 266019
rect 368560 265967 368566 266019
rect 368618 266007 368624 266019
rect 378160 266007 378166 266019
rect 368618 265979 378166 266007
rect 368618 265967 368624 265979
rect 378160 265967 378166 265979
rect 378218 265967 378224 266019
rect 378832 265967 378838 266019
rect 378890 265967 378896 266019
rect 286864 265893 286870 265945
rect 286922 265933 286928 265945
rect 378850 265933 378878 265967
rect 286922 265905 378878 265933
rect 378946 265933 378974 266201
rect 379408 266189 379414 266241
rect 379466 266229 379472 266241
rect 399184 266229 399190 266241
rect 379466 266201 399190 266229
rect 379466 266189 379472 266201
rect 399184 266189 399190 266201
rect 399242 266189 399248 266241
rect 405136 266189 405142 266241
rect 405194 266229 405200 266241
rect 430480 266229 430486 266241
rect 405194 266201 430486 266229
rect 405194 266189 405200 266201
rect 430480 266189 430486 266201
rect 430538 266189 430544 266241
rect 485200 266189 485206 266241
rect 485258 266229 485264 266241
rect 495280 266229 495286 266241
rect 485258 266201 495286 266229
rect 485258 266189 485264 266201
rect 495280 266189 495286 266201
rect 495338 266189 495344 266241
rect 535696 266189 535702 266241
rect 535754 266229 535760 266241
rect 545680 266229 545686 266241
rect 535754 266201 545686 266229
rect 535754 266189 535760 266201
rect 545680 266189 545686 266201
rect 545738 266189 545744 266241
rect 379024 266115 379030 266167
rect 379082 266155 379088 266167
rect 383152 266155 383158 266167
rect 379082 266127 383158 266155
rect 379082 266115 379088 266127
rect 383152 266115 383158 266127
rect 383210 266115 383216 266167
rect 383344 266115 383350 266167
rect 383402 266155 383408 266167
rect 388528 266155 388534 266167
rect 383402 266127 388534 266155
rect 383402 266115 383408 266127
rect 388528 266115 388534 266127
rect 388586 266115 388592 266167
rect 389008 266115 389014 266167
rect 389066 266155 389072 266167
rect 392272 266155 392278 266167
rect 389066 266127 392278 266155
rect 389066 266115 389072 266127
rect 392272 266115 392278 266127
rect 392330 266115 392336 266167
rect 541456 266115 541462 266167
rect 541514 266155 541520 266167
rect 542032 266155 542038 266167
rect 541514 266127 542038 266155
rect 541514 266115 541520 266127
rect 542032 266115 542038 266127
rect 542090 266115 542096 266167
rect 381616 266041 381622 266093
rect 381674 266081 381680 266093
rect 622480 266081 622486 266093
rect 381674 266053 622486 266081
rect 381674 266041 381680 266053
rect 622480 266041 622486 266053
rect 622538 266041 622544 266093
rect 379120 265967 379126 266019
rect 379178 266007 379184 266019
rect 383440 266007 383446 266019
rect 379178 265979 383446 266007
rect 379178 265967 379184 265979
rect 383440 265967 383446 265979
rect 383498 265967 383504 266019
rect 398512 265967 398518 266019
rect 398570 266007 398576 266019
rect 597520 266007 597526 266019
rect 398570 265979 597526 266007
rect 398570 265967 398576 265979
rect 597520 265967 597526 265979
rect 597578 265967 597584 266019
rect 383056 265933 383062 265945
rect 378946 265905 383062 265933
rect 286922 265893 286928 265905
rect 383056 265893 383062 265905
rect 383114 265893 383120 265945
rect 386992 265893 386998 265945
rect 387050 265933 387056 265945
rect 396688 265933 396694 265945
rect 387050 265905 396694 265933
rect 387050 265893 387056 265905
rect 396688 265893 396694 265905
rect 396746 265893 396752 265945
rect 265648 265819 265654 265871
rect 265706 265859 265712 265871
rect 265706 265831 267902 265859
rect 265706 265819 265712 265831
rect 267874 265637 267902 265831
rect 282736 265819 282742 265871
rect 282794 265859 282800 265871
rect 394096 265859 394102 265871
rect 282794 265831 394102 265859
rect 282794 265819 282800 265831
rect 394096 265819 394102 265831
rect 394154 265819 394160 265871
rect 279952 265745 279958 265797
rect 280010 265785 280016 265797
rect 378640 265785 378646 265797
rect 280010 265757 378646 265785
rect 280010 265745 280016 265757
rect 378640 265745 378646 265757
rect 378698 265745 378704 265797
rect 384208 265745 384214 265797
rect 384266 265785 384272 265797
rect 398800 265785 398806 265797
rect 384266 265757 398806 265785
rect 384266 265745 384272 265757
rect 398800 265745 398806 265757
rect 398858 265745 398864 265797
rect 287152 265671 287158 265723
rect 287210 265711 287216 265723
rect 392848 265711 392854 265723
rect 287210 265683 392854 265711
rect 287210 265671 287216 265683
rect 392848 265671 392854 265683
rect 392906 265671 392912 265723
rect 427504 265671 427510 265723
rect 427562 265711 427568 265723
rect 438640 265711 438646 265723
rect 427562 265683 438646 265711
rect 427562 265671 427568 265683
rect 438640 265671 438646 265683
rect 438698 265671 438704 265723
rect 287920 265637 287926 265649
rect 267874 265609 287926 265637
rect 287920 265597 287926 265609
rect 287978 265597 287984 265649
rect 328240 265597 328246 265649
rect 328298 265637 328304 265649
rect 429328 265637 429334 265649
rect 328298 265609 429334 265637
rect 328298 265597 328304 265609
rect 429328 265597 429334 265609
rect 429386 265597 429392 265649
rect 327856 265523 327862 265575
rect 327914 265563 327920 265575
rect 429424 265563 429430 265575
rect 327914 265535 429430 265563
rect 327914 265523 327920 265535
rect 429424 265523 429430 265535
rect 429482 265523 429488 265575
rect 287056 265449 287062 265501
rect 287114 265489 287120 265501
rect 375184 265489 375190 265501
rect 287114 265461 375190 265489
rect 287114 265449 287120 265461
rect 375184 265449 375190 265461
rect 375242 265449 375248 265501
rect 386896 265489 386902 265501
rect 375298 265461 386902 265489
rect 286768 265375 286774 265427
rect 286826 265415 286832 265427
rect 375298 265415 375326 265461
rect 386896 265449 386902 265461
rect 386954 265449 386960 265501
rect 286826 265387 375326 265415
rect 286826 265375 286832 265387
rect 375376 265375 375382 265427
rect 375434 265415 375440 265427
rect 389584 265415 389590 265427
rect 375434 265387 389590 265415
rect 375434 265375 375440 265387
rect 389584 265375 389590 265387
rect 389642 265375 389648 265427
rect 389776 265375 389782 265427
rect 389834 265415 389840 265427
rect 593872 265415 593878 265427
rect 389834 265387 593878 265415
rect 389834 265375 389840 265387
rect 593872 265375 593878 265387
rect 593930 265375 593936 265427
rect 329296 265301 329302 265353
rect 329354 265341 329360 265353
rect 424816 265341 424822 265353
rect 329354 265313 424822 265341
rect 329354 265301 329360 265313
rect 424816 265301 424822 265313
rect 424874 265301 424880 265353
rect 294160 265227 294166 265279
rect 294218 265267 294224 265279
rect 390736 265267 390742 265279
rect 294218 265239 390742 265267
rect 294218 265227 294224 265239
rect 390736 265227 390742 265239
rect 390794 265227 390800 265279
rect 405904 265227 405910 265279
rect 405962 265267 405968 265279
rect 423280 265267 423286 265279
rect 405962 265239 423286 265267
rect 405962 265227 405968 265239
rect 423280 265227 423286 265239
rect 423338 265227 423344 265279
rect 301264 265153 301270 265205
rect 301322 265193 301328 265205
rect 301322 265165 375038 265193
rect 301322 265153 301328 265165
rect 329872 265079 329878 265131
rect 329930 265119 329936 265131
rect 374896 265119 374902 265131
rect 329930 265091 374902 265119
rect 329930 265079 329936 265091
rect 374896 265079 374902 265091
rect 374954 265079 374960 265131
rect 375010 265119 375038 265165
rect 378064 265153 378070 265205
rect 378122 265193 378128 265205
rect 378544 265193 378550 265205
rect 378122 265165 378550 265193
rect 378122 265153 378128 265165
rect 378544 265153 378550 265165
rect 378602 265153 378608 265205
rect 378640 265153 378646 265205
rect 378698 265193 378704 265205
rect 389104 265193 389110 265205
rect 378698 265165 389110 265193
rect 378698 265153 378704 265165
rect 389104 265153 389110 265165
rect 389162 265153 389168 265205
rect 391888 265193 391894 265205
rect 389218 265165 391894 265193
rect 389218 265119 389246 265165
rect 391888 265153 391894 265165
rect 391946 265153 391952 265205
rect 394576 265153 394582 265205
rect 394634 265193 394640 265205
rect 398896 265193 398902 265205
rect 394634 265165 398902 265193
rect 394634 265153 394640 265165
rect 398896 265153 398902 265165
rect 398954 265153 398960 265205
rect 375010 265091 389246 265119
rect 283120 265005 283126 265057
rect 283178 265045 283184 265057
rect 425584 265045 425590 265057
rect 283178 265017 425590 265045
rect 283178 265005 283184 265017
rect 425584 265005 425590 265017
rect 425642 265005 425648 265057
rect 429232 265005 429238 265057
rect 429290 265045 429296 265057
rect 443440 265045 443446 265057
rect 429290 265017 443446 265045
rect 429290 265005 429296 265017
rect 443440 265005 443446 265017
rect 443498 265005 443504 265057
rect 251344 264931 251350 264983
rect 251402 264971 251408 264983
rect 386032 264971 386038 264983
rect 251402 264943 386038 264971
rect 251402 264931 251408 264943
rect 386032 264931 386038 264943
rect 386090 264931 386096 264983
rect 421648 264931 421654 264983
rect 421706 264971 421712 264983
rect 432496 264971 432502 264983
rect 421706 264943 432502 264971
rect 421706 264931 421712 264943
rect 432496 264931 432502 264943
rect 432554 264931 432560 264983
rect 271600 264857 271606 264909
rect 271658 264897 271664 264909
rect 318256 264897 318262 264909
rect 271658 264869 318262 264897
rect 271658 264857 271664 264869
rect 318256 264857 318262 264869
rect 318314 264857 318320 264909
rect 325072 264857 325078 264909
rect 325130 264897 325136 264909
rect 329392 264897 329398 264909
rect 325130 264869 329398 264897
rect 325130 264857 325136 264869
rect 329392 264857 329398 264869
rect 329450 264857 329456 264909
rect 329488 264857 329494 264909
rect 329546 264897 329552 264909
rect 344368 264897 344374 264909
rect 329546 264869 344374 264897
rect 329546 264857 329552 264869
rect 344368 264857 344374 264869
rect 344426 264857 344432 264909
rect 359536 264857 359542 264909
rect 359594 264897 359600 264909
rect 499888 264897 499894 264909
rect 359594 264869 499894 264897
rect 359594 264857 359600 264869
rect 499888 264857 499894 264869
rect 499946 264857 499952 264909
rect 267952 264783 267958 264835
rect 268010 264823 268016 264835
rect 318064 264823 318070 264835
rect 268010 264795 318070 264823
rect 268010 264783 268016 264795
rect 318064 264783 318070 264795
rect 318122 264783 318128 264835
rect 329200 264823 329206 264835
rect 318178 264795 329206 264823
rect 264496 264709 264502 264761
rect 264554 264749 264560 264761
rect 318178 264749 318206 264795
rect 329200 264783 329206 264795
rect 329258 264783 329264 264835
rect 339952 264823 339958 264835
rect 333634 264795 339958 264823
rect 333634 264749 333662 264795
rect 339952 264783 339958 264795
rect 340010 264783 340016 264835
rect 359920 264783 359926 264835
rect 359978 264823 359984 264835
rect 506896 264823 506902 264835
rect 359978 264795 506902 264823
rect 359978 264783 359984 264795
rect 506896 264783 506902 264795
rect 506954 264783 506960 264835
rect 264554 264721 318206 264749
rect 318370 264721 333662 264749
rect 264554 264709 264560 264721
rect 257296 264635 257302 264687
rect 257354 264675 257360 264687
rect 318160 264675 318166 264687
rect 257354 264647 318166 264675
rect 257354 264635 257360 264647
rect 318160 264635 318166 264647
rect 318218 264635 318224 264687
rect 260848 264561 260854 264613
rect 260906 264601 260912 264613
rect 318370 264601 318398 264721
rect 333712 264709 333718 264761
rect 333770 264749 333776 264761
rect 340336 264749 340342 264761
rect 333770 264721 340342 264749
rect 333770 264709 333776 264721
rect 340336 264709 340342 264721
rect 340394 264709 340400 264761
rect 360976 264709 360982 264761
rect 361034 264749 361040 264761
rect 524944 264749 524950 264761
rect 361034 264721 524950 264749
rect 361034 264709 361040 264721
rect 524944 264709 524950 264721
rect 525002 264709 525008 264761
rect 318448 264635 318454 264687
rect 318506 264675 318512 264687
rect 339568 264675 339574 264687
rect 318506 264647 339574 264675
rect 318506 264635 318512 264647
rect 339568 264635 339574 264647
rect 339626 264635 339632 264687
rect 360592 264635 360598 264687
rect 360650 264675 360656 264687
rect 517744 264675 517750 264687
rect 360650 264647 517750 264675
rect 360650 264635 360656 264647
rect 517744 264635 517750 264647
rect 517802 264635 517808 264687
rect 260906 264573 318398 264601
rect 260906 264561 260912 264573
rect 318640 264561 318646 264613
rect 318698 264601 318704 264613
rect 333712 264601 333718 264613
rect 318698 264573 333718 264601
rect 318698 264561 318704 264573
rect 333712 264561 333718 264573
rect 333770 264561 333776 264613
rect 339280 264601 339286 264613
rect 333826 264573 339286 264601
rect 253744 264487 253750 264539
rect 253802 264527 253808 264539
rect 333826 264527 333854 264573
rect 339280 264561 339286 264573
rect 339338 264561 339344 264613
rect 361360 264561 361366 264613
rect 361418 264601 361424 264613
rect 532048 264601 532054 264613
rect 361418 264573 532054 264601
rect 361418 264561 361424 264573
rect 532048 264561 532054 264573
rect 532106 264561 532112 264613
rect 253802 264499 333854 264527
rect 253802 264487 253808 264499
rect 335248 264487 335254 264539
rect 335306 264527 335312 264539
rect 356176 264527 356182 264539
rect 335306 264499 356182 264527
rect 335306 264487 335312 264499
rect 356176 264487 356182 264499
rect 356234 264487 356240 264539
rect 361744 264487 361750 264539
rect 361802 264527 361808 264539
rect 539152 264527 539158 264539
rect 361802 264499 539158 264527
rect 361802 264487 361808 264499
rect 539152 264487 539158 264499
rect 539210 264487 539216 264539
rect 283312 264413 283318 264465
rect 283370 264453 283376 264465
rect 371440 264453 371446 264465
rect 283370 264425 371446 264453
rect 283370 264413 283376 264425
rect 371440 264413 371446 264425
rect 371498 264413 371504 264465
rect 374224 264413 374230 264465
rect 374282 264453 374288 264465
rect 558256 264453 558262 264465
rect 374282 264425 558262 264453
rect 374282 264413 374288 264425
rect 558256 264413 558262 264425
rect 558314 264413 558320 264465
rect 250096 264339 250102 264391
rect 250154 264379 250160 264391
rect 338896 264379 338902 264391
rect 250154 264351 338902 264379
rect 250154 264339 250160 264351
rect 338896 264339 338902 264351
rect 338954 264339 338960 264391
rect 347344 264379 347350 264391
rect 339586 264351 347350 264379
rect 42256 264265 42262 264317
rect 42314 264305 42320 264317
rect 53296 264305 53302 264317
rect 42314 264277 53302 264305
rect 42314 264265 42320 264277
rect 53296 264265 53302 264277
rect 53354 264265 53360 264317
rect 246640 264265 246646 264317
rect 246698 264305 246704 264317
rect 338512 264305 338518 264317
rect 246698 264277 338518 264305
rect 246698 264265 246704 264277
rect 338512 264265 338518 264277
rect 338570 264265 338576 264317
rect 338608 264265 338614 264317
rect 338666 264305 338672 264317
rect 339586 264305 339614 264351
rect 347344 264339 347350 264351
rect 347402 264339 347408 264391
rect 362128 264339 362134 264391
rect 362186 264379 362192 264391
rect 546352 264379 546358 264391
rect 362186 264351 546358 264379
rect 362186 264339 362192 264351
rect 546352 264339 546358 264351
rect 546410 264339 546416 264391
rect 341680 264305 341686 264317
rect 338666 264277 339614 264305
rect 339682 264277 341686 264305
rect 338666 264265 338672 264277
rect 243088 264191 243094 264243
rect 243146 264231 243152 264243
rect 338128 264231 338134 264243
rect 243146 264203 338134 264231
rect 243146 264191 243152 264203
rect 338128 264191 338134 264203
rect 338186 264191 338192 264243
rect 339682 264231 339710 264277
rect 341680 264265 341686 264277
rect 341738 264265 341744 264317
rect 375376 264265 375382 264317
rect 375434 264305 375440 264317
rect 568912 264305 568918 264317
rect 375434 264277 568918 264305
rect 375434 264265 375440 264277
rect 568912 264265 568918 264277
rect 568970 264265 568976 264317
rect 338242 264203 339710 264231
rect 214480 264117 214486 264169
rect 214538 264157 214544 264169
rect 335248 264157 335254 264169
rect 214538 264129 335254 264157
rect 214538 264117 214544 264129
rect 335248 264117 335254 264129
rect 335306 264117 335312 264169
rect 335344 264117 335350 264169
rect 335402 264157 335408 264169
rect 338032 264157 338038 264169
rect 335402 264129 338038 264157
rect 335402 264117 335408 264129
rect 338032 264117 338038 264129
rect 338090 264117 338096 264169
rect 196720 264043 196726 264095
rect 196778 264083 196784 264095
rect 312400 264083 312406 264095
rect 196778 264055 312406 264083
rect 196778 264043 196784 264055
rect 312400 264043 312406 264055
rect 312458 264043 312464 264095
rect 318448 264043 318454 264095
rect 318506 264083 318512 264095
rect 338242 264083 338270 264203
rect 339760 264191 339766 264243
rect 339818 264231 339824 264243
rect 368656 264231 368662 264243
rect 339818 264203 368662 264231
rect 339818 264191 339824 264203
rect 368656 264191 368662 264203
rect 368714 264191 368720 264243
rect 374992 264191 374998 264243
rect 375050 264231 375056 264243
rect 565360 264231 565366 264243
rect 375050 264203 565366 264231
rect 375050 264191 375056 264203
rect 565360 264191 565366 264203
rect 565418 264191 565424 264243
rect 352144 264157 352150 264169
rect 318506 264055 338270 264083
rect 338338 264129 352150 264157
rect 318506 264043 318512 264055
rect 200176 263969 200182 264021
rect 200234 264009 200240 264021
rect 329488 264009 329494 264021
rect 200234 263981 329494 264009
rect 200234 263969 200240 263981
rect 329488 263969 329494 263981
rect 329546 263969 329552 264021
rect 329584 263969 329590 264021
rect 329642 264009 329648 264021
rect 338224 264009 338230 264021
rect 329642 263981 338230 264009
rect 329642 263969 329648 263981
rect 338224 263969 338230 263981
rect 338282 263969 338288 264021
rect 207376 263895 207382 263947
rect 207434 263935 207440 263947
rect 338338 263935 338366 264129
rect 352144 264117 352150 264129
rect 352202 264117 352208 264169
rect 375664 264117 375670 264169
rect 375722 264157 375728 264169
rect 572464 264157 572470 264169
rect 375722 264129 572470 264157
rect 375722 264117 375728 264129
rect 572464 264117 572470 264129
rect 572522 264117 572528 264169
rect 340528 264043 340534 264095
rect 340586 264083 340592 264095
rect 360016 264083 360022 264095
rect 340586 264055 360022 264083
rect 340586 264043 340592 264055
rect 360016 264043 360022 264055
rect 360074 264043 360080 264095
rect 376048 264043 376054 264095
rect 376106 264083 376112 264095
rect 576112 264083 576118 264095
rect 376106 264055 576118 264083
rect 376106 264043 376112 264055
rect 576112 264043 576118 264055
rect 576170 264043 576176 264095
rect 338416 263969 338422 264021
rect 338474 264009 338480 264021
rect 346480 264009 346486 264021
rect 338474 263981 346486 264009
rect 338474 263969 338480 263981
rect 346480 263969 346486 263981
rect 346538 263969 346544 264021
rect 347728 263969 347734 264021
rect 347786 264009 347792 264021
rect 368464 264009 368470 264021
rect 347786 263981 368470 264009
rect 347786 263969 347792 263981
rect 368464 263969 368470 263981
rect 368522 263969 368528 264021
rect 376432 263969 376438 264021
rect 376490 264009 376496 264021
rect 579664 264009 579670 264021
rect 376490 263981 579670 264009
rect 376490 263969 376496 263981
rect 579664 263969 579670 263981
rect 579722 263969 579728 264021
rect 207434 263907 338366 263935
rect 207434 263895 207440 263907
rect 338704 263895 338710 263947
rect 338762 263935 338768 263947
rect 340720 263935 340726 263947
rect 338762 263907 340726 263935
rect 338762 263895 338768 263907
rect 340720 263895 340726 263907
rect 340778 263895 340784 263947
rect 377584 263895 377590 263947
rect 377642 263935 377648 263947
rect 586768 263935 586774 263947
rect 377642 263907 586774 263935
rect 377642 263895 377648 263907
rect 586768 263895 586774 263907
rect 586826 263895 586832 263947
rect 203728 263821 203734 263873
rect 203786 263861 203792 263873
rect 348496 263861 348502 263873
rect 203786 263833 348502 263861
rect 203786 263821 203792 263833
rect 348496 263821 348502 263833
rect 348554 263821 348560 263873
rect 352528 263821 352534 263873
rect 352586 263861 352592 263873
rect 375088 263861 375094 263873
rect 352586 263833 375094 263861
rect 352586 263821 352592 263833
rect 375088 263821 375094 263833
rect 375146 263821 375152 263873
rect 376816 263821 376822 263873
rect 376874 263861 376880 263873
rect 583120 263861 583126 263873
rect 376874 263833 583126 263861
rect 376874 263821 376880 263833
rect 583120 263821 583126 263833
rect 583178 263821 583184 263873
rect 239440 263747 239446 263799
rect 239498 263787 239504 263799
rect 337744 263787 337750 263799
rect 239498 263759 337750 263787
rect 239498 263747 239504 263759
rect 337744 263747 337750 263759
rect 337802 263747 337808 263799
rect 337840 263747 337846 263799
rect 337898 263787 337904 263799
rect 592720 263787 592726 263799
rect 337898 263759 592726 263787
rect 337898 263747 337904 263759
rect 592720 263747 592726 263759
rect 592778 263747 592784 263799
rect 228784 263673 228790 263725
rect 228842 263713 228848 263725
rect 228842 263685 314462 263713
rect 228842 263673 228848 263685
rect 232336 263599 232342 263651
rect 232394 263639 232400 263651
rect 314320 263639 314326 263651
rect 232394 263611 314326 263639
rect 232394 263599 232400 263611
rect 314320 263599 314326 263611
rect 314378 263599 314384 263651
rect 314434 263639 314462 263685
rect 318064 263673 318070 263725
rect 318122 263713 318128 263725
rect 318122 263685 333566 263713
rect 318122 263673 318128 263685
rect 330064 263639 330070 263651
rect 314434 263611 330070 263639
rect 330064 263599 330070 263611
rect 330122 263599 330128 263651
rect 330160 263599 330166 263651
rect 330218 263639 330224 263651
rect 333538 263639 333566 263685
rect 339664 263673 339670 263725
rect 339722 263713 339728 263725
rect 624784 263713 624790 263725
rect 339722 263685 624790 263713
rect 339722 263673 339728 263685
rect 624784 263673 624790 263685
rect 624842 263673 624848 263725
rect 330218 263611 333470 263639
rect 333538 263611 335006 263639
rect 330218 263599 330224 263611
rect 42256 263525 42262 263577
rect 42314 263565 42320 263577
rect 53392 263565 53398 263577
rect 42314 263537 53398 263565
rect 42314 263525 42320 263537
rect 53392 263525 53398 263537
rect 53450 263525 53456 263577
rect 275152 263525 275158 263577
rect 275210 263565 275216 263577
rect 318448 263565 318454 263577
rect 275210 263537 318454 263565
rect 275210 263525 275216 263537
rect 318448 263525 318454 263537
rect 318506 263525 318512 263577
rect 318544 263525 318550 263577
rect 318602 263565 318608 263577
rect 329584 263565 329590 263577
rect 318602 263537 329590 263565
rect 318602 263525 318608 263537
rect 329584 263525 329590 263537
rect 329642 263525 329648 263577
rect 329680 263525 329686 263577
rect 329738 263565 329744 263577
rect 333232 263565 333238 263577
rect 329738 263537 333238 263565
rect 329738 263525 329744 263537
rect 333232 263525 333238 263537
rect 333290 263525 333296 263577
rect 333442 263565 333470 263611
rect 334864 263565 334870 263577
rect 333442 263537 334870 263565
rect 334864 263525 334870 263537
rect 334922 263525 334928 263577
rect 334978 263565 335006 263611
rect 335344 263599 335350 263651
rect 335402 263639 335408 263651
rect 628432 263639 628438 263651
rect 335402 263611 628438 263639
rect 335402 263599 335408 263611
rect 628432 263599 628438 263611
rect 628490 263599 628496 263651
rect 341104 263565 341110 263577
rect 334978 263537 341110 263565
rect 341104 263525 341110 263537
rect 341162 263525 341168 263577
rect 368560 263565 368566 263577
rect 357922 263537 368566 263565
rect 318160 263451 318166 263503
rect 318218 263491 318224 263503
rect 342544 263491 342550 263503
rect 318218 263463 342550 263491
rect 318218 263451 318224 263463
rect 342544 263451 342550 263463
rect 342602 263451 342608 263503
rect 285808 263377 285814 263429
rect 285866 263417 285872 263429
rect 342832 263417 342838 263429
rect 285866 263389 342838 263417
rect 285866 263377 285872 263389
rect 342832 263377 342838 263389
rect 342890 263377 342896 263429
rect 278704 263303 278710 263355
rect 278762 263343 278768 263355
rect 342160 263343 342166 263355
rect 278762 263315 342166 263343
rect 278762 263303 278768 263315
rect 342160 263303 342166 263315
rect 342218 263303 342224 263355
rect 282928 263229 282934 263281
rect 282986 263269 282992 263281
rect 318160 263269 318166 263281
rect 282986 263241 318166 263269
rect 282986 263229 282992 263241
rect 318160 263229 318166 263241
rect 318218 263229 318224 263281
rect 319120 263229 319126 263281
rect 319178 263269 319184 263281
rect 333136 263269 333142 263281
rect 319178 263241 333142 263269
rect 319178 263229 319184 263241
rect 333136 263229 333142 263241
rect 333194 263229 333200 263281
rect 333232 263229 333238 263281
rect 333290 263269 333296 263281
rect 357922 263269 357950 263537
rect 368560 263525 368566 263537
rect 368618 263525 368624 263577
rect 383152 263525 383158 263577
rect 383210 263565 383216 263577
rect 386800 263565 386806 263577
rect 383210 263537 386806 263565
rect 383210 263525 383216 263537
rect 386800 263525 386806 263537
rect 386858 263525 386864 263577
rect 423568 263525 423574 263577
rect 423626 263565 423632 263577
rect 430384 263565 430390 263577
rect 423626 263537 430390 263565
rect 423626 263525 423632 263537
rect 430384 263525 430390 263537
rect 430442 263525 430448 263577
rect 535696 263525 535702 263577
rect 535754 263565 535760 263577
rect 536176 263565 536182 263577
rect 535754 263537 536182 263565
rect 535754 263525 535760 263537
rect 536176 263525 536182 263537
rect 536234 263525 536240 263577
rect 359152 263451 359158 263503
rect 359210 263491 359216 263503
rect 492784 263491 492790 263503
rect 359210 263463 492790 263491
rect 359210 263451 359216 263463
rect 492784 263451 492790 263463
rect 492842 263451 492848 263503
rect 358768 263377 358774 263429
rect 358826 263417 358832 263429
rect 485584 263417 485590 263429
rect 358826 263389 485590 263417
rect 358826 263377 358832 263389
rect 485584 263377 485590 263389
rect 485642 263377 485648 263429
rect 358384 263303 358390 263355
rect 358442 263343 358448 263355
rect 478576 263343 478582 263355
rect 358442 263315 478582 263343
rect 358442 263303 358448 263315
rect 478576 263303 478582 263315
rect 478634 263303 478640 263355
rect 333290 263241 357950 263269
rect 333290 263229 333296 263241
rect 358000 263229 358006 263281
rect 358058 263269 358064 263281
rect 474928 263269 474934 263281
rect 358058 263241 474934 263269
rect 358058 263229 358064 263241
rect 474928 263229 474934 263241
rect 474986 263229 474992 263281
rect 289456 263155 289462 263207
rect 289514 263195 289520 263207
rect 343312 263195 343318 263207
rect 289514 263167 343318 263195
rect 289514 263155 289520 263167
rect 343312 263155 343318 263167
rect 343370 263155 343376 263207
rect 357712 263155 357718 263207
rect 357770 263195 357776 263207
rect 467824 263195 467830 263207
rect 357770 263167 467830 263195
rect 357770 263155 357776 263167
rect 467824 263155 467830 263167
rect 467882 263155 467888 263207
rect 236176 263121 236182 263133
rect 167074 263093 189662 263121
rect 124048 263007 124054 263059
rect 124106 263047 124112 263059
rect 141136 263047 141142 263059
rect 124106 263019 141142 263047
rect 124106 263007 124112 263019
rect 141136 263007 141142 263019
rect 141194 263007 141200 263059
rect 149392 263007 149398 263059
rect 149450 263047 149456 263059
rect 167074 263047 167102 263093
rect 149450 263019 167102 263047
rect 189634 263047 189662 263093
rect 236098 263093 236182 263121
rect 189634 263019 201662 263047
rect 149450 263007 149456 263019
rect 141136 262859 141142 262911
rect 141194 262899 141200 262911
rect 149392 262899 149398 262911
rect 141194 262871 149398 262899
rect 141194 262859 141200 262871
rect 149392 262859 149398 262871
rect 149450 262859 149456 262911
rect 201634 262899 201662 263019
rect 221680 262973 221686 262985
rect 216034 262945 221686 262973
rect 216034 262899 216062 262945
rect 221680 262933 221686 262945
rect 221738 262933 221744 262985
rect 221776 262933 221782 262985
rect 221834 262973 221840 262985
rect 236098 262973 236126 263093
rect 236176 263081 236182 263093
rect 236234 263081 236240 263133
rect 262096 263081 262102 263133
rect 262154 263081 262160 263133
rect 262288 263081 262294 263133
rect 262346 263121 262352 263133
rect 262346 263093 287774 263121
rect 262346 263081 262352 263093
rect 236272 263007 236278 263059
rect 236330 263047 236336 263059
rect 262114 263047 262142 263081
rect 236330 263019 262142 263047
rect 287746 263047 287774 263093
rect 293008 263081 293014 263133
rect 293066 263121 293072 263133
rect 343696 263121 343702 263133
rect 293066 263093 343702 263121
rect 293066 263081 293072 263093
rect 343696 263081 343702 263093
rect 343754 263081 343760 263133
rect 357328 263081 357334 263133
rect 357386 263121 357392 263133
rect 460720 263121 460726 263133
rect 357386 263093 460726 263121
rect 357386 263081 357392 263093
rect 460720 263081 460726 263093
rect 460778 263081 460784 263133
rect 325456 263047 325462 263059
rect 287746 263019 325462 263047
rect 236330 263007 236336 263019
rect 325456 263007 325462 263019
rect 325514 263007 325520 263059
rect 328048 263007 328054 263059
rect 328106 263047 328112 263059
rect 333520 263047 333526 263059
rect 328106 263019 333526 263047
rect 328106 263007 328112 263019
rect 333520 263007 333526 263019
rect 333578 263007 333584 263059
rect 333616 263007 333622 263059
rect 333674 263047 333680 263059
rect 333674 263019 341726 263047
rect 333674 263007 333680 263019
rect 221834 262945 236126 262973
rect 221834 262933 221840 262945
rect 331504 262933 331510 262985
rect 331562 262973 331568 262985
rect 341698 262973 341726 263019
rect 368560 263007 368566 263059
rect 368618 263047 368624 263059
rect 427792 263047 427798 263059
rect 368618 263019 427798 263047
rect 368618 263007 368624 263019
rect 427792 263007 427798 263019
rect 427850 263007 427856 263059
rect 429520 262973 429526 262985
rect 331562 262945 341630 262973
rect 341698 262945 429526 262973
rect 331562 262933 331568 262945
rect 201634 262871 216062 262899
rect 318256 262859 318262 262911
rect 318314 262899 318320 262911
rect 341488 262899 341494 262911
rect 318314 262871 341494 262899
rect 318314 262859 318320 262871
rect 341488 262859 341494 262871
rect 341546 262859 341552 262911
rect 341602 262899 341630 262945
rect 429520 262933 429526 262945
rect 429578 262933 429584 262985
rect 429616 262899 429622 262911
rect 341602 262871 429622 262899
rect 429616 262859 429622 262871
rect 429674 262859 429680 262911
rect 296560 262785 296566 262837
rect 296618 262825 296624 262837
rect 344080 262825 344086 262837
rect 296618 262797 344086 262825
rect 296618 262785 296624 262797
rect 344080 262785 344086 262797
rect 344138 262785 344144 262837
rect 356944 262785 356950 262837
rect 357002 262825 357008 262837
rect 453520 262825 453526 262837
rect 357002 262797 453526 262825
rect 357002 262785 357008 262797
rect 453520 262785 453526 262797
rect 453578 262785 453584 262837
rect 286384 262711 286390 262763
rect 286442 262751 286448 262763
rect 369040 262751 369046 262763
rect 286442 262723 369046 262751
rect 286442 262711 286448 262723
rect 369040 262711 369046 262723
rect 369098 262711 369104 262763
rect 383440 262711 383446 262763
rect 383498 262751 383504 262763
rect 384016 262751 384022 262763
rect 383498 262723 384022 262751
rect 383498 262711 383504 262723
rect 384016 262711 384022 262723
rect 384074 262711 384080 262763
rect 426256 262711 426262 262763
rect 426314 262751 426320 262763
rect 434896 262751 434902 262763
rect 426314 262723 434902 262751
rect 426314 262711 426320 262723
rect 434896 262711 434902 262723
rect 434954 262711 434960 262763
rect 300112 262637 300118 262689
rect 300170 262677 300176 262689
rect 344752 262677 344758 262689
rect 300170 262649 344758 262677
rect 300170 262637 300176 262649
rect 344752 262637 344758 262649
rect 344810 262637 344816 262689
rect 355792 262637 355798 262689
rect 355850 262677 355856 262689
rect 435664 262677 435670 262689
rect 355850 262649 435670 262677
rect 355850 262637 355856 262649
rect 435664 262637 435670 262649
rect 435722 262637 435728 262689
rect 303664 262563 303670 262615
rect 303722 262603 303728 262615
rect 345136 262603 345142 262615
rect 303722 262575 345142 262603
rect 303722 262563 303728 262575
rect 345136 262563 345142 262575
rect 345194 262563 345200 262615
rect 355504 262563 355510 262615
rect 355562 262603 355568 262615
rect 428560 262603 428566 262615
rect 355562 262575 428566 262603
rect 355562 262563 355568 262575
rect 428560 262563 428566 262575
rect 428618 262563 428624 262615
rect 310864 262489 310870 262541
rect 310922 262529 310928 262541
rect 345904 262529 345910 262541
rect 310922 262501 345910 262529
rect 310922 262489 310928 262501
rect 345904 262489 345910 262501
rect 345962 262489 345968 262541
rect 355120 262489 355126 262541
rect 355178 262529 355184 262541
rect 421456 262529 421462 262541
rect 355178 262501 421462 262529
rect 355178 262489 355184 262501
rect 421456 262489 421462 262501
rect 421514 262489 421520 262541
rect 426448 262489 426454 262541
rect 426506 262529 426512 262541
rect 437488 262529 437494 262541
rect 426506 262501 437494 262529
rect 426506 262489 426512 262501
rect 437488 262489 437494 262501
rect 437546 262489 437552 262541
rect 307216 262415 307222 262467
rect 307274 262455 307280 262467
rect 345520 262455 345526 262467
rect 307274 262427 345526 262455
rect 307274 262415 307280 262427
rect 345520 262415 345526 262427
rect 345578 262415 345584 262467
rect 354736 262415 354742 262467
rect 354794 262455 354800 262467
rect 414352 262455 414358 262467
rect 354794 262427 414358 262455
rect 354794 262415 354800 262427
rect 414352 262415 414358 262427
rect 414410 262415 414416 262467
rect 312016 262341 312022 262393
rect 312074 262381 312080 262393
rect 366832 262381 366838 262393
rect 312074 262353 366838 262381
rect 312074 262341 312080 262353
rect 366832 262341 366838 262353
rect 366890 262341 366896 262393
rect 383056 262341 383062 262393
rect 383114 262381 383120 262393
rect 397648 262381 397654 262393
rect 383114 262353 397654 262381
rect 383114 262341 383120 262353
rect 397648 262341 397654 262353
rect 397706 262341 397712 262393
rect 42832 262267 42838 262319
rect 42890 262307 42896 262319
rect 58960 262307 58966 262319
rect 42890 262279 58966 262307
rect 42890 262267 42896 262279
rect 58960 262267 58966 262279
rect 59018 262267 59024 262319
rect 314416 262267 314422 262319
rect 314474 262307 314480 262319
rect 346288 262307 346294 262319
rect 314474 262279 346294 262307
rect 314474 262267 314480 262279
rect 346288 262267 346294 262279
rect 346346 262267 346352 262319
rect 353968 262267 353974 262319
rect 354026 262307 354032 262319
rect 391792 262307 391798 262319
rect 354026 262279 391798 262307
rect 354026 262267 354032 262279
rect 391792 262267 391798 262279
rect 391850 262267 391856 262319
rect 314320 262193 314326 262245
rect 314378 262233 314384 262245
rect 334096 262233 334102 262245
rect 314378 262205 334102 262233
rect 314378 262193 314384 262205
rect 334096 262193 334102 262205
rect 334154 262193 334160 262245
rect 346960 262233 346966 262245
rect 336994 262205 346966 262233
rect 301840 262119 301846 262171
rect 301898 262159 301904 262171
rect 302032 262159 302038 262171
rect 301898 262131 302038 262159
rect 301898 262119 301904 262131
rect 302032 262119 302038 262131
rect 302090 262119 302096 262171
rect 321520 262119 321526 262171
rect 321578 262159 321584 262171
rect 336994 262159 337022 262205
rect 346960 262193 346966 262205
rect 347018 262193 347024 262245
rect 353680 262193 353686 262245
rect 353738 262233 353744 262245
rect 388912 262233 388918 262245
rect 353738 262205 388918 262233
rect 353738 262193 353744 262205
rect 388912 262193 388918 262205
rect 388970 262193 388976 262245
rect 321578 262131 337022 262159
rect 321578 262119 321584 262131
rect 337072 262119 337078 262171
rect 337130 262159 337136 262171
rect 646288 262159 646294 262171
rect 337130 262131 646294 262159
rect 337130 262119 337136 262131
rect 646288 262119 646294 262131
rect 646346 262119 646352 262171
rect 256144 262045 256150 262097
rect 256202 262085 256208 262097
rect 296944 262085 296950 262097
rect 256202 262057 296950 262085
rect 256202 262045 256208 262057
rect 296944 262045 296950 262057
rect 297002 262045 297008 262097
rect 310288 262045 310294 262097
rect 310346 262085 310352 262097
rect 466576 262085 466582 262097
rect 310346 262057 466582 262085
rect 310346 262045 310352 262057
rect 466576 262045 466582 262057
rect 466634 262045 466640 262097
rect 249040 261971 249046 262023
rect 249098 262011 249104 262023
rect 296560 262011 296566 262023
rect 249098 261983 296566 262011
rect 249098 261971 249104 261983
rect 296560 261971 296566 261983
rect 296618 261971 296624 262023
rect 311344 261971 311350 262023
rect 311402 262011 311408 262023
rect 477328 262011 477334 262023
rect 311402 261983 477334 262011
rect 311402 261971 311408 261983
rect 477328 261971 477334 261983
rect 477386 261971 477392 262023
rect 231184 261897 231190 261949
rect 231242 261937 231248 261949
rect 231242 261909 234206 261937
rect 231242 261897 231248 261909
rect 175216 261823 175222 261875
rect 175274 261863 175280 261875
rect 234064 261863 234070 261875
rect 175274 261835 234070 261863
rect 175274 261823 175280 261835
rect 234064 261823 234070 261835
rect 234122 261823 234128 261875
rect 168016 261749 168022 261801
rect 168074 261789 168080 261801
rect 233200 261789 233206 261801
rect 168074 261761 233206 261789
rect 168074 261749 168080 261761
rect 233200 261749 233206 261761
rect 233258 261749 233264 261801
rect 234178 261789 234206 261909
rect 245392 261897 245398 261949
rect 245450 261937 245456 261949
rect 296176 261937 296182 261949
rect 245450 261909 296182 261937
rect 245450 261897 245456 261909
rect 296176 261897 296182 261909
rect 296234 261897 296240 261949
rect 310096 261897 310102 261949
rect 310154 261937 310160 261949
rect 473776 261937 473782 261949
rect 310154 261909 473782 261937
rect 310154 261897 310160 261909
rect 473776 261897 473782 261909
rect 473834 261897 473840 261949
rect 238288 261823 238294 261875
rect 238346 261863 238352 261875
rect 295792 261863 295798 261875
rect 238346 261835 295798 261863
rect 238346 261823 238352 261835
rect 295792 261823 295798 261835
rect 295850 261823 295856 261875
rect 311632 261823 311638 261875
rect 311690 261863 311696 261875
rect 484432 261863 484438 261875
rect 311690 261835 484438 261863
rect 311690 261823 311696 261835
rect 484432 261823 484438 261835
rect 484490 261823 484496 261875
rect 277072 261789 277078 261801
rect 234178 261761 277078 261789
rect 277072 261749 277078 261761
rect 277130 261749 277136 261801
rect 312016 261749 312022 261801
rect 312074 261789 312080 261801
rect 491632 261789 491638 261801
rect 312074 261761 491638 261789
rect 312074 261749 312080 261761
rect 491632 261749 491638 261761
rect 491690 261749 491696 261801
rect 303184 261675 303190 261727
rect 303242 261715 303248 261727
rect 334576 261715 334582 261727
rect 303242 261687 334582 261715
rect 303242 261675 303248 261687
rect 334576 261675 334582 261687
rect 334634 261675 334640 261727
rect 373840 261675 373846 261727
rect 373898 261715 373904 261727
rect 554608 261715 554614 261727
rect 373898 261687 554614 261715
rect 373898 261675 373904 261687
rect 554608 261675 554614 261687
rect 554666 261675 554672 261727
rect 303952 261601 303958 261653
rect 304010 261641 304016 261653
rect 348880 261641 348886 261653
rect 304010 261613 348886 261641
rect 304010 261601 304016 261613
rect 348880 261601 348886 261613
rect 348938 261601 348944 261653
rect 353296 261601 353302 261653
rect 353354 261641 353360 261653
rect 366256 261641 366262 261653
rect 353354 261613 366262 261641
rect 353354 261601 353360 261613
rect 366256 261601 366262 261613
rect 366314 261601 366320 261653
rect 374608 261601 374614 261653
rect 374666 261641 374672 261653
rect 561808 261641 561814 261653
rect 374666 261613 561814 261641
rect 374666 261601 374672 261613
rect 561808 261601 561814 261613
rect 561866 261601 561872 261653
rect 185872 261527 185878 261579
rect 185930 261567 185936 261579
rect 201616 261567 201622 261579
rect 185930 261539 201622 261567
rect 185930 261527 185936 261539
rect 201616 261527 201622 261539
rect 201674 261527 201680 261579
rect 206128 261527 206134 261579
rect 206186 261567 206192 261579
rect 305008 261567 305014 261579
rect 206186 261539 305014 261567
rect 206186 261527 206192 261539
rect 305008 261527 305014 261539
rect 305066 261527 305072 261579
rect 312784 261527 312790 261579
rect 312842 261567 312848 261579
rect 312842 261539 326270 261567
rect 312842 261527 312848 261539
rect 191920 261453 191926 261505
rect 191978 261493 191984 261505
rect 288784 261493 288790 261505
rect 191978 261465 288790 261493
rect 191978 261453 191984 261465
rect 288784 261453 288790 261465
rect 288842 261453 288848 261505
rect 313552 261453 313558 261505
rect 313610 261493 313616 261505
rect 326242 261493 326270 261539
rect 326320 261527 326326 261579
rect 326378 261567 326384 261579
rect 498832 261567 498838 261579
rect 326378 261539 498838 261567
rect 326378 261527 326384 261539
rect 498832 261527 498838 261539
rect 498890 261527 498896 261579
rect 505840 261493 505846 261505
rect 313610 261465 326174 261493
rect 326242 261465 505846 261493
rect 313610 261453 313616 261465
rect 80656 261379 80662 261431
rect 80714 261419 80720 261431
rect 83536 261419 83542 261431
rect 80714 261391 83542 261419
rect 80714 261379 80720 261391
rect 83536 261379 83542 261391
rect 83594 261379 83600 261431
rect 199024 261379 199030 261431
rect 199082 261419 199088 261431
rect 299920 261419 299926 261431
rect 199082 261391 299926 261419
rect 199082 261379 199088 261391
rect 299920 261379 299926 261391
rect 299978 261379 299984 261431
rect 326032 261419 326038 261431
rect 314338 261391 326038 261419
rect 193072 261305 193078 261357
rect 193130 261345 193136 261357
rect 314338 261345 314366 261391
rect 326032 261379 326038 261391
rect 326090 261379 326096 261431
rect 326146 261419 326174 261465
rect 505840 261453 505846 261465
rect 505898 261453 505904 261505
rect 516496 261419 516502 261431
rect 326146 261391 516502 261419
rect 516496 261379 516502 261391
rect 516554 261379 516560 261431
rect 331024 261345 331030 261357
rect 193130 261317 314366 261345
rect 314434 261317 331030 261345
rect 193130 261305 193136 261317
rect 195472 261231 195478 261283
rect 195530 261271 195536 261283
rect 297328 261271 297334 261283
rect 195530 261243 297334 261271
rect 195530 261231 195536 261243
rect 297328 261231 297334 261243
rect 297386 261231 297392 261283
rect 302800 261231 302806 261283
rect 302858 261271 302864 261283
rect 314434 261271 314462 261317
rect 331024 261305 331030 261317
rect 331082 261305 331088 261357
rect 354256 261305 354262 261357
rect 354314 261345 354320 261357
rect 366160 261345 366166 261357
rect 354314 261317 366166 261345
rect 354314 261305 354320 261317
rect 366160 261305 366166 261317
rect 366218 261305 366224 261357
rect 366256 261305 366262 261357
rect 366314 261345 366320 261357
rect 389296 261345 389302 261357
rect 366314 261317 389302 261345
rect 366314 261305 366320 261317
rect 389296 261305 389302 261317
rect 389354 261305 389360 261357
rect 424240 261305 424246 261357
rect 424298 261345 424304 261357
rect 430864 261345 430870 261357
rect 424298 261317 430870 261345
rect 424298 261305 424304 261317
rect 430864 261305 430870 261317
rect 430922 261305 430928 261357
rect 302858 261243 314462 261271
rect 302858 261231 302864 261243
rect 314512 261231 314518 261283
rect 314570 261271 314576 261283
rect 314570 261243 324062 261271
rect 314570 261231 314576 261243
rect 177616 261157 177622 261209
rect 177674 261197 177680 261209
rect 288880 261197 288886 261209
rect 177674 261169 288886 261197
rect 177674 261157 177680 261169
rect 288880 261157 288886 261169
rect 288938 261157 288944 261209
rect 302608 261157 302614 261209
rect 302666 261197 302672 261209
rect 323920 261197 323926 261209
rect 302666 261169 323926 261197
rect 302666 261157 302672 261169
rect 323920 261157 323926 261169
rect 323978 261157 323984 261209
rect 324034 261197 324062 261243
rect 324112 261231 324118 261283
rect 324170 261271 324176 261283
rect 523696 261271 523702 261283
rect 324170 261243 523702 261271
rect 324170 261231 324176 261243
rect 523696 261231 523702 261243
rect 523754 261231 523760 261283
rect 530896 261197 530902 261209
rect 324034 261169 530902 261197
rect 530896 261157 530902 261169
rect 530954 261157 530960 261209
rect 181264 261083 181270 261135
rect 181322 261123 181328 261135
rect 302416 261123 302422 261135
rect 181322 261095 302422 261123
rect 181322 261083 181328 261095
rect 302416 261083 302422 261095
rect 302474 261083 302480 261135
rect 314608 261083 314614 261135
rect 314666 261123 314672 261135
rect 538000 261123 538006 261135
rect 314666 261095 538006 261123
rect 314666 261083 314672 261095
rect 538000 261083 538006 261095
rect 538058 261083 538064 261135
rect 170416 261009 170422 261061
rect 170474 261049 170480 261061
rect 302512 261049 302518 261061
rect 170474 261021 302518 261049
rect 170474 261009 170480 261021
rect 302512 261009 302518 261021
rect 302570 261009 302576 261061
rect 313840 261009 313846 261061
rect 313898 261049 313904 261061
rect 324112 261049 324118 261061
rect 313898 261021 324118 261049
rect 313898 261009 313904 261021
rect 324112 261009 324118 261021
rect 324170 261009 324176 261061
rect 326416 261009 326422 261061
rect 326474 261049 326480 261061
rect 549808 261049 549814 261061
rect 326474 261021 549814 261049
rect 326474 261009 326480 261021
rect 549808 261009 549814 261021
rect 549866 261009 549872 261061
rect 279472 260935 279478 260987
rect 279530 260975 279536 260987
rect 299440 260975 299446 260987
rect 279530 260947 299446 260975
rect 279530 260935 279536 260947
rect 299440 260935 299446 260947
rect 299498 260935 299504 260987
rect 312400 260935 312406 260987
rect 312458 260975 312464 260987
rect 326320 260975 326326 260987
rect 312458 260947 326326 260975
rect 312458 260935 312464 260947
rect 326320 260935 326326 260947
rect 326378 260935 326384 260987
rect 326800 260935 326806 260987
rect 326858 260975 326864 260987
rect 553456 260975 553462 260987
rect 326858 260947 553462 260975
rect 326858 260935 326864 260947
rect 553456 260935 553462 260947
rect 553514 260935 553520 260987
rect 149104 260861 149110 260913
rect 149162 260901 149168 260913
rect 305488 260901 305494 260913
rect 149162 260873 305494 260901
rect 149162 260861 149168 260873
rect 305488 260861 305494 260873
rect 305546 260861 305552 260913
rect 305680 260861 305686 260913
rect 305738 260901 305744 260913
rect 373552 260901 373558 260913
rect 305738 260873 373558 260901
rect 305738 260861 305744 260873
rect 373552 260861 373558 260873
rect 373610 260861 373616 260913
rect 380464 260861 380470 260913
rect 380522 260901 380528 260913
rect 615376 260901 615382 260913
rect 380522 260873 615382 260901
rect 380522 260861 380528 260873
rect 615376 260861 615382 260873
rect 615434 260861 615440 260913
rect 158434 260799 178526 260827
rect 138352 260713 138358 260765
rect 138410 260753 138416 260765
rect 158434 260753 158462 260799
rect 138410 260725 158462 260753
rect 178498 260753 178526 260799
rect 298210 260799 299486 260827
rect 298210 260753 298238 260799
rect 178498 260725 298238 260753
rect 299458 260753 299486 260799
rect 303568 260787 303574 260839
rect 303626 260827 303632 260839
rect 341776 260827 341782 260839
rect 303626 260799 341782 260827
rect 303626 260787 303632 260799
rect 341776 260787 341782 260799
rect 341834 260787 341840 260839
rect 341872 260787 341878 260839
rect 341930 260827 341936 260839
rect 574864 260827 574870 260839
rect 341930 260799 574870 260827
rect 341930 260787 341936 260799
rect 574864 260787 574870 260799
rect 574922 260787 574928 260839
rect 305584 260753 305590 260765
rect 299458 260725 305590 260753
rect 138410 260713 138416 260725
rect 305584 260713 305590 260725
rect 305642 260713 305648 260765
rect 305776 260713 305782 260765
rect 305834 260753 305840 260765
rect 380752 260753 380758 260765
rect 305834 260725 380758 260753
rect 305834 260713 305840 260725
rect 380752 260713 380758 260725
rect 380810 260713 380816 260765
rect 380848 260713 380854 260765
rect 380906 260753 380912 260765
rect 618832 260753 618838 260765
rect 380906 260725 618838 260753
rect 380906 260713 380912 260725
rect 618832 260713 618838 260725
rect 618890 260713 618896 260765
rect 131248 260639 131254 260691
rect 131306 260679 131312 260691
rect 198736 260679 198742 260691
rect 131306 260651 198742 260679
rect 131306 260639 131312 260651
rect 198736 260639 198742 260651
rect 198794 260639 198800 260691
rect 279376 260679 279382 260691
rect 218818 260651 279382 260679
rect 218818 260617 218846 260651
rect 279376 260639 279382 260651
rect 279434 260639 279440 260691
rect 299440 260639 299446 260691
rect 299498 260679 299504 260691
rect 299632 260679 299638 260691
rect 299498 260651 299638 260679
rect 299498 260639 299504 260651
rect 299632 260639 299638 260651
rect 299690 260639 299696 260691
rect 304720 260639 304726 260691
rect 304778 260679 304784 260691
rect 304778 260651 308702 260679
rect 304778 260639 304784 260651
rect 218032 260565 218038 260617
rect 218090 260605 218096 260617
rect 218704 260605 218710 260617
rect 218090 260577 218710 260605
rect 218090 260565 218096 260577
rect 218704 260565 218710 260577
rect 218762 260565 218768 260617
rect 218800 260565 218806 260617
rect 218858 260565 218864 260617
rect 263248 260565 263254 260617
rect 263306 260605 263312 260617
rect 297712 260605 297718 260617
rect 263306 260577 297718 260605
rect 263306 260565 263312 260577
rect 297712 260565 297718 260577
rect 297770 260565 297776 260617
rect 308674 260605 308702 260651
rect 308752 260639 308758 260691
rect 308810 260679 308816 260691
rect 313264 260679 313270 260691
rect 308810 260651 313270 260679
rect 308810 260639 308816 260651
rect 313264 260639 313270 260651
rect 313322 260639 313328 260691
rect 328624 260639 328630 260691
rect 328682 260679 328688 260691
rect 571312 260679 571318 260691
rect 328682 260651 571318 260679
rect 328682 260639 328688 260651
rect 571312 260639 571318 260651
rect 571370 260639 571376 260691
rect 363184 260605 363190 260617
rect 308674 260577 363190 260605
rect 363184 260565 363190 260577
rect 363242 260565 363248 260617
rect 373456 260565 373462 260617
rect 373514 260605 373520 260617
rect 521968 260605 521974 260617
rect 373514 260577 521974 260605
rect 373514 260565 373520 260577
rect 521968 260565 521974 260577
rect 522026 260565 522032 260617
rect 270352 260491 270358 260543
rect 270410 260531 270416 260543
rect 298000 260531 298006 260543
rect 270410 260503 298006 260531
rect 270410 260491 270416 260503
rect 298000 260491 298006 260503
rect 298058 260491 298064 260543
rect 310192 260491 310198 260543
rect 310250 260531 310256 260543
rect 459472 260531 459478 260543
rect 310250 260503 459478 260531
rect 310250 260491 310256 260503
rect 459472 260491 459478 260503
rect 459530 260491 459536 260543
rect 277552 260417 277558 260469
rect 277610 260457 277616 260469
rect 298384 260457 298390 260469
rect 277610 260429 298390 260457
rect 277610 260417 277616 260429
rect 298384 260417 298390 260429
rect 298442 260417 298448 260469
rect 309808 260417 309814 260469
rect 309866 260457 309872 260469
rect 452368 260457 452374 260469
rect 309866 260429 452374 260457
rect 309866 260417 309872 260429
rect 452368 260417 452374 260429
rect 452426 260417 452432 260469
rect 216784 260343 216790 260395
rect 216842 260383 216848 260395
rect 218800 260383 218806 260395
rect 216842 260355 218806 260383
rect 216842 260343 216848 260355
rect 218800 260343 218806 260355
rect 218858 260343 218864 260395
rect 220432 260343 220438 260395
rect 220490 260383 220496 260395
rect 313168 260383 313174 260395
rect 220490 260355 313174 260383
rect 220490 260343 220496 260355
rect 313168 260343 313174 260355
rect 313226 260343 313232 260395
rect 313264 260343 313270 260395
rect 313322 260383 313328 260395
rect 434512 260383 434518 260395
rect 313322 260355 434518 260383
rect 313322 260343 313328 260355
rect 434512 260343 434518 260355
rect 434570 260343 434576 260395
rect 213328 260269 213334 260321
rect 213386 260309 213392 260321
rect 309040 260309 309046 260321
rect 213386 260281 309046 260309
rect 213386 260269 213392 260281
rect 309040 260269 309046 260281
rect 309098 260269 309104 260321
rect 309424 260269 309430 260321
rect 309482 260309 309488 260321
rect 445264 260309 445270 260321
rect 309482 260281 445270 260309
rect 309482 260269 309488 260281
rect 445264 260269 445270 260281
rect 445322 260269 445328 260321
rect 269200 260195 269206 260247
rect 269258 260235 269264 260247
rect 388240 260235 388246 260247
rect 269258 260207 388246 260235
rect 269258 260195 269264 260207
rect 388240 260195 388246 260207
rect 388298 260195 388304 260247
rect 403696 260195 403702 260247
rect 403754 260235 403760 260247
rect 447664 260235 447670 260247
rect 403754 260207 447670 260235
rect 403754 260195 403760 260207
rect 447664 260195 447670 260207
rect 447722 260195 447728 260247
rect 156208 260121 156214 260173
rect 156266 260161 156272 260173
rect 305392 260161 305398 260173
rect 156266 260133 305398 260161
rect 156266 260121 156272 260133
rect 305392 260121 305398 260133
rect 305450 260121 305456 260173
rect 308368 260121 308374 260173
rect 308426 260161 308432 260173
rect 427408 260161 427414 260173
rect 308426 260133 427414 260161
rect 308426 260121 308432 260133
rect 427408 260121 427414 260133
rect 427466 260121 427472 260173
rect 431152 260121 431158 260173
rect 431210 260161 431216 260173
rect 443248 260161 443254 260173
rect 431210 260133 443254 260161
rect 431210 260121 431216 260133
rect 443248 260121 443254 260133
rect 443306 260121 443312 260173
rect 145552 260047 145558 260099
rect 145610 260087 145616 260099
rect 305296 260087 305302 260099
rect 145610 260059 305302 260087
rect 145610 260047 145616 260059
rect 305296 260047 305302 260059
rect 305354 260047 305360 260099
rect 307984 260047 307990 260099
rect 308042 260087 308048 260099
rect 420208 260087 420214 260099
rect 308042 260059 420214 260087
rect 308042 260047 308048 260059
rect 420208 260047 420214 260059
rect 420266 260047 420272 260099
rect 426352 260047 426358 260099
rect 426410 260087 426416 260099
rect 436048 260087 436054 260099
rect 426410 260059 436054 260087
rect 426410 260047 426416 260059
rect 436048 260047 436054 260059
rect 436106 260047 436112 260099
rect 307216 259973 307222 260025
rect 307274 260013 307280 260025
rect 307274 259985 399038 260013
rect 307274 259973 307280 259985
rect 307600 259899 307606 259951
rect 307658 259939 307664 259951
rect 399010 259939 399038 259985
rect 405520 259973 405526 260025
rect 405578 260013 405584 260025
rect 424912 260013 424918 260025
rect 405578 259985 424918 260013
rect 405578 259973 405584 259985
rect 424912 259973 424918 259985
rect 424970 259973 424976 260025
rect 432784 259973 432790 260025
rect 432842 260013 432848 260025
rect 443152 260013 443158 260025
rect 432842 259985 443158 260013
rect 432842 259973 432848 259985
rect 443152 259973 443158 259985
rect 443210 259973 443216 260025
rect 406000 259939 406006 259951
rect 307658 259911 398942 259939
rect 399010 259911 406006 259939
rect 307658 259899 307664 259911
rect 306928 259825 306934 259877
rect 306986 259865 306992 259877
rect 398914 259865 398942 259911
rect 406000 259899 406006 259911
rect 406058 259899 406064 259951
rect 306986 259837 395582 259865
rect 398914 259837 402494 259865
rect 306986 259825 306992 259837
rect 306544 259751 306550 259803
rect 306602 259791 306608 259803
rect 395248 259791 395254 259803
rect 306602 259763 395254 259791
rect 306602 259751 306608 259763
rect 395248 259751 395254 259763
rect 395306 259751 395312 259803
rect 306160 259677 306166 259729
rect 306218 259717 306224 259729
rect 388144 259717 388150 259729
rect 306218 259689 388150 259717
rect 306218 259677 306224 259689
rect 388144 259677 388150 259689
rect 388202 259677 388208 259729
rect 395554 259717 395582 259837
rect 402352 259717 402358 259729
rect 395554 259689 402358 259717
rect 402352 259677 402358 259689
rect 402410 259677 402416 259729
rect 402466 259717 402494 259837
rect 408784 259825 408790 259877
rect 408842 259865 408848 259877
rect 427888 259865 427894 259877
rect 408842 259837 427894 259865
rect 408842 259825 408848 259837
rect 427888 259825 427894 259837
rect 427946 259825 427952 259877
rect 406288 259751 406294 259803
rect 406346 259791 406352 259803
rect 425680 259791 425686 259803
rect 406346 259763 425686 259791
rect 406346 259751 406352 259763
rect 425680 259751 425686 259763
rect 425738 259751 425744 259803
rect 413104 259717 413110 259729
rect 402466 259689 413110 259717
rect 413104 259677 413110 259689
rect 413162 259677 413168 259729
rect 304336 259603 304342 259655
rect 304394 259643 304400 259655
rect 355984 259643 355990 259655
rect 304394 259615 355990 259643
rect 304394 259603 304400 259615
rect 355984 259603 355990 259615
rect 356042 259603 356048 259655
rect 356560 259603 356566 259655
rect 356618 259643 356624 259655
rect 430000 259643 430006 259655
rect 356618 259615 430006 259643
rect 356618 259603 356624 259615
rect 430000 259603 430006 259615
rect 430058 259603 430064 259655
rect 286000 259529 286006 259581
rect 286058 259569 286064 259581
rect 354256 259569 354262 259581
rect 286058 259541 354262 259569
rect 286058 259529 286064 259541
rect 354256 259529 354262 259541
rect 354314 259529 354320 259581
rect 354448 259529 354454 259581
rect 354506 259569 354512 259581
rect 407152 259569 407158 259581
rect 354506 259541 407158 259569
rect 354506 259529 354512 259541
rect 407152 259529 407158 259541
rect 407210 259529 407216 259581
rect 286672 259455 286678 259507
rect 286730 259495 286736 259507
rect 369424 259495 369430 259507
rect 286730 259467 369430 259495
rect 286730 259455 286736 259467
rect 369424 259455 369430 259467
rect 369482 259455 369488 259507
rect 377872 259455 377878 259507
rect 377930 259495 377936 259507
rect 590320 259495 590326 259507
rect 377930 259467 590326 259495
rect 377930 259455 377936 259467
rect 590320 259455 590326 259467
rect 590378 259455 590384 259507
rect 286096 259381 286102 259433
rect 286154 259421 286160 259433
rect 370864 259421 370870 259433
rect 286154 259393 370870 259421
rect 286154 259381 286160 259393
rect 370864 259381 370870 259393
rect 370922 259381 370928 259433
rect 378352 259381 378358 259433
rect 378410 259421 378416 259433
rect 378410 259393 379358 259421
rect 378410 259381 378416 259393
rect 282448 259307 282454 259359
rect 282506 259347 282512 259359
rect 369040 259347 369046 259359
rect 282506 259319 369046 259347
rect 282506 259307 282512 259319
rect 369040 259307 369046 259319
rect 369098 259307 369104 259359
rect 378256 259307 378262 259359
rect 378314 259347 378320 259359
rect 379120 259347 379126 259359
rect 378314 259319 379126 259347
rect 378314 259307 378320 259319
rect 379120 259307 379126 259319
rect 379178 259307 379184 259359
rect 379330 259347 379358 259393
rect 383632 259381 383638 259433
rect 383690 259421 383696 259433
rect 385264 259421 385270 259433
rect 383690 259393 385270 259421
rect 383690 259381 383696 259393
rect 385264 259381 385270 259393
rect 385322 259381 385328 259433
rect 384880 259347 384886 259359
rect 379330 259319 384886 259347
rect 384880 259307 384886 259319
rect 384938 259307 384944 259359
rect 389584 259307 389590 259359
rect 389642 259347 389648 259359
rect 390064 259347 390070 259359
rect 389642 259319 390070 259347
rect 389642 259307 389648 259319
rect 390064 259307 390070 259319
rect 390122 259307 390128 259359
rect 284560 259233 284566 259285
rect 284618 259273 284624 259285
rect 425008 259273 425014 259285
rect 284618 259245 425014 259273
rect 284618 259233 284624 259245
rect 425008 259233 425014 259245
rect 425066 259233 425072 259285
rect 305296 259159 305302 259211
rect 305354 259199 305360 259211
rect 429808 259199 429814 259211
rect 305354 259171 429814 259199
rect 305354 259159 305360 259171
rect 429808 259159 429814 259171
rect 429866 259159 429872 259211
rect 433840 259199 433846 259211
rect 429922 259171 433846 259199
rect 305392 259085 305398 259137
rect 305450 259125 305456 259137
rect 429712 259125 429718 259137
rect 305450 259097 429718 259125
rect 305450 259085 305456 259097
rect 429712 259085 429718 259097
rect 429770 259085 429776 259137
rect 302416 259011 302422 259063
rect 302474 259051 302480 259063
rect 429922 259051 429950 259171
rect 433840 259159 433846 259171
rect 433898 259159 433904 259211
rect 440560 259159 440566 259211
rect 440618 259199 440624 259211
rect 445648 259199 445654 259211
rect 440618 259171 445654 259199
rect 440618 259159 440624 259171
rect 445648 259159 445654 259171
rect 445706 259159 445712 259211
rect 430096 259085 430102 259137
rect 430154 259125 430160 259137
rect 447856 259125 447862 259137
rect 430154 259097 447862 259125
rect 430154 259085 430160 259097
rect 447856 259085 447862 259097
rect 447914 259085 447920 259137
rect 447952 259085 447958 259137
rect 448010 259125 448016 259137
rect 451888 259125 451894 259137
rect 448010 259097 451894 259125
rect 448010 259085 448016 259097
rect 451888 259085 451894 259097
rect 451946 259085 451952 259137
rect 302474 259023 429950 259051
rect 302474 259011 302480 259023
rect 435952 259011 435958 259063
rect 436010 259051 436016 259063
rect 449392 259051 449398 259063
rect 436010 259023 449398 259051
rect 436010 259011 436016 259023
rect 449392 259011 449398 259023
rect 449450 259011 449456 259063
rect 305488 258937 305494 258989
rect 305546 258977 305552 258989
rect 430480 258977 430486 258989
rect 305546 258949 430486 258977
rect 305546 258937 305552 258949
rect 430480 258937 430486 258949
rect 430538 258937 430544 258989
rect 433456 258937 433462 258989
rect 433514 258977 433520 258989
rect 447952 258977 447958 258989
rect 433514 258949 447958 258977
rect 433514 258937 433520 258949
rect 447952 258937 447958 258949
rect 448010 258937 448016 258989
rect 452944 258977 452950 258989
rect 448162 258949 452950 258977
rect 302512 258863 302518 258915
rect 302570 258903 302576 258915
rect 432688 258903 432694 258915
rect 302570 258875 432694 258903
rect 302570 258863 302576 258875
rect 432688 258863 432694 258875
rect 432746 258863 432752 258915
rect 288880 258789 288886 258841
rect 288938 258829 288944 258841
rect 433456 258829 433462 258841
rect 288938 258801 433462 258829
rect 288938 258789 288944 258801
rect 433456 258789 433462 258801
rect 433514 258789 433520 258841
rect 443248 258789 443254 258841
rect 443306 258829 443312 258841
rect 448162 258829 448190 258949
rect 452944 258937 452950 258949
rect 453002 258937 453008 258989
rect 443306 258801 448190 258829
rect 443306 258789 443312 258801
rect 282256 258715 282262 258767
rect 282314 258755 282320 258767
rect 418768 258755 418774 258767
rect 282314 258727 418774 258755
rect 282314 258715 282320 258727
rect 418768 258715 418774 258727
rect 418826 258715 418832 258767
rect 418864 258715 418870 258767
rect 418922 258755 418928 258767
rect 443056 258755 443062 258767
rect 418922 258727 443062 258755
rect 418922 258715 418928 258727
rect 443056 258715 443062 258727
rect 443114 258715 443120 258767
rect 443152 258715 443158 258767
rect 443210 258755 443216 258767
rect 451120 258755 451126 258767
rect 443210 258727 451126 258755
rect 443210 258715 443216 258727
rect 451120 258715 451126 258727
rect 451178 258715 451184 258767
rect 277840 258641 277846 258693
rect 277898 258681 277904 258693
rect 439696 258681 439702 258693
rect 277898 258653 439702 258681
rect 277898 258641 277904 258653
rect 439696 258641 439702 258653
rect 439754 258641 439760 258693
rect 277936 258567 277942 258619
rect 277994 258607 278000 258619
rect 430096 258607 430102 258619
rect 277994 258579 430102 258607
rect 277994 258567 278000 258579
rect 430096 258567 430102 258579
rect 430154 258567 430160 258619
rect 430192 258567 430198 258619
rect 430250 258607 430256 258619
rect 447088 258607 447094 258619
rect 430250 258579 447094 258607
rect 430250 258567 430256 258579
rect 447088 258567 447094 258579
rect 447146 258567 447152 258619
rect 234064 258493 234070 258545
rect 234122 258533 234128 258545
rect 445264 258533 445270 258545
rect 234122 258505 445270 258533
rect 234122 258493 234128 258505
rect 445264 258493 445270 258505
rect 445322 258493 445328 258545
rect 233200 258419 233206 258471
rect 233258 258459 233264 258471
rect 444496 258459 444502 258471
rect 233258 258431 444502 258459
rect 233258 258419 233264 258431
rect 444496 258419 444502 258431
rect 444554 258419 444560 258471
rect 201616 258345 201622 258397
rect 201674 258385 201680 258397
rect 446704 258385 446710 258397
rect 201674 258357 446710 258385
rect 201674 258345 201680 258357
rect 446704 258345 446710 258357
rect 446762 258345 446768 258397
rect 161008 258271 161014 258323
rect 161066 258311 161072 258323
rect 443728 258311 443734 258323
rect 161066 258283 443734 258311
rect 161066 258271 161072 258283
rect 443728 258271 443734 258283
rect 443786 258271 443792 258323
rect 153808 258197 153814 258249
rect 153866 258237 153872 258249
rect 418864 258237 418870 258249
rect 153866 258209 418870 258237
rect 153866 258197 153872 258209
rect 418864 258197 418870 258209
rect 418922 258197 418928 258249
rect 441520 258237 441526 258249
rect 418978 258209 441526 258237
rect 143152 258123 143158 258175
rect 143210 258163 143216 258175
rect 418978 258163 419006 258209
rect 441520 258197 441526 258209
rect 441578 258197 441584 258249
rect 143210 258135 419006 258163
rect 143210 258123 143216 258135
rect 423376 258123 423382 258175
rect 423434 258163 423440 258175
rect 427984 258163 427990 258175
rect 423434 258135 427990 258163
rect 423434 258123 423440 258135
rect 427984 258123 427990 258135
rect 428042 258123 428048 258175
rect 428176 258123 428182 258175
rect 428234 258163 428240 258175
rect 441232 258163 441238 258175
rect 428234 258135 441238 258163
rect 428234 258123 428240 258135
rect 441232 258123 441238 258135
rect 441290 258123 441296 258175
rect 83632 258049 83638 258101
rect 83690 258089 83696 258101
rect 96304 258089 96310 258101
rect 83690 258061 96310 258089
rect 83690 258049 83696 258061
rect 96304 258049 96310 258061
rect 96362 258049 96368 258101
rect 118096 258049 118102 258101
rect 118154 258089 118160 258101
rect 438832 258089 438838 258101
rect 118154 258061 438838 258089
rect 118154 258049 118160 258061
rect 438832 258049 438838 258061
rect 438890 258049 438896 258101
rect 106192 257975 106198 258027
rect 106250 258015 106256 258027
rect 437104 258015 437110 258027
rect 106250 257987 437110 258015
rect 106250 257975 106256 257987
rect 437104 257975 437110 257987
rect 437162 257975 437168 258027
rect 437200 257975 437206 258027
rect 437258 258015 437264 258027
rect 450352 258015 450358 258027
rect 437258 257987 450358 258015
rect 437258 257975 437264 257987
rect 450352 257975 450358 257987
rect 450410 257975 450416 258027
rect 99184 257901 99190 257953
rect 99242 257941 99248 257953
rect 436432 257941 436438 257953
rect 99242 257913 436438 257941
rect 99242 257901 99248 257913
rect 436432 257901 436438 257913
rect 436490 257901 436496 257953
rect 110992 257827 110998 257879
rect 111050 257867 111056 257879
rect 449584 257867 449590 257879
rect 111050 257839 449590 257867
rect 111050 257827 111056 257839
rect 449584 257827 449590 257839
rect 449642 257827 449648 257879
rect 103888 257753 103894 257805
rect 103946 257793 103952 257805
rect 448912 257793 448918 257805
rect 103946 257765 448918 257793
rect 103946 257753 103952 257765
rect 448912 257753 448918 257765
rect 448970 257753 448976 257805
rect 455440 257753 455446 257805
rect 455498 257793 455504 257805
rect 456784 257793 456790 257805
rect 455498 257765 456790 257793
rect 455498 257753 455504 257765
rect 456784 257753 456790 257765
rect 456842 257753 456848 257805
rect 460816 257753 460822 257805
rect 460874 257793 460880 257805
rect 462832 257793 462838 257805
rect 460874 257765 462838 257793
rect 460874 257753 460880 257765
rect 462832 257753 462838 257765
rect 462890 257753 462896 257805
rect 469456 257753 469462 257805
rect 469514 257793 469520 257805
rect 471088 257793 471094 257805
rect 469514 257765 471094 257793
rect 469514 257753 469520 257765
rect 471088 257753 471094 257765
rect 471146 257753 471152 257805
rect 480976 257753 480982 257805
rect 481034 257793 481040 257805
rect 482992 257793 482998 257805
rect 481034 257765 482998 257793
rect 481034 257753 481040 257765
rect 482992 257753 482998 257765
rect 483050 257753 483056 257805
rect 486832 257753 486838 257805
rect 486890 257793 486896 257805
rect 488944 257793 488950 257805
rect 486890 257765 488950 257793
rect 486890 257753 486896 257765
rect 488944 257753 488950 257765
rect 489002 257753 489008 257805
rect 492688 257753 492694 257805
rect 492746 257793 492752 257805
rect 494800 257793 494806 257805
rect 492746 257765 494806 257793
rect 492746 257753 492752 257765
rect 494800 257753 494806 257765
rect 494858 257753 494864 257805
rect 495376 257753 495382 257805
rect 495434 257793 495440 257805
rect 497296 257793 497302 257805
rect 495434 257765 497302 257793
rect 495434 257753 495440 257765
rect 497296 257753 497302 257765
rect 497354 257753 497360 257805
rect 501232 257753 501238 257805
rect 501290 257793 501296 257805
rect 503152 257793 503158 257805
rect 501290 257765 503158 257793
rect 501290 257753 501296 257765
rect 503152 257753 503158 257765
rect 503210 257753 503216 257805
rect 507088 257753 507094 257805
rect 507146 257793 507152 257805
rect 509200 257793 509206 257805
rect 507146 257765 509206 257793
rect 507146 257753 507152 257765
rect 509200 257753 509206 257765
rect 509258 257753 509264 257805
rect 509776 257753 509782 257805
rect 509834 257793 509840 257805
rect 511600 257793 511606 257805
rect 509834 257765 511606 257793
rect 509834 257753 509840 257765
rect 511600 257753 511606 257765
rect 511658 257753 511664 257805
rect 512848 257753 512854 257805
rect 512906 257793 512912 257805
rect 514000 257793 514006 257805
rect 512906 257765 514006 257793
rect 512906 257753 512912 257765
rect 514000 257753 514006 257765
rect 514058 257753 514064 257805
rect 527056 257753 527062 257805
rect 527114 257793 527120 257805
rect 528208 257793 528214 257805
rect 527114 257765 528214 257793
rect 527114 257753 527120 257765
rect 528208 257753 528214 257765
rect 528266 257753 528272 257805
rect 533008 257753 533014 257805
rect 533066 257793 533072 257805
rect 535312 257793 535318 257805
rect 533066 257765 535318 257793
rect 533066 257753 533072 257765
rect 535312 257753 535318 257765
rect 535370 257753 535376 257805
rect 541648 257753 541654 257805
rect 541706 257793 541712 257805
rect 543664 257793 543670 257805
rect 541706 257765 543670 257793
rect 541706 257753 541712 257765
rect 543664 257753 543670 257765
rect 543722 257753 543728 257805
rect 282256 257679 282262 257731
rect 282314 257719 282320 257731
rect 284368 257719 284374 257731
rect 282314 257691 284374 257719
rect 282314 257679 282320 257691
rect 284368 257679 284374 257691
rect 284426 257679 284432 257731
rect 305584 257679 305590 257731
rect 305642 257719 305648 257731
rect 429040 257719 429046 257731
rect 305642 257691 429046 257719
rect 305642 257679 305648 257691
rect 429040 257679 429046 257691
rect 429098 257679 429104 257731
rect 430096 257679 430102 257731
rect 430154 257719 430160 257731
rect 445936 257719 445942 257731
rect 430154 257691 445942 257719
rect 430154 257679 430160 257691
rect 445936 257679 445942 257691
rect 445994 257679 446000 257731
rect 512656 257679 512662 257731
rect 512714 257719 512720 257731
rect 515152 257719 515158 257731
rect 512714 257691 515158 257719
rect 512714 257679 512720 257691
rect 515152 257679 515158 257691
rect 515210 257679 515216 257731
rect 527152 257679 527158 257731
rect 527210 257719 527216 257731
rect 529456 257719 529462 257731
rect 527210 257691 529462 257719
rect 527210 257679 527216 257691
rect 529456 257679 529462 257691
rect 529514 257679 529520 257731
rect 309136 257605 309142 257657
rect 309194 257645 309200 257657
rect 428272 257645 428278 257657
rect 309194 257617 428278 257645
rect 309194 257605 309200 257617
rect 428272 257605 428278 257617
rect 428330 257605 428336 257657
rect 428464 257605 428470 257657
rect 428522 257645 428528 257657
rect 446320 257645 446326 257657
rect 428522 257617 446326 257645
rect 428522 257605 428528 257617
rect 446320 257605 446326 257617
rect 446378 257605 446384 257657
rect 427600 257571 427606 257583
rect 330658 257543 427606 257571
rect 325456 257235 325462 257287
rect 325514 257275 325520 257287
rect 330658 257275 330686 257543
rect 427600 257531 427606 257543
rect 427658 257531 427664 257583
rect 430288 257531 430294 257583
rect 430346 257571 430352 257583
rect 448528 257571 448534 257583
rect 430346 257543 448534 257571
rect 430346 257531 430352 257543
rect 448528 257531 448534 257543
rect 448586 257531 448592 257583
rect 331888 257457 331894 257509
rect 331946 257497 331952 257509
rect 333616 257497 333622 257509
rect 331946 257469 333622 257497
rect 331946 257457 331952 257469
rect 333616 257457 333622 257469
rect 333674 257457 333680 257509
rect 334864 257457 334870 257509
rect 334922 257497 334928 257509
rect 339664 257497 339670 257509
rect 334922 257469 339670 257497
rect 334922 257457 334928 257469
rect 339664 257457 339670 257469
rect 339722 257457 339728 257509
rect 426832 257497 426838 257509
rect 339778 257469 426838 257497
rect 331120 257383 331126 257435
rect 331178 257423 331184 257435
rect 339778 257423 339806 257469
rect 426832 257457 426838 257469
rect 426890 257457 426896 257509
rect 426928 257457 426934 257509
rect 426986 257497 426992 257509
rect 426986 257469 427358 257497
rect 426986 257457 426992 257469
rect 427216 257423 427222 257435
rect 331178 257395 339806 257423
rect 339874 257395 427222 257423
rect 331178 257383 331184 257395
rect 330736 257309 330742 257361
rect 330794 257349 330800 257361
rect 339874 257349 339902 257395
rect 427216 257383 427222 257395
rect 427274 257383 427280 257435
rect 427330 257423 427358 257469
rect 427888 257457 427894 257509
rect 427946 257497 427952 257509
rect 444112 257497 444118 257509
rect 427946 257469 444118 257497
rect 427946 257457 427952 257469
rect 444112 257457 444118 257469
rect 444170 257457 444176 257509
rect 444880 257423 444886 257435
rect 427330 257395 444886 257423
rect 444880 257383 444886 257395
rect 444938 257383 444944 257435
rect 330794 257321 339902 257349
rect 330794 257309 330800 257321
rect 351088 257309 351094 257361
rect 351146 257349 351152 257361
rect 357424 257349 357430 257361
rect 351146 257321 357430 257349
rect 351146 257309 351152 257321
rect 357424 257309 357430 257321
rect 357482 257309 357488 257361
rect 358480 257309 358486 257361
rect 358538 257349 358544 257361
rect 426448 257349 426454 257361
rect 358538 257321 426454 257349
rect 358538 257309 358544 257321
rect 426448 257309 426454 257321
rect 426506 257309 426512 257361
rect 325514 257247 330686 257275
rect 325514 257235 325520 257247
rect 333520 257235 333526 257287
rect 333578 257275 333584 257287
rect 394480 257275 394486 257287
rect 333578 257247 394486 257275
rect 333578 257235 333584 257247
rect 394480 257235 394486 257247
rect 394538 257235 394544 257287
rect 401104 257235 401110 257287
rect 401162 257275 401168 257287
rect 404752 257275 404758 257287
rect 401162 257247 404758 257275
rect 401162 257235 401168 257247
rect 404752 257235 404758 257247
rect 404810 257235 404816 257287
rect 406960 257235 406966 257287
rect 407018 257275 407024 257287
rect 408688 257275 408694 257287
rect 407018 257247 408694 257275
rect 407018 257235 407024 257247
rect 408688 257235 408694 257247
rect 408746 257235 408752 257287
rect 409168 257235 409174 257287
rect 409226 257275 409232 257287
rect 423664 257275 423670 257287
rect 409226 257247 423670 257275
rect 409226 257235 409232 257247
rect 423664 257235 423670 257247
rect 423722 257235 423728 257287
rect 425968 257235 425974 257287
rect 426026 257275 426032 257287
rect 438928 257275 438934 257287
rect 426026 257247 438934 257275
rect 426026 257235 426032 257247
rect 438928 257235 438934 257247
rect 438986 257235 438992 257287
rect 333136 257161 333142 257213
rect 333194 257201 333200 257213
rect 393712 257201 393718 257213
rect 333194 257173 393718 257201
rect 333194 257161 333200 257173
rect 393712 257161 393718 257173
rect 393770 257161 393776 257213
rect 427312 257161 427318 257213
rect 427370 257201 427376 257213
rect 442672 257201 442678 257213
rect 427370 257173 442678 257201
rect 427370 257161 427376 257173
rect 442672 257161 442678 257173
rect 442730 257161 442736 257213
rect 331216 257087 331222 257139
rect 331274 257127 331280 257139
rect 337840 257127 337846 257139
rect 331274 257099 337846 257127
rect 331274 257087 331280 257099
rect 337840 257087 337846 257099
rect 337898 257087 337904 257139
rect 350704 257087 350710 257139
rect 350762 257127 350768 257139
rect 353584 257127 353590 257139
rect 350762 257099 353590 257127
rect 350762 257087 350768 257099
rect 353584 257087 353590 257099
rect 353642 257087 353648 257139
rect 360016 257087 360022 257139
rect 360074 257127 360080 257139
rect 396304 257127 396310 257139
rect 360074 257099 396310 257127
rect 360074 257087 360080 257099
rect 396304 257087 396310 257099
rect 396362 257087 396368 257139
rect 418768 257087 418774 257139
rect 418826 257127 418832 257139
rect 440848 257127 440854 257139
rect 418826 257099 440854 257127
rect 418826 257087 418832 257099
rect 440848 257087 440854 257099
rect 440906 257087 440912 257139
rect 346576 257013 346582 257065
rect 346634 257053 346640 257065
rect 349936 257053 349942 257065
rect 346634 257025 349942 257053
rect 346634 257013 346640 257025
rect 349936 257013 349942 257025
rect 349994 257013 350000 257065
rect 378736 257013 378742 257065
rect 378794 257053 378800 257065
rect 379216 257053 379222 257065
rect 378794 257025 379222 257053
rect 378794 257013 378800 257025
rect 379216 257013 379222 257025
rect 379274 257013 379280 257065
rect 383056 257013 383062 257065
rect 383114 257053 383120 257065
rect 393040 257053 393046 257065
rect 383114 257025 393046 257053
rect 383114 257013 383120 257025
rect 393040 257013 393046 257025
rect 393098 257013 393104 257065
rect 423184 257013 423190 257065
rect 423242 257053 423248 257065
rect 440464 257053 440470 257065
rect 423242 257025 440470 257053
rect 423242 257013 423248 257025
rect 440464 257013 440470 257025
rect 440522 257013 440528 257065
rect 342928 256939 342934 256991
rect 342986 256979 342992 256991
rect 349552 256979 349558 256991
rect 342986 256951 349558 256979
rect 342986 256939 342992 256951
rect 349552 256939 349558 256951
rect 349610 256939 349616 256991
rect 351760 256939 351766 256991
rect 351818 256979 351824 256991
rect 364336 256979 364342 256991
rect 351818 256951 364342 256979
rect 351818 256939 351824 256951
rect 364336 256939 364342 256951
rect 364394 256939 364400 256991
rect 368656 256939 368662 256991
rect 368714 256979 368720 256991
rect 368714 256951 378686 256979
rect 368714 256939 368720 256951
rect 322288 256865 322294 256917
rect 322346 256905 322352 256917
rect 327184 256905 327190 256917
rect 322346 256877 327190 256905
rect 322346 256865 322352 256877
rect 327184 256865 327190 256877
rect 327242 256865 327248 256917
rect 330928 256865 330934 256917
rect 330986 256905 330992 256917
rect 330986 256877 342014 256905
rect 330986 256865 330992 256877
rect 282544 256791 282550 256843
rect 282602 256831 282608 256843
rect 325648 256831 325654 256843
rect 282602 256803 325654 256831
rect 282602 256791 282608 256803
rect 325648 256791 325654 256803
rect 325706 256791 325712 256843
rect 329008 256791 329014 256843
rect 329066 256831 329072 256843
rect 341872 256831 341878 256843
rect 329066 256803 341878 256831
rect 329066 256791 329072 256803
rect 341872 256791 341878 256803
rect 341930 256791 341936 256843
rect 341986 256831 342014 256877
rect 366832 256865 366838 256917
rect 366890 256905 366896 256917
rect 378448 256905 378454 256917
rect 366890 256877 378454 256905
rect 366890 256865 366896 256877
rect 378448 256865 378454 256877
rect 378506 256865 378512 256917
rect 358480 256831 358486 256843
rect 341986 256803 358486 256831
rect 358480 256791 358486 256803
rect 358538 256791 358544 256843
rect 365584 256791 365590 256843
rect 365642 256831 365648 256843
rect 365642 256803 367742 256831
rect 365642 256791 365648 256803
rect 285904 256717 285910 256769
rect 285962 256757 285968 256769
rect 366832 256757 366838 256769
rect 285962 256729 366838 256757
rect 285962 256717 285968 256729
rect 366832 256717 366838 256729
rect 366890 256717 366896 256769
rect 367714 256757 367742 256803
rect 367792 256791 367798 256843
rect 367850 256831 367856 256843
rect 378544 256831 378550 256843
rect 367850 256803 378550 256831
rect 367850 256791 367856 256803
rect 378544 256791 378550 256803
rect 378602 256791 378608 256843
rect 378658 256831 378686 256951
rect 378832 256939 378838 256991
rect 378890 256979 378896 256991
rect 388720 256979 388726 256991
rect 378890 256951 388726 256979
rect 378890 256939 378896 256951
rect 388720 256939 388726 256951
rect 388778 256939 388784 256991
rect 423472 256939 423478 256991
rect 423530 256979 423536 256991
rect 428656 256979 428662 256991
rect 423530 256951 428662 256979
rect 423530 256939 423536 256951
rect 428656 256939 428662 256951
rect 428714 256939 428720 256991
rect 428944 256939 428950 256991
rect 429002 256979 429008 256991
rect 441904 256979 441910 256991
rect 429002 256951 441910 256979
rect 429002 256939 429008 256951
rect 441904 256939 441910 256951
rect 441962 256939 441968 256991
rect 425776 256865 425782 256917
rect 425834 256905 425840 256917
rect 428176 256905 428182 256917
rect 425834 256877 428182 256905
rect 425834 256865 425840 256877
rect 428176 256865 428182 256877
rect 428234 256865 428240 256917
rect 429712 256865 429718 256917
rect 429770 256905 429776 256917
rect 431248 256905 431254 256917
rect 429770 256877 431254 256905
rect 429770 256865 429776 256877
rect 431248 256865 431254 256877
rect 431306 256865 431312 256917
rect 395920 256831 395926 256843
rect 378658 256803 395926 256831
rect 395920 256791 395926 256803
rect 395978 256791 395984 256843
rect 425872 256791 425878 256843
rect 425930 256831 425936 256843
rect 437872 256831 437878 256843
rect 425930 256803 437878 256831
rect 425930 256791 425936 256803
rect 437872 256791 437878 256803
rect 437930 256791 437936 256843
rect 368368 256757 368374 256769
rect 367714 256729 368374 256757
rect 368368 256717 368374 256729
rect 368426 256717 368432 256769
rect 368464 256717 368470 256769
rect 368522 256757 368528 256769
rect 383152 256757 383158 256769
rect 368522 256729 383158 256757
rect 368522 256717 368528 256729
rect 383152 256717 383158 256729
rect 383210 256717 383216 256769
rect 383266 256729 383582 256757
rect 286480 256643 286486 256695
rect 286538 256683 286544 256695
rect 365872 256683 365878 256695
rect 286538 256655 365878 256683
rect 286538 256643 286544 256655
rect 365872 256643 365878 256655
rect 365930 256643 365936 256695
rect 367120 256643 367126 256695
rect 367178 256683 367184 256695
rect 383266 256683 383294 256729
rect 367178 256655 383294 256683
rect 383554 256683 383582 256729
rect 391600 256717 391606 256769
rect 391658 256757 391664 256769
rect 452272 256757 452278 256769
rect 391658 256729 452278 256757
rect 391658 256717 391664 256729
rect 452272 256717 452278 256729
rect 452330 256717 452336 256769
rect 438256 256683 438262 256695
rect 383554 256655 438262 256683
rect 367178 256643 367184 256655
rect 438256 256643 438262 256655
rect 438314 256643 438320 256695
rect 285808 256569 285814 256621
rect 285866 256609 285872 256621
rect 365584 256609 365590 256621
rect 285866 256581 365590 256609
rect 285866 256569 285872 256581
rect 365584 256569 365590 256581
rect 365642 256569 365648 256621
rect 367504 256609 367510 256621
rect 365698 256581 367510 256609
rect 285232 256495 285238 256547
rect 285290 256535 285296 256547
rect 365698 256535 365726 256581
rect 367504 256569 367510 256581
rect 367562 256569 367568 256621
rect 367600 256569 367606 256621
rect 367658 256609 367664 256621
rect 442288 256609 442294 256621
rect 367658 256581 442294 256609
rect 367658 256569 367664 256581
rect 442288 256569 442294 256581
rect 442346 256569 442352 256621
rect 383632 256535 383638 256547
rect 285290 256507 301022 256535
rect 285290 256495 285296 256507
rect 285136 256421 285142 256473
rect 285194 256461 285200 256473
rect 300994 256461 301022 256507
rect 310690 256507 365726 256535
rect 378466 256507 383638 256535
rect 310690 256461 310718 256507
rect 369808 256461 369814 256473
rect 285194 256433 300926 256461
rect 300994 256433 310718 256461
rect 310786 256433 369814 256461
rect 285194 256421 285200 256433
rect 283600 256347 283606 256399
rect 283658 256387 283664 256399
rect 300784 256387 300790 256399
rect 283658 256359 300790 256387
rect 283658 256347 283664 256359
rect 300784 256347 300790 256359
rect 300842 256347 300848 256399
rect 300898 256387 300926 256433
rect 310786 256387 310814 256433
rect 369808 256421 369814 256433
rect 369866 256421 369872 256473
rect 371440 256421 371446 256473
rect 371498 256461 371504 256473
rect 378466 256461 378494 256507
rect 383632 256495 383638 256507
rect 383690 256495 383696 256547
rect 383728 256495 383734 256547
rect 383786 256535 383792 256547
rect 451504 256535 451510 256547
rect 383786 256507 451510 256535
rect 383786 256495 383792 256507
rect 451504 256495 451510 256507
rect 451562 256495 451568 256547
rect 371498 256433 378494 256461
rect 371498 256421 371504 256433
rect 378544 256421 378550 256473
rect 378602 256461 378608 256473
rect 383056 256461 383062 256473
rect 378602 256433 383062 256461
rect 378602 256421 378608 256433
rect 383056 256421 383062 256433
rect 383114 256421 383120 256473
rect 393040 256421 393046 256473
rect 393098 256461 393104 256473
rect 450064 256461 450070 256473
rect 393098 256433 450070 256461
rect 393098 256421 393104 256433
rect 450064 256421 450070 256433
rect 450122 256421 450128 256473
rect 300898 256359 310814 256387
rect 310864 256347 310870 256399
rect 310922 256387 310928 256399
rect 370192 256387 370198 256399
rect 310922 256359 370198 256387
rect 310922 256347 310928 256359
rect 370192 256347 370198 256359
rect 370250 256347 370256 256399
rect 370288 256347 370294 256399
rect 370346 256387 370352 256399
rect 450736 256387 450742 256399
rect 370346 256359 450742 256387
rect 370346 256347 370352 256359
rect 450736 256347 450742 256359
rect 450794 256347 450800 256399
rect 640720 256347 640726 256399
rect 640778 256387 640784 256399
rect 679696 256387 679702 256399
rect 640778 256359 679702 256387
rect 640778 256347 640784 256359
rect 679696 256347 679702 256359
rect 679754 256347 679760 256399
rect 310960 256273 310966 256325
rect 311018 256313 311024 256325
rect 322384 256313 322390 256325
rect 311018 256285 322390 256313
rect 311018 256273 311024 256285
rect 322384 256273 322390 256285
rect 322442 256273 322448 256325
rect 322576 256273 322582 256325
rect 322634 256313 322640 256325
rect 637648 256313 637654 256325
rect 322634 256285 637654 256313
rect 322634 256273 322640 256285
rect 637648 256273 637654 256285
rect 637706 256273 637712 256325
rect 288880 256199 288886 256251
rect 288938 256239 288944 256251
rect 322480 256239 322486 256251
rect 288938 256211 322486 256239
rect 288938 256199 288944 256211
rect 322480 256199 322486 256211
rect 322538 256199 322544 256251
rect 322672 256199 322678 256251
rect 322730 256239 322736 256251
rect 630736 256239 630742 256251
rect 322730 256211 630742 256239
rect 322730 256199 322736 256211
rect 630736 256199 630742 256211
rect 630794 256199 630800 256251
rect 300400 256125 300406 256177
rect 300458 256165 300464 256177
rect 310384 256165 310390 256177
rect 300458 256137 310390 256165
rect 300458 256125 300464 256137
rect 310384 256125 310390 256137
rect 310442 256125 310448 256177
rect 422416 256165 422422 256177
rect 310498 256137 422422 256165
rect 282640 256051 282646 256103
rect 282698 256091 282704 256103
rect 293104 256091 293110 256103
rect 282698 256063 293110 256091
rect 282698 256051 282704 256063
rect 293104 256051 293110 256063
rect 293162 256051 293168 256103
rect 293200 256051 293206 256103
rect 293258 256091 293264 256103
rect 310498 256091 310526 256137
rect 422416 256125 422422 256137
rect 422474 256125 422480 256177
rect 495280 256125 495286 256177
rect 495338 256165 495344 256177
rect 508432 256165 508438 256177
rect 495338 256137 508438 256165
rect 495338 256125 495344 256137
rect 508432 256125 508438 256137
rect 508490 256125 508496 256177
rect 293258 256063 310526 256091
rect 293258 256051 293264 256063
rect 310576 256051 310582 256103
rect 310634 256091 310640 256103
rect 362800 256091 362806 256103
rect 310634 256063 362806 256091
rect 310634 256051 310640 256063
rect 362800 256051 362806 256063
rect 362858 256051 362864 256103
rect 285328 255977 285334 256029
rect 285386 256017 285392 256029
rect 363184 256017 363190 256029
rect 285386 255989 363190 256017
rect 285386 255977 285392 255989
rect 363184 255977 363190 255989
rect 363242 255977 363248 256029
rect 259312 255903 259318 255955
rect 259370 255943 259376 255955
rect 259370 255915 283742 255943
rect 259370 255903 259376 255915
rect 141136 255829 141142 255881
rect 141194 255869 141200 255881
rect 141194 255841 151262 255869
rect 141194 255829 141200 255841
rect 80656 255721 80662 255733
rect 80578 255693 80662 255721
rect 60592 255533 60598 255585
rect 60650 255573 60656 255585
rect 80578 255573 80606 255693
rect 80656 255681 80662 255693
rect 80714 255681 80720 255733
rect 106672 255681 106678 255733
rect 106730 255721 106736 255733
rect 118096 255721 118102 255733
rect 106730 255693 118102 255721
rect 106730 255681 106736 255693
rect 118096 255681 118102 255693
rect 118154 255681 118160 255733
rect 138160 255681 138166 255733
rect 138218 255721 138224 255733
rect 141136 255721 141142 255733
rect 138218 255693 141142 255721
rect 138218 255681 138224 255693
rect 141136 255681 141142 255693
rect 141194 255681 141200 255733
rect 151234 255721 151262 255841
rect 178576 255795 178582 255807
rect 166882 255767 178582 255795
rect 166882 255721 166910 255767
rect 178576 255755 178582 255767
rect 178634 255755 178640 255807
rect 178672 255755 178678 255807
rect 178730 255795 178736 255807
rect 178730 255767 191774 255795
rect 178730 255755 178736 255767
rect 151234 255693 166910 255721
rect 191746 255721 191774 255767
rect 218416 255755 218422 255807
rect 218474 255795 218480 255807
rect 218800 255795 218806 255807
rect 218474 255767 218806 255795
rect 218474 255755 218480 255767
rect 218800 255755 218806 255767
rect 218858 255755 218864 255807
rect 283714 255795 283742 255915
rect 284080 255903 284086 255955
rect 284138 255943 284144 255955
rect 300400 255943 300406 255955
rect 284138 255915 300406 255943
rect 284138 255903 284144 255915
rect 300400 255903 300406 255915
rect 300458 255903 300464 255955
rect 300496 255903 300502 255955
rect 300554 255943 300560 255955
rect 310576 255943 310582 255955
rect 300554 255915 310582 255943
rect 300554 255903 300560 255915
rect 310576 255903 310582 255915
rect 310634 255903 310640 255955
rect 310912 255903 310918 255955
rect 310970 255943 310976 255955
rect 363952 255943 363958 255955
rect 310970 255915 363958 255943
rect 310970 255903 310976 255915
rect 363952 255903 363958 255915
rect 364010 255903 364016 255955
rect 421552 255903 421558 255955
rect 421610 255943 421616 255955
rect 424432 255943 424438 255955
rect 421610 255915 424438 255943
rect 421610 255903 421616 255915
rect 424432 255903 424438 255915
rect 424490 255903 424496 255955
rect 288016 255829 288022 255881
rect 288074 255869 288080 255881
rect 288074 255841 300830 255869
rect 288074 255829 288080 255841
rect 300688 255795 300694 255807
rect 283714 255767 300694 255795
rect 300688 255755 300694 255767
rect 300746 255755 300752 255807
rect 300802 255795 300830 255841
rect 300880 255829 300886 255881
rect 300938 255869 300944 255881
rect 365392 255869 365398 255881
rect 300938 255841 365398 255869
rect 300938 255829 300944 255841
rect 365392 255829 365398 255841
rect 365450 255829 365456 255881
rect 423472 255829 423478 255881
rect 423530 255869 423536 255881
rect 423530 255841 433502 255869
rect 423530 255829 423536 255841
rect 423856 255795 423862 255807
rect 300802 255767 423862 255795
rect 423856 255755 423862 255767
rect 423914 255755 423920 255807
rect 218896 255721 218902 255733
rect 191746 255693 218902 255721
rect 218896 255681 218902 255693
rect 218954 255681 218960 255733
rect 259138 255693 259262 255721
rect 86704 255607 86710 255659
rect 86762 255647 86768 255659
rect 106480 255647 106486 255659
rect 86762 255619 106486 255647
rect 86762 255607 86768 255619
rect 106480 255607 106486 255619
rect 106538 255607 106544 255659
rect 259138 255647 259166 255693
rect 259234 255659 259262 255693
rect 293104 255681 293110 255733
rect 293162 255721 293168 255733
rect 300496 255721 300502 255733
rect 293162 255693 300502 255721
rect 293162 255681 293168 255693
rect 300496 255681 300502 255693
rect 300554 255681 300560 255733
rect 300784 255681 300790 255733
rect 300842 255721 300848 255733
rect 433474 255721 433502 255841
rect 541456 255755 541462 255807
rect 541514 255795 541520 255807
rect 541840 255795 541846 255807
rect 541514 255767 541846 255795
rect 541514 255755 541520 255767
rect 541840 255755 541846 255767
rect 541898 255755 541904 255807
rect 443536 255721 443542 255733
rect 300842 255693 383102 255721
rect 433474 255693 443542 255721
rect 300842 255681 300848 255693
rect 256258 255619 259166 255647
rect 256258 255573 256286 255619
rect 259216 255607 259222 255659
rect 259274 255607 259280 255659
rect 289456 255607 289462 255659
rect 289514 255647 289520 255659
rect 322288 255647 322294 255659
rect 289514 255619 322294 255647
rect 289514 255607 289520 255619
rect 322288 255607 322294 255619
rect 322346 255607 322352 255659
rect 322384 255607 322390 255659
rect 322442 255647 322448 255659
rect 324208 255647 324214 255659
rect 322442 255619 324214 255647
rect 322442 255607 322448 255619
rect 324208 255607 324214 255619
rect 324266 255607 324272 255659
rect 383074 255647 383102 255693
rect 443536 255681 443542 255693
rect 443594 255681 443600 255733
rect 443632 255681 443638 255733
rect 443690 255721 443696 255733
rect 443690 255693 463742 255721
rect 443690 255681 443696 255693
rect 423376 255647 423382 255659
rect 383074 255619 406334 255647
rect 60650 255545 80606 255573
rect 236194 255545 256286 255573
rect 60650 255533 60656 255545
rect 43600 255459 43606 255511
rect 43658 255499 43664 255511
rect 60496 255499 60502 255511
rect 43658 255471 60502 255499
rect 43658 255459 43664 255471
rect 60496 255459 60502 255471
rect 60554 255459 60560 255511
rect 218896 255459 218902 255511
rect 218954 255499 218960 255511
rect 236194 255499 236222 255545
rect 288592 255533 288598 255585
rect 288650 255573 288656 255585
rect 310768 255573 310774 255585
rect 288650 255545 310774 255573
rect 288650 255533 288656 255545
rect 310768 255533 310774 255545
rect 310826 255533 310832 255585
rect 310864 255533 310870 255585
rect 310922 255573 310928 255585
rect 337264 255573 337270 255585
rect 310922 255545 337270 255573
rect 310922 255533 310928 255545
rect 337264 255533 337270 255545
rect 337322 255533 337328 255585
rect 406306 255573 406334 255619
rect 408994 255619 423382 255647
rect 408994 255573 409022 255619
rect 423376 255607 423382 255619
rect 423434 255607 423440 255659
rect 463714 255647 463742 255693
rect 490960 255681 490966 255733
rect 491018 255721 491024 255733
rect 501136 255721 501142 255733
rect 491018 255693 501142 255721
rect 491018 255681 491024 255693
rect 501136 255681 501142 255693
rect 501194 255681 501200 255733
rect 570160 255721 570166 255733
rect 541474 255693 570166 255721
rect 469360 255647 469366 255659
rect 463714 255619 469366 255647
rect 469360 255607 469366 255619
rect 469418 255607 469424 255659
rect 538480 255607 538486 255659
rect 538538 255647 538544 255659
rect 541474 255647 541502 255693
rect 570160 255681 570166 255693
rect 570218 255681 570224 255733
rect 590512 255681 590518 255733
rect 590570 255721 590576 255733
rect 601936 255721 601942 255733
rect 590570 255693 601942 255721
rect 590570 255681 590576 255693
rect 601936 255681 601942 255693
rect 601994 255681 602000 255733
rect 622000 255681 622006 255733
rect 622058 255721 622064 255733
rect 630640 255721 630646 255733
rect 622058 255693 630646 255721
rect 622058 255681 622064 255693
rect 630640 255681 630646 255693
rect 630698 255681 630704 255733
rect 671056 255721 671062 255733
rect 665218 255693 671062 255721
rect 538538 255619 541502 255647
rect 538538 255607 538544 255619
rect 570352 255607 570358 255659
rect 570410 255647 570416 255659
rect 590320 255647 590326 255659
rect 570410 255619 590326 255647
rect 570410 255607 570416 255619
rect 590320 255607 590326 255619
rect 590378 255607 590384 255659
rect 630832 255607 630838 255659
rect 630890 255647 630896 255659
rect 642256 255647 642262 255659
rect 630890 255619 642262 255647
rect 630890 255607 630896 255619
rect 642256 255607 642262 255619
rect 642314 255607 642320 255659
rect 662320 255607 662326 255659
rect 662378 255647 662384 255659
rect 665218 255647 665246 255693
rect 671056 255681 671062 255693
rect 671114 255681 671120 255733
rect 662378 255619 665246 255647
rect 662378 255607 662384 255619
rect 490960 255573 490966 255585
rect 406306 255545 409022 255573
rect 480994 255545 490966 255573
rect 218954 255471 236222 255499
rect 218954 255459 218960 255471
rect 286288 255459 286294 255511
rect 286346 255499 286352 255511
rect 363568 255499 363574 255511
rect 286346 255471 363574 255499
rect 286346 255459 286352 255471
rect 363568 255459 363574 255471
rect 363626 255459 363632 255511
rect 469360 255459 469366 255511
rect 469418 255499 469424 255511
rect 480994 255499 481022 255545
rect 490960 255533 490966 255545
rect 491018 255533 491024 255585
rect 469418 255471 481022 255499
rect 469418 255459 469424 255471
rect 301072 255385 301078 255437
rect 301130 255425 301136 255437
rect 364240 255425 364246 255437
rect 301130 255397 364246 255425
rect 301130 255385 301136 255397
rect 364240 255385 364246 255397
rect 364298 255385 364304 255437
rect 283216 255311 283222 255363
rect 283274 255351 283280 255363
rect 364624 255351 364630 255363
rect 283274 255323 364630 255351
rect 283274 255311 283280 255323
rect 364624 255311 364630 255323
rect 364682 255311 364688 255363
rect 284176 255237 284182 255289
rect 284234 255277 284240 255289
rect 365008 255277 365014 255289
rect 284234 255249 365014 255277
rect 284234 255237 284240 255249
rect 365008 255237 365014 255249
rect 365066 255237 365072 255289
rect 518416 255237 518422 255289
rect 518474 255277 518480 255289
rect 519856 255277 519862 255289
rect 518474 255249 519862 255277
rect 518474 255237 518480 255249
rect 519856 255237 519862 255249
rect 519914 255237 519920 255289
rect 286960 255163 286966 255215
rect 287018 255203 287024 255215
rect 367984 255203 367990 255215
rect 287018 255175 367990 255203
rect 287018 255163 287024 255175
rect 367984 255163 367990 255175
rect 368042 255163 368048 255215
rect 287824 255089 287830 255141
rect 287882 255129 287888 255141
rect 366448 255129 366454 255141
rect 287882 255101 366454 255129
rect 287882 255089 287888 255101
rect 366448 255089 366454 255101
rect 366506 255089 366512 255141
rect 283408 255015 283414 255067
rect 283466 255055 283472 255067
rect 368656 255055 368662 255067
rect 283466 255027 300926 255055
rect 283466 255015 283472 255027
rect 83536 254941 83542 254993
rect 83594 254981 83600 254993
rect 112144 254981 112150 254993
rect 83594 254953 112150 254981
rect 83594 254941 83600 254953
rect 112144 254941 112150 254953
rect 112202 254941 112208 254993
rect 277072 254941 277078 254993
rect 277130 254981 277136 254993
rect 293584 254981 293590 254993
rect 277130 254953 293590 254981
rect 277130 254941 277136 254953
rect 293584 254941 293590 254953
rect 293642 254941 293648 254993
rect 300898 254981 300926 255027
rect 310978 255027 368662 255055
rect 310978 254981 311006 255027
rect 368656 255015 368662 255027
rect 368714 255015 368720 255067
rect 388720 255015 388726 255067
rect 388778 255055 388784 255067
rect 391504 255055 391510 255067
rect 388778 255027 391510 255055
rect 388778 255015 388784 255027
rect 391504 255015 391510 255027
rect 391562 255015 391568 255067
rect 300898 254953 311006 254981
rect 319792 254941 319798 254993
rect 319850 254981 319856 254993
rect 440752 254981 440758 254993
rect 319850 254953 440758 254981
rect 319850 254941 319856 254953
rect 440752 254941 440758 254953
rect 440810 254941 440816 254993
rect 65200 254867 65206 254919
rect 65258 254907 65264 254919
rect 200272 254907 200278 254919
rect 65258 254879 200278 254907
rect 65258 254867 65264 254879
rect 200272 254867 200278 254879
rect 200330 254867 200336 254919
rect 288112 254867 288118 254919
rect 288170 254907 288176 254919
rect 319888 254907 319894 254919
rect 288170 254879 319894 254907
rect 288170 254867 288176 254879
rect 319888 254867 319894 254879
rect 319946 254867 319952 254919
rect 321616 254867 321622 254919
rect 321674 254907 321680 254919
rect 443632 254907 443638 254919
rect 321674 254879 443638 254907
rect 321674 254867 321680 254879
rect 443632 254867 443638 254879
rect 443690 254867 443696 254919
rect 295312 254793 295318 254845
rect 295370 254833 295376 254845
rect 320848 254833 320854 254845
rect 295370 254805 320854 254833
rect 295370 254793 295376 254805
rect 320848 254793 320854 254805
rect 320906 254793 320912 254845
rect 322384 254793 322390 254845
rect 322442 254833 322448 254845
rect 443536 254833 443542 254845
rect 322442 254805 443542 254833
rect 322442 254793 322448 254805
rect 443536 254793 443542 254805
rect 443594 254793 443600 254845
rect 316816 254719 316822 254771
rect 316874 254759 316880 254771
rect 440656 254759 440662 254771
rect 316874 254731 440662 254759
rect 316874 254719 316880 254731
rect 440656 254719 440662 254731
rect 440714 254719 440720 254771
rect 285424 254645 285430 254697
rect 285482 254685 285488 254697
rect 414352 254685 414358 254697
rect 285482 254657 414358 254685
rect 285482 254645 285488 254657
rect 414352 254645 414358 254657
rect 414410 254645 414416 254697
rect 285520 254571 285526 254623
rect 285578 254611 285584 254623
rect 412144 254611 412150 254623
rect 285578 254583 412150 254611
rect 285578 254571 285584 254583
rect 412144 254571 412150 254583
rect 412202 254571 412208 254623
rect 282928 254497 282934 254549
rect 282986 254537 282992 254549
rect 413968 254537 413974 254549
rect 282986 254509 413974 254537
rect 282986 254497 282992 254509
rect 413968 254497 413974 254509
rect 414026 254497 414032 254549
rect 283984 254423 283990 254475
rect 284042 254463 284048 254475
rect 301072 254463 301078 254475
rect 284042 254435 301078 254463
rect 284042 254423 284048 254435
rect 301072 254423 301078 254435
rect 301130 254423 301136 254475
rect 310096 254423 310102 254475
rect 310154 254463 310160 254475
rect 310960 254463 310966 254475
rect 310154 254435 310966 254463
rect 310154 254423 310160 254435
rect 310960 254423 310966 254435
rect 311018 254423 311024 254475
rect 316048 254423 316054 254475
rect 316106 254463 316112 254475
rect 446416 254463 446422 254475
rect 316106 254435 446422 254463
rect 316106 254423 316112 254435
rect 446416 254423 446422 254435
rect 446474 254423 446480 254475
rect 318256 254349 318262 254401
rect 318314 254389 318320 254401
rect 445360 254389 445366 254401
rect 318314 254361 445366 254389
rect 318314 254349 318320 254361
rect 445360 254349 445366 254361
rect 445418 254349 445424 254401
rect 317584 254275 317590 254327
rect 317642 254315 317648 254327
rect 444304 254315 444310 254327
rect 317642 254287 444310 254315
rect 317642 254275 317648 254287
rect 444304 254275 444310 254287
rect 444362 254275 444368 254327
rect 284272 254201 284278 254253
rect 284330 254241 284336 254253
rect 298288 254241 298294 254253
rect 284330 254213 298294 254241
rect 284330 254201 284336 254213
rect 298288 254201 298294 254213
rect 298346 254201 298352 254253
rect 315376 254201 315382 254253
rect 315434 254241 315440 254253
rect 446416 254241 446422 254253
rect 315434 254213 446422 254241
rect 315434 254201 315440 254213
rect 446416 254201 446422 254213
rect 446474 254201 446480 254253
rect 287248 254127 287254 254179
rect 287306 254167 287312 254179
rect 421360 254167 421366 254179
rect 287306 254139 421366 254167
rect 287306 254127 287312 254139
rect 421360 254127 421366 254139
rect 421418 254127 421424 254179
rect 287344 254053 287350 254105
rect 287402 254093 287408 254105
rect 422032 254093 422038 254105
rect 287402 254065 422038 254093
rect 287402 254053 287408 254065
rect 422032 254053 422038 254065
rect 422090 254053 422096 254105
rect 284848 253979 284854 254031
rect 284906 254019 284912 254031
rect 420208 254019 420214 254031
rect 284906 253991 420214 254019
rect 284906 253979 284912 253991
rect 420208 253979 420214 253991
rect 420266 253979 420272 254031
rect 287152 253905 287158 253957
rect 287210 253945 287216 253957
rect 423184 253945 423190 253957
rect 287210 253917 423190 253945
rect 287210 253905 287216 253917
rect 423184 253905 423190 253917
rect 423242 253905 423248 253957
rect 285712 253831 285718 253883
rect 285770 253871 285776 253883
rect 290992 253871 290998 253883
rect 285770 253843 290998 253871
rect 285770 253831 285776 253843
rect 290992 253831 290998 253843
rect 291050 253831 291056 253883
rect 298288 253831 298294 253883
rect 298346 253871 298352 253883
rect 420592 253871 420598 253883
rect 298346 253843 420598 253871
rect 298346 253831 298352 253843
rect 420592 253831 420598 253843
rect 420650 253831 420656 253883
rect 288304 253757 288310 253809
rect 288362 253797 288368 253809
rect 322480 253797 322486 253809
rect 288362 253769 322486 253797
rect 288362 253757 288368 253769
rect 322480 253757 322486 253769
rect 322538 253757 322544 253809
rect 322576 253757 322582 253809
rect 322634 253797 322640 253809
rect 338320 253797 338326 253809
rect 322634 253769 338326 253797
rect 322634 253757 322640 253769
rect 338320 253757 338326 253769
rect 338378 253757 338384 253809
rect 351376 253757 351382 253809
rect 351434 253797 351440 253809
rect 360784 253797 360790 253809
rect 351434 253769 360790 253797
rect 351434 253757 351440 253769
rect 360784 253757 360790 253769
rect 360842 253757 360848 253809
rect 285040 253683 285046 253735
rect 285098 253723 285104 253735
rect 422800 253723 422806 253735
rect 285098 253695 422806 253723
rect 285098 253683 285104 253695
rect 422800 253683 422806 253695
rect 422858 253683 422864 253735
rect 284944 253609 284950 253661
rect 285002 253649 285008 253661
rect 290896 253649 290902 253661
rect 285002 253621 290902 253649
rect 285002 253609 285008 253621
rect 290896 253609 290902 253621
rect 290954 253609 290960 253661
rect 290992 253609 290998 253661
rect 291050 253649 291056 253661
rect 362416 253649 362422 253661
rect 291050 253621 362422 253649
rect 291050 253609 291056 253621
rect 362416 253609 362422 253621
rect 362474 253609 362480 253661
rect 204400 253535 204406 253587
rect 204458 253575 204464 253587
rect 316720 253575 316726 253587
rect 204458 253547 316726 253575
rect 204458 253535 204464 253547
rect 316720 253535 316726 253547
rect 316778 253535 316784 253587
rect 322480 253535 322486 253587
rect 322538 253575 322544 253587
rect 323056 253575 323062 253587
rect 322538 253547 323062 253575
rect 322538 253535 322544 253547
rect 323056 253535 323062 253547
rect 323114 253535 323120 253587
rect 338320 253535 338326 253587
rect 338378 253575 338384 253587
rect 495280 253575 495286 253587
rect 338378 253547 495286 253575
rect 338378 253535 338384 253547
rect 495280 253535 495286 253547
rect 495338 253535 495344 253587
rect 287632 253461 287638 253513
rect 287690 253501 287696 253513
rect 367216 253501 367222 253513
rect 287690 253473 367222 253501
rect 287690 253461 287696 253473
rect 367216 253461 367222 253473
rect 367274 253461 367280 253513
rect 288496 253387 288502 253439
rect 288554 253427 288560 253439
rect 508336 253427 508342 253439
rect 288554 253399 508342 253427
rect 288554 253387 288560 253399
rect 508336 253387 508342 253399
rect 508394 253387 508400 253439
rect 674800 253387 674806 253439
rect 674858 253427 674864 253439
rect 676816 253427 676822 253439
rect 674858 253399 676822 253427
rect 674858 253387 674864 253399
rect 676816 253387 676822 253399
rect 676874 253387 676880 253439
rect 287920 253313 287926 253365
rect 287978 253353 287984 253365
rect 370576 253353 370582 253365
rect 287978 253325 370582 253353
rect 287978 253313 287984 253325
rect 370576 253313 370582 253325
rect 370634 253313 370640 253365
rect 283024 253239 283030 253291
rect 283082 253279 283088 253291
rect 300880 253279 300886 253291
rect 283082 253251 300886 253279
rect 283082 253239 283088 253251
rect 300880 253239 300886 253251
rect 300938 253239 300944 253291
rect 282832 253165 282838 253217
rect 282890 253205 282896 253217
rect 371248 253205 371254 253217
rect 282890 253177 371254 253205
rect 282890 253165 282896 253177
rect 371248 253165 371254 253177
rect 371306 253165 371312 253217
rect 418000 253165 418006 253217
rect 418058 253205 418064 253217
rect 440272 253205 440278 253217
rect 418058 253177 440278 253205
rect 418058 253165 418064 253177
rect 440272 253165 440278 253177
rect 440330 253165 440336 253217
rect 140176 253091 140182 253143
rect 140234 253131 140240 253143
rect 141520 253131 141526 253143
rect 140234 253103 141526 253131
rect 140234 253091 140240 253103
rect 141520 253091 141526 253103
rect 141578 253091 141584 253143
rect 287440 253091 287446 253143
rect 287498 253131 287504 253143
rect 372400 253131 372406 253143
rect 287498 253103 372406 253131
rect 287498 253091 287504 253103
rect 372400 253091 372406 253103
rect 372458 253091 372464 253143
rect 416944 253091 416950 253143
rect 417002 253131 417008 253143
rect 446416 253131 446422 253143
rect 417002 253103 446422 253131
rect 417002 253091 417008 253103
rect 446416 253091 446422 253103
rect 446474 253091 446480 253143
rect 287728 253017 287734 253069
rect 287786 253057 287792 253069
rect 371632 253057 371638 253069
rect 287786 253029 371638 253057
rect 287786 253017 287792 253029
rect 371632 253017 371638 253029
rect 371690 253017 371696 253069
rect 423568 253017 423574 253069
rect 423626 253057 423632 253069
rect 423626 253029 435422 253057
rect 423626 253017 423632 253029
rect 112144 252943 112150 252995
rect 112202 252983 112208 252995
rect 142480 252983 142486 252995
rect 112202 252955 142486 252983
rect 112202 252943 112208 252955
rect 142480 252943 142486 252955
rect 142538 252943 142544 252995
rect 287536 252943 287542 252995
rect 287594 252983 287600 252995
rect 372736 252983 372742 252995
rect 287594 252955 372742 252983
rect 287594 252943 287600 252955
rect 372736 252943 372742 252955
rect 372794 252943 372800 252995
rect 388432 252943 388438 252995
rect 388490 252983 388496 252995
rect 392992 252983 392998 252995
rect 388490 252955 392998 252983
rect 388490 252943 388496 252955
rect 392992 252943 392998 252955
rect 393050 252943 393056 252995
rect 435394 252983 435422 253029
rect 445360 252983 445366 252995
rect 435394 252955 445366 252983
rect 445360 252943 445366 252955
rect 445418 252943 445424 252995
rect 96304 252869 96310 252921
rect 96362 252909 96368 252921
rect 141136 252909 141142 252921
rect 96362 252881 141142 252909
rect 96362 252869 96368 252881
rect 141136 252869 141142 252881
rect 141194 252869 141200 252921
rect 287824 252869 287830 252921
rect 287882 252909 287888 252921
rect 372016 252909 372022 252921
rect 287882 252881 372022 252909
rect 287882 252869 287888 252881
rect 372016 252869 372022 252881
rect 372074 252869 372080 252921
rect 416560 252869 416566 252921
rect 416618 252909 416624 252921
rect 444976 252909 444982 252921
rect 416618 252881 444982 252909
rect 416618 252869 416624 252881
rect 444976 252869 444982 252881
rect 445034 252869 445040 252921
rect 446224 252869 446230 252921
rect 446282 252869 446288 252921
rect 80848 252795 80854 252847
rect 80906 252835 80912 252847
rect 146800 252835 146806 252847
rect 80906 252807 146806 252835
rect 80906 252795 80912 252807
rect 146800 252795 146806 252807
rect 146858 252795 146864 252847
rect 284368 252795 284374 252847
rect 284426 252835 284432 252847
rect 411376 252835 411382 252847
rect 284426 252807 411382 252835
rect 284426 252795 284432 252807
rect 411376 252795 411382 252807
rect 411434 252795 411440 252847
rect 417280 252795 417286 252847
rect 417338 252835 417344 252847
rect 446242 252835 446270 252869
rect 417338 252807 446270 252835
rect 417338 252795 417344 252807
rect 67600 252721 67606 252773
rect 67658 252761 67664 252773
rect 146896 252761 146902 252773
rect 67658 252733 146902 252761
rect 67658 252721 67664 252733
rect 146896 252721 146902 252733
rect 146954 252721 146960 252773
rect 45328 252647 45334 252699
rect 45386 252687 45392 252699
rect 200368 252687 200374 252699
rect 45386 252659 200374 252687
rect 45386 252647 45392 252659
rect 200368 252647 200374 252659
rect 200426 252647 200432 252699
rect 45040 252573 45046 252625
rect 45098 252613 45104 252625
rect 200176 252613 200182 252625
rect 45098 252585 200182 252613
rect 45098 252573 45104 252585
rect 200176 252573 200182 252585
rect 200234 252573 200240 252625
rect 45424 252499 45430 252551
rect 45482 252539 45488 252551
rect 200560 252539 200566 252551
rect 45482 252511 200566 252539
rect 45482 252499 45488 252511
rect 200560 252499 200566 252511
rect 200618 252499 200624 252551
rect 44848 252425 44854 252477
rect 44906 252465 44912 252477
rect 200464 252465 200470 252477
rect 44906 252437 200470 252465
rect 44906 252425 44912 252437
rect 200464 252425 200470 252437
rect 200522 252425 200528 252477
rect 45232 252351 45238 252403
rect 45290 252391 45296 252403
rect 204496 252391 204502 252403
rect 45290 252363 204502 252391
rect 45290 252351 45296 252363
rect 204496 252351 204502 252363
rect 204554 252351 204560 252403
rect 45136 252277 45142 252329
rect 45194 252317 45200 252329
rect 204688 252317 204694 252329
rect 45194 252289 204694 252317
rect 45194 252277 45200 252289
rect 204688 252277 204694 252289
rect 204746 252277 204752 252329
rect 44944 252203 44950 252255
rect 45002 252243 45008 252255
rect 204880 252243 204886 252255
rect 45002 252215 204886 252243
rect 45002 252203 45008 252215
rect 204880 252203 204886 252215
rect 204938 252203 204944 252255
rect 44752 252129 44758 252181
rect 44810 252169 44816 252181
rect 204784 252169 204790 252181
rect 44810 252141 204790 252169
rect 44810 252129 44816 252141
rect 204784 252129 204790 252141
rect 204842 252129 204848 252181
rect 44560 252055 44566 252107
rect 44618 252095 44624 252107
rect 204592 252095 204598 252107
rect 44618 252067 204598 252095
rect 44618 252055 44624 252067
rect 204592 252055 204598 252067
rect 204650 252055 204656 252107
rect 44656 251981 44662 252033
rect 44714 252021 44720 252033
rect 204208 252021 204214 252033
rect 44714 251993 204214 252021
rect 44714 251981 44720 251993
rect 204208 251981 204214 251993
rect 204266 251981 204272 252033
rect 675376 251167 675382 251219
rect 675434 251167 675440 251219
rect 283312 251093 283318 251145
rect 283370 251133 283376 251145
rect 283696 251133 283702 251145
rect 283370 251105 283702 251133
rect 283370 251093 283376 251105
rect 283696 251093 283702 251105
rect 283754 251093 283760 251145
rect 675394 250997 675422 251167
rect 283120 250945 283126 250997
rect 283178 250985 283184 250997
rect 283312 250985 283318 250997
rect 283178 250957 283318 250985
rect 283178 250945 283184 250957
rect 283312 250945 283318 250957
rect 283370 250945 283376 250997
rect 675376 250945 675382 250997
rect 675434 250945 675440 250997
rect 282736 250797 282742 250849
rect 282794 250837 282800 250849
rect 283120 250837 283126 250849
rect 282794 250809 283126 250837
rect 282794 250797 282800 250809
rect 283120 250797 283126 250809
rect 283178 250797 283184 250849
rect 139216 250723 139222 250775
rect 139274 250763 139280 250775
rect 140176 250763 140182 250775
rect 139274 250735 140182 250763
rect 139274 250723 139280 250735
rect 140176 250723 140182 250735
rect 140234 250723 140240 250775
rect 42160 250575 42166 250627
rect 42218 250615 42224 250627
rect 42218 250587 139166 250615
rect 42218 250575 42224 250587
rect 139138 250541 139166 250587
rect 145360 250575 145366 250627
rect 145418 250615 145424 250627
rect 182320 250615 182326 250627
rect 145418 250587 182326 250615
rect 145418 250575 145424 250587
rect 182320 250575 182326 250587
rect 182378 250575 182384 250627
rect 139138 250513 139262 250541
rect 139234 250319 139262 250513
rect 230128 250501 230134 250553
rect 230186 250541 230192 250553
rect 282736 250541 282742 250553
rect 230186 250513 282742 250541
rect 230186 250501 230192 250513
rect 282736 250501 282742 250513
rect 282794 250501 282800 250553
rect 145360 250393 145366 250405
rect 139810 250365 145366 250393
rect 139810 250319 139838 250365
rect 145360 250353 145366 250365
rect 145418 250353 145424 250405
rect 139234 250291 139838 250319
rect 141136 250279 141142 250331
rect 141194 250319 141200 250331
rect 144400 250319 144406 250331
rect 141194 250291 144406 250319
rect 141194 250279 141200 250291
rect 144400 250279 144406 250291
rect 144458 250279 144464 250331
rect 139312 250205 139318 250257
rect 139370 250245 139376 250257
rect 144304 250245 144310 250257
rect 139370 250217 144310 250245
rect 139370 250205 139376 250217
rect 144304 250205 144310 250217
rect 144362 250205 144368 250257
rect 674800 250205 674806 250257
rect 674858 250245 674864 250257
rect 675280 250245 675286 250257
rect 674858 250217 675286 250245
rect 674858 250205 674864 250217
rect 675280 250205 675286 250217
rect 675338 250205 675344 250257
rect 139792 250131 139798 250183
rect 139850 250171 139856 250183
rect 141328 250171 141334 250183
rect 139850 250143 141334 250171
rect 139850 250131 139856 250143
rect 141328 250131 141334 250143
rect 141386 250131 141392 250183
rect 139888 250057 139894 250109
rect 139946 250097 139952 250109
rect 141232 250097 141238 250109
rect 139946 250069 141238 250097
rect 139946 250057 139952 250069
rect 141232 250057 141238 250069
rect 141290 250057 141296 250109
rect 44560 249983 44566 250035
rect 44618 250023 44624 250035
rect 200080 250023 200086 250035
rect 44618 249995 200086 250023
rect 44618 249983 44624 249995
rect 200080 249983 200086 249995
rect 200138 249983 200144 250035
rect 218416 249095 218422 249147
rect 218474 249135 218480 249147
rect 218800 249135 218806 249147
rect 218474 249107 218806 249135
rect 218474 249095 218480 249107
rect 218800 249095 218806 249107
rect 218858 249095 218864 249147
rect 541456 249095 541462 249147
rect 541514 249135 541520 249147
rect 541840 249135 541846 249147
rect 541514 249107 541846 249135
rect 541514 249095 541520 249107
rect 541840 249095 541846 249107
rect 541898 249095 541904 249147
rect 282352 248873 282358 248925
rect 282410 248913 282416 248925
rect 283888 248913 283894 248925
rect 282410 248885 283894 248913
rect 282410 248873 282416 248885
rect 283888 248873 283894 248885
rect 283946 248873 283952 248925
rect 288304 248355 288310 248407
rect 288362 248355 288368 248407
rect 288112 248281 288118 248333
rect 288170 248281 288176 248333
rect 288016 248133 288022 248185
rect 288074 248173 288080 248185
rect 288130 248173 288158 248281
rect 288074 248145 288158 248173
rect 288074 248133 288080 248145
rect 144016 247763 144022 247815
rect 144074 247803 144080 247815
rect 191440 247803 191446 247815
rect 144074 247775 191446 247803
rect 144074 247763 144080 247775
rect 191440 247763 191446 247775
rect 191498 247763 191504 247815
rect 285616 247763 285622 247815
rect 285674 247803 285680 247815
rect 285674 247775 286046 247803
rect 285674 247763 285680 247775
rect 286018 247741 286046 247775
rect 145456 247689 145462 247741
rect 145514 247729 145520 247741
rect 148240 247729 148246 247741
rect 145514 247701 148246 247729
rect 145514 247689 145520 247701
rect 148240 247689 148246 247701
rect 148298 247689 148304 247741
rect 286000 247689 286006 247741
rect 286058 247689 286064 247741
rect 288322 247667 288350 248355
rect 532912 247689 532918 247741
rect 532970 247729 532976 247741
rect 533392 247729 533398 247741
rect 532970 247701 533398 247729
rect 532970 247689 532976 247701
rect 533392 247689 533398 247701
rect 533450 247689 533456 247741
rect 541552 247689 541558 247741
rect 541610 247729 541616 247741
rect 541744 247729 541750 247741
rect 541610 247701 541750 247729
rect 541610 247689 541616 247701
rect 541744 247689 541750 247701
rect 541802 247689 541808 247741
rect 34576 247615 34582 247667
rect 34634 247655 34640 247667
rect 42160 247655 42166 247667
rect 34634 247627 42166 247655
rect 34634 247615 34640 247627
rect 42160 247615 42166 247627
rect 42218 247615 42224 247667
rect 235888 247615 235894 247667
rect 235946 247655 235952 247667
rect 282352 247655 282358 247667
rect 235946 247627 282358 247655
rect 235946 247615 235952 247627
rect 282352 247615 282358 247627
rect 282410 247615 282416 247667
rect 285616 247615 285622 247667
rect 285674 247655 285680 247667
rect 285904 247655 285910 247667
rect 285674 247627 285910 247655
rect 285674 247615 285680 247627
rect 285904 247615 285910 247627
rect 285962 247615 285968 247667
rect 288304 247615 288310 247667
rect 288362 247615 288368 247667
rect 182320 247541 182326 247593
rect 182378 247581 182384 247593
rect 200752 247581 200758 247593
rect 182378 247553 200758 247581
rect 182378 247541 182384 247553
rect 200752 247541 200758 247553
rect 200810 247541 200816 247593
rect 674416 246727 674422 246779
rect 674474 246767 674480 246779
rect 675184 246767 675190 246779
rect 674474 246739 675190 246767
rect 674474 246727 674480 246739
rect 675184 246727 675190 246739
rect 675242 246727 675248 246779
rect 282736 245247 282742 245299
rect 282794 245287 282800 245299
rect 282794 245259 284414 245287
rect 282794 245247 282800 245259
rect 282736 245099 282742 245151
rect 282794 245139 282800 245151
rect 283312 245139 283318 245151
rect 282794 245111 283318 245139
rect 282794 245099 282800 245111
rect 283312 245099 283318 245111
rect 283370 245099 283376 245151
rect 144112 244877 144118 244929
rect 144170 244917 144176 244929
rect 148432 244917 148438 244929
rect 144170 244889 148438 244917
rect 144170 244877 144176 244889
rect 148432 244877 148438 244889
rect 148490 244877 148496 244929
rect 144016 244803 144022 244855
rect 144074 244843 144080 244855
rect 197200 244843 197206 244855
rect 144074 244815 197206 244843
rect 144074 244803 144080 244815
rect 197200 244803 197206 244815
rect 197258 244803 197264 244855
rect 282160 244803 282166 244855
rect 282218 244843 282224 244855
rect 282640 244843 282646 244855
rect 282218 244815 282646 244843
rect 282218 244803 282224 244815
rect 282640 244803 282646 244815
rect 282698 244803 282704 244855
rect 283792 244803 283798 244855
rect 283850 244843 283856 244855
rect 284272 244843 284278 244855
rect 283850 244815 284278 244843
rect 283850 244803 283856 244815
rect 284272 244803 284278 244815
rect 284330 244803 284336 244855
rect 42064 244729 42070 244781
rect 42122 244769 42128 244781
rect 42544 244769 42550 244781
rect 42122 244741 42550 244769
rect 42122 244729 42128 244741
rect 42544 244729 42550 244741
rect 42602 244729 42608 244781
rect 241648 244729 241654 244781
rect 241706 244769 241712 244781
rect 282256 244769 282262 244781
rect 241706 244741 282262 244769
rect 241706 244729 241712 244741
rect 282256 244729 282262 244741
rect 282314 244729 282320 244781
rect 253360 244655 253366 244707
rect 253418 244695 253424 244707
rect 284272 244695 284278 244707
rect 253418 244667 284278 244695
rect 253418 244655 253424 244667
rect 284272 244655 284278 244667
rect 284330 244655 284336 244707
rect 262000 244581 262006 244633
rect 262058 244621 262064 244633
rect 282256 244621 282262 244633
rect 262058 244593 282262 244621
rect 262058 244581 262064 244593
rect 282256 244581 282262 244593
rect 282314 244581 282320 244633
rect 282448 244581 282454 244633
rect 282506 244621 282512 244633
rect 282640 244621 282646 244633
rect 282506 244593 282646 244621
rect 282506 244581 282512 244593
rect 282640 244581 282646 244593
rect 282698 244581 282704 244633
rect 284386 244621 284414 245259
rect 288304 244729 288310 244781
rect 288362 244729 288368 244781
rect 284290 244593 284414 244621
rect 267760 244507 267766 244559
rect 267818 244547 267824 244559
rect 283024 244547 283030 244559
rect 267818 244519 283030 244547
rect 267818 244507 267824 244519
rect 283024 244507 283030 244519
rect 283082 244507 283088 244559
rect 37264 244433 37270 244485
rect 37322 244473 37328 244485
rect 41776 244473 41782 244485
rect 37322 244445 41782 244473
rect 37322 244433 37328 244445
rect 41776 244433 41782 244445
rect 41834 244433 41840 244485
rect 144400 244433 144406 244485
rect 144458 244473 144464 244485
rect 149584 244473 149590 244485
rect 144458 244445 149590 244473
rect 144458 244433 144464 244445
rect 149584 244433 149590 244445
rect 149642 244433 149648 244485
rect 276400 244433 276406 244485
rect 276458 244473 276464 244485
rect 282448 244473 282454 244485
rect 276458 244445 282454 244473
rect 276458 244433 276464 244445
rect 282448 244433 282454 244445
rect 282506 244433 282512 244485
rect 284290 244041 284318 244593
rect 288322 244559 288350 244729
rect 288304 244507 288310 244559
rect 288362 244507 288368 244559
rect 284272 243989 284278 244041
rect 284330 243989 284336 244041
rect 139984 243619 139990 243671
rect 140042 243659 140048 243671
rect 142192 243659 142198 243671
rect 140042 243631 142198 243659
rect 140042 243619 140048 243631
rect 142192 243619 142198 243631
rect 142250 243619 142256 243671
rect 674992 242953 674998 243005
rect 675050 242993 675056 243005
rect 675376 242993 675382 243005
rect 675050 242965 675382 242993
rect 675050 242953 675056 242965
rect 675376 242953 675382 242965
rect 675434 242953 675440 243005
rect 674128 242361 674134 242413
rect 674186 242401 674192 242413
rect 675376 242401 675382 242413
rect 674186 242373 675382 242401
rect 674186 242361 674192 242373
rect 675376 242361 675382 242373
rect 675434 242361 675440 242413
rect 41968 242287 41974 242339
rect 42026 242327 42032 242339
rect 42736 242327 42742 242339
rect 42026 242299 42742 242327
rect 42026 242287 42032 242299
rect 42736 242287 42742 242299
rect 42794 242287 42800 242339
rect 43120 242065 43126 242117
rect 43178 242105 43184 242117
rect 43504 242105 43510 242117
rect 43178 242077 43510 242105
rect 43178 242065 43184 242077
rect 43504 242065 43510 242077
rect 43562 242065 43568 242117
rect 37168 241991 37174 242043
rect 37226 242031 37232 242043
rect 42640 242031 42646 242043
rect 37226 242003 42646 242031
rect 37226 241991 37232 242003
rect 42640 241991 42646 242003
rect 42698 241991 42704 242043
rect 144016 241991 144022 242043
rect 144074 242031 144080 242043
rect 151120 242031 151126 242043
rect 144074 242003 151126 242031
rect 144074 241991 144080 242003
rect 151120 241991 151126 242003
rect 151178 241991 151184 242043
rect 288304 241991 288310 242043
rect 288362 241991 288368 242043
rect 37360 241917 37366 241969
rect 37418 241957 37424 241969
rect 43120 241957 43126 241969
rect 37418 241929 43126 241957
rect 37418 241917 37424 241929
rect 43120 241917 43126 241929
rect 43178 241917 43184 241969
rect 145744 241917 145750 241969
rect 145802 241957 145808 241969
rect 148624 241957 148630 241969
rect 145802 241929 148630 241957
rect 145802 241917 145808 241929
rect 148624 241917 148630 241929
rect 148682 241917 148688 241969
rect 204208 241917 204214 241969
rect 204266 241957 204272 241969
rect 207376 241957 207382 241969
rect 204266 241929 207382 241957
rect 204266 241917 204272 241929
rect 207376 241917 207382 241929
rect 207434 241917 207440 241969
rect 146800 241843 146806 241895
rect 146858 241883 146864 241895
rect 152080 241883 152086 241895
rect 146858 241855 152086 241883
rect 146858 241843 146864 241855
rect 152080 241843 152086 241855
rect 152138 241843 152144 241895
rect 288322 241821 288350 241991
rect 288304 241769 288310 241821
rect 288362 241769 288368 241821
rect 674320 241695 674326 241747
rect 674378 241735 674384 241747
rect 675472 241735 675478 241747
rect 674378 241707 675478 241735
rect 674378 241695 674384 241707
rect 675472 241695 675478 241707
rect 675530 241695 675536 241747
rect 42736 240733 42742 240785
rect 42794 240773 42800 240785
rect 43216 240773 43222 240785
rect 42794 240745 43222 240773
rect 42794 240733 42800 240745
rect 43216 240733 43222 240745
rect 43274 240733 43280 240785
rect 41776 240585 41782 240637
rect 41834 240585 41840 240637
rect 41794 240415 41822 240585
rect 674896 240511 674902 240563
rect 674954 240551 674960 240563
rect 675472 240551 675478 240563
rect 674954 240523 675478 240551
rect 674954 240511 674960 240523
rect 675472 240511 675478 240523
rect 675530 240511 675536 240563
rect 140176 240437 140182 240489
rect 140234 240477 140240 240489
rect 141424 240477 141430 240489
rect 140234 240449 141430 240477
rect 140234 240437 140240 240449
rect 141424 240437 141430 240449
rect 141482 240437 141488 240489
rect 41776 240363 41782 240415
rect 41834 240363 41840 240415
rect 288592 239623 288598 239675
rect 288650 239663 288656 239675
rect 290512 239663 290518 239675
rect 288650 239635 290518 239663
rect 288650 239623 288656 239635
rect 290512 239623 290518 239635
rect 290570 239623 290576 239675
rect 366688 239623 366694 239675
rect 366746 239663 366752 239675
rect 373936 239663 373942 239675
rect 366746 239635 373942 239663
rect 366746 239623 366752 239635
rect 373936 239623 373942 239635
rect 373994 239623 374000 239675
rect 381520 239623 381526 239675
rect 381578 239663 381584 239675
rect 388912 239663 388918 239675
rect 381578 239635 388918 239663
rect 381578 239623 381584 239635
rect 388912 239623 388918 239635
rect 388970 239623 388976 239675
rect 396112 239623 396118 239675
rect 396170 239663 396176 239675
rect 541648 239663 541654 239675
rect 396170 239635 541654 239663
rect 396170 239623 396176 239635
rect 541648 239623 541654 239635
rect 541706 239623 541712 239675
rect 288112 239549 288118 239601
rect 288170 239589 288176 239601
rect 289408 239589 289414 239601
rect 288170 239561 289414 239589
rect 288170 239549 288176 239561
rect 289408 239549 289414 239561
rect 289466 239549 289472 239601
rect 409264 239589 409270 239601
rect 289570 239561 409270 239589
rect 288208 239475 288214 239527
rect 288266 239515 288272 239527
rect 289570 239515 289598 239561
rect 409264 239549 409270 239561
rect 409322 239549 409328 239601
rect 409456 239549 409462 239601
rect 409514 239589 409520 239601
rect 414544 239589 414550 239601
rect 409514 239561 414550 239589
rect 409514 239549 409520 239561
rect 414544 239549 414550 239561
rect 414602 239549 414608 239601
rect 437776 239549 437782 239601
rect 437834 239589 437840 239601
rect 443728 239589 443734 239601
rect 437834 239561 443734 239589
rect 437834 239549 437840 239561
rect 443728 239549 443734 239561
rect 443786 239549 443792 239601
rect 443968 239549 443974 239601
rect 444026 239589 444032 239601
rect 454000 239589 454006 239601
rect 444026 239561 454006 239589
rect 444026 239549 444032 239561
rect 454000 239549 454006 239561
rect 454058 239549 454064 239601
rect 288266 239487 289598 239515
rect 288266 239475 288272 239487
rect 291184 239475 291190 239527
rect 291242 239515 291248 239527
rect 381520 239515 381526 239527
rect 291242 239487 381526 239515
rect 291242 239475 291248 239487
rect 381520 239475 381526 239487
rect 381578 239475 381584 239527
rect 401872 239475 401878 239527
rect 401930 239515 401936 239527
rect 401930 239487 406526 239515
rect 401930 239475 401936 239487
rect 348418 239413 381566 239441
rect 293104 239253 293110 239305
rect 293162 239293 293168 239305
rect 348418 239293 348446 239413
rect 381538 239367 381566 239413
rect 401392 239401 401398 239453
rect 401450 239441 401456 239453
rect 406384 239441 406390 239453
rect 401450 239413 406390 239441
rect 401450 239401 401456 239413
rect 406384 239401 406390 239413
rect 406442 239401 406448 239453
rect 406498 239441 406526 239487
rect 406576 239475 406582 239527
rect 406634 239515 406640 239527
rect 408880 239515 408886 239527
rect 406634 239487 408886 239515
rect 406634 239475 406640 239487
rect 408880 239475 408886 239487
rect 408938 239475 408944 239527
rect 410320 239475 410326 239527
rect 410378 239515 410384 239527
rect 410378 239487 410846 239515
rect 410378 239475 410384 239487
rect 410818 239441 410846 239487
rect 410992 239475 410998 239527
rect 411050 239515 411056 239527
rect 411568 239515 411574 239527
rect 411050 239487 411574 239515
rect 411050 239475 411056 239487
rect 411568 239475 411574 239487
rect 411626 239475 411632 239527
rect 412048 239475 412054 239527
rect 412106 239515 412112 239527
rect 445264 239515 445270 239527
rect 412106 239487 445270 239515
rect 412106 239475 412112 239487
rect 445264 239475 445270 239487
rect 445322 239475 445328 239527
rect 444400 239441 444406 239453
rect 406498 239413 410366 239441
rect 410818 239413 444406 239441
rect 381538 239339 402014 239367
rect 293162 239265 348446 239293
rect 293162 239253 293168 239265
rect 388912 239253 388918 239305
rect 388970 239293 388976 239305
rect 401872 239293 401878 239305
rect 388970 239265 401878 239293
rect 388970 239253 388976 239265
rect 401872 239253 401878 239265
rect 401930 239253 401936 239305
rect 401986 239293 402014 239339
rect 405328 239327 405334 239379
rect 405386 239367 405392 239379
rect 410224 239367 410230 239379
rect 405386 239339 410230 239367
rect 405386 239327 405392 239339
rect 410224 239327 410230 239339
rect 410282 239327 410288 239379
rect 410338 239367 410366 239413
rect 444400 239401 444406 239413
rect 444458 239401 444464 239453
rect 411088 239367 411094 239379
rect 410338 239339 411094 239367
rect 411088 239327 411094 239339
rect 411146 239327 411152 239379
rect 414064 239327 414070 239379
rect 414122 239367 414128 239379
rect 444112 239367 444118 239379
rect 414122 239339 444118 239367
rect 414122 239327 414128 239339
rect 444112 239327 444118 239339
rect 444170 239327 444176 239379
rect 446320 239327 446326 239379
rect 446378 239367 446384 239379
rect 447952 239367 447958 239379
rect 446378 239339 447958 239367
rect 446378 239327 446384 239339
rect 447952 239327 447958 239339
rect 448010 239327 448016 239379
rect 406576 239293 406582 239305
rect 401986 239265 406582 239293
rect 406576 239253 406582 239265
rect 406634 239253 406640 239305
rect 407536 239253 407542 239305
rect 407594 239293 407600 239305
rect 408880 239293 408886 239305
rect 407594 239265 408886 239293
rect 407594 239253 407600 239265
rect 408880 239253 408886 239265
rect 408938 239253 408944 239305
rect 412144 239253 412150 239305
rect 412202 239293 412208 239305
rect 444304 239293 444310 239305
rect 412202 239265 444310 239293
rect 412202 239253 412208 239265
rect 444304 239253 444310 239265
rect 444362 239253 444368 239305
rect 140368 239179 140374 239231
rect 140426 239219 140432 239231
rect 141136 239219 141142 239231
rect 140426 239191 141142 239219
rect 140426 239179 140432 239191
rect 141136 239179 141142 239191
rect 141194 239179 141200 239231
rect 288400 239179 288406 239231
rect 288458 239219 288464 239231
rect 406288 239219 406294 239231
rect 288458 239191 406294 239219
rect 288458 239179 288464 239191
rect 406288 239179 406294 239191
rect 406346 239179 406352 239231
rect 408496 239179 408502 239231
rect 408554 239219 408560 239231
rect 443536 239219 443542 239231
rect 408554 239191 443542 239219
rect 408554 239179 408560 239191
rect 443536 239179 443542 239191
rect 443594 239179 443600 239231
rect 149584 239105 149590 239157
rect 149642 239145 149648 239157
rect 155344 239145 155350 239157
rect 149642 239117 155350 239145
rect 149642 239105 149648 239117
rect 155344 239105 155350 239117
rect 155402 239105 155408 239157
rect 391312 239105 391318 239157
rect 391370 239145 391376 239157
rect 457936 239145 457942 239157
rect 391370 239117 457942 239145
rect 391370 239105 391376 239117
rect 457936 239105 457942 239117
rect 457994 239105 458000 239157
rect 144016 239031 144022 239083
rect 144074 239071 144080 239083
rect 188560 239071 188566 239083
rect 144074 239043 188566 239071
rect 144074 239031 144080 239043
rect 188560 239031 188566 239043
rect 188618 239031 188624 239083
rect 325456 239031 325462 239083
rect 325514 239071 325520 239083
rect 341584 239071 341590 239083
rect 325514 239043 341590 239071
rect 325514 239031 325520 239043
rect 341584 239031 341590 239043
rect 341642 239031 341648 239083
rect 345808 239031 345814 239083
rect 345866 239071 345872 239083
rect 365488 239071 365494 239083
rect 345866 239043 365494 239071
rect 345866 239031 345872 239043
rect 365488 239031 365494 239043
rect 365546 239031 365552 239083
rect 391696 239031 391702 239083
rect 391754 239071 391760 239083
rect 392656 239071 392662 239083
rect 391754 239043 392662 239071
rect 391754 239031 391760 239043
rect 392656 239031 392662 239043
rect 392714 239031 392720 239083
rect 397456 239031 397462 239083
rect 397514 239071 397520 239083
rect 413680 239071 413686 239083
rect 397514 239043 413686 239071
rect 397514 239031 397520 239043
rect 413680 239031 413686 239043
rect 413738 239031 413744 239083
rect 413872 239031 413878 239083
rect 413930 239071 413936 239083
rect 419632 239071 419638 239083
rect 413930 239043 419638 239071
rect 413930 239031 413936 239043
rect 419632 239031 419638 239043
rect 419690 239031 419696 239083
rect 146896 238957 146902 239009
rect 146954 238997 146960 239009
rect 149776 238997 149782 239009
rect 146954 238969 149782 238997
rect 146954 238957 146960 238969
rect 149776 238957 149782 238969
rect 149834 238957 149840 239009
rect 218704 238957 218710 239009
rect 218762 238997 218768 239009
rect 342736 238997 342742 239009
rect 218762 238969 342742 238997
rect 218762 238957 218768 238969
rect 342736 238957 342742 238969
rect 342794 238957 342800 239009
rect 344272 238957 344278 239009
rect 344330 238997 344336 239009
rect 354736 238997 354742 239009
rect 344330 238969 354742 238997
rect 344330 238957 344336 238969
rect 354736 238957 354742 238969
rect 354794 238957 354800 239009
rect 354832 238957 354838 239009
rect 354890 238997 354896 239009
rect 518416 238997 518422 239009
rect 354890 238969 518422 238997
rect 354890 238957 354896 238969
rect 518416 238957 518422 238969
rect 518474 238957 518480 239009
rect 227344 238883 227350 238935
rect 227402 238923 227408 238935
rect 349360 238923 349366 238935
rect 227402 238895 349366 238923
rect 227402 238883 227408 238895
rect 349360 238883 349366 238895
rect 349418 238883 349424 238935
rect 350704 238883 350710 238935
rect 350762 238923 350768 238935
rect 353200 238923 353206 238935
rect 350762 238895 353206 238923
rect 350762 238883 350768 238895
rect 353200 238883 353206 238895
rect 353258 238883 353264 238935
rect 354448 238923 354454 238935
rect 354370 238895 354454 238923
rect 283888 238809 283894 238861
rect 283946 238849 283952 238861
rect 340144 238849 340150 238861
rect 283946 238821 340150 238849
rect 283946 238809 283952 238821
rect 340144 238809 340150 238821
rect 340202 238809 340208 238861
rect 342736 238809 342742 238861
rect 342794 238849 342800 238861
rect 345328 238849 345334 238861
rect 342794 238821 345334 238849
rect 342794 238809 342800 238821
rect 345328 238809 345334 238821
rect 345386 238809 345392 238861
rect 346864 238809 346870 238861
rect 346922 238849 346928 238861
rect 354370 238849 354398 238895
rect 354448 238883 354454 238895
rect 354506 238883 354512 238935
rect 354544 238883 354550 238935
rect 354602 238923 354608 238935
rect 512944 238923 512950 238935
rect 354602 238895 512950 238923
rect 354602 238883 354608 238895
rect 512944 238883 512950 238895
rect 513002 238883 513008 238935
rect 501232 238849 501238 238861
rect 346922 238821 354398 238849
rect 354562 238821 501238 238849
rect 346922 238809 346928 238821
rect 140560 238735 140566 238787
rect 140618 238775 140624 238787
rect 140944 238775 140950 238787
rect 140618 238747 140950 238775
rect 140618 238735 140624 238747
rect 140944 238735 140950 238747
rect 141002 238735 141008 238787
rect 289552 238735 289558 238787
rect 289610 238775 289616 238787
rect 354352 238775 354358 238787
rect 289610 238747 354358 238775
rect 289610 238735 289616 238747
rect 354352 238735 354358 238747
rect 354410 238735 354416 238787
rect 354448 238735 354454 238787
rect 354506 238775 354512 238787
rect 354562 238775 354590 238821
rect 501232 238809 501238 238821
rect 501290 238809 501296 238861
rect 354506 238747 354590 238775
rect 358498 238747 358718 238775
rect 354506 238735 354512 238747
rect 283696 238661 283702 238713
rect 283754 238701 283760 238713
rect 339472 238701 339478 238713
rect 283754 238673 339478 238701
rect 283754 238661 283760 238673
rect 339472 238661 339478 238673
rect 339530 238661 339536 238713
rect 346480 238661 346486 238713
rect 346538 238701 346544 238713
rect 358498 238701 358526 238747
rect 346538 238673 358526 238701
rect 358690 238701 358718 238747
rect 359152 238735 359158 238787
rect 359210 238775 359216 238787
rect 507088 238775 507094 238787
rect 359210 238747 507094 238775
rect 359210 238735 359216 238747
rect 507088 238735 507094 238747
rect 507146 238735 507152 238787
rect 495472 238701 495478 238713
rect 358690 238673 495478 238701
rect 346538 238661 346544 238673
rect 495472 238661 495478 238673
rect 495530 238661 495536 238713
rect 285040 238587 285046 238639
rect 285098 238627 285104 238639
rect 337168 238627 337174 238639
rect 285098 238599 337174 238627
rect 285098 238587 285104 238599
rect 337168 238587 337174 238599
rect 337226 238587 337232 238639
rect 337264 238587 337270 238639
rect 337322 238627 337328 238639
rect 358480 238627 358486 238639
rect 337322 238599 358486 238627
rect 337322 238587 337328 238599
rect 358480 238587 358486 238599
rect 358538 238587 358544 238639
rect 360496 238587 360502 238639
rect 360554 238627 360560 238639
rect 501328 238627 501334 238639
rect 360554 238599 501334 238627
rect 360554 238587 360560 238599
rect 501328 238587 501334 238599
rect 501386 238587 501392 238639
rect 42160 238513 42166 238565
rect 42218 238553 42224 238565
rect 42352 238553 42358 238565
rect 42218 238525 42358 238553
rect 42218 238513 42224 238525
rect 42352 238513 42358 238525
rect 42410 238513 42416 238565
rect 287056 238513 287062 238565
rect 287114 238553 287120 238565
rect 340528 238553 340534 238565
rect 287114 238525 340534 238553
rect 287114 238513 287120 238525
rect 340528 238513 340534 238525
rect 340586 238513 340592 238565
rect 346096 238513 346102 238565
rect 346154 238553 346160 238565
rect 486832 238553 486838 238565
rect 346154 238525 486838 238553
rect 346154 238513 346160 238525
rect 486832 238513 486838 238525
rect 486890 238513 486896 238565
rect 42544 238439 42550 238491
rect 42602 238439 42608 238491
rect 286576 238439 286582 238491
rect 286634 238479 286640 238491
rect 339856 238479 339862 238491
rect 286634 238451 339862 238479
rect 286634 238439 286640 238451
rect 339856 238439 339862 238451
rect 339914 238439 339920 238491
rect 345712 238439 345718 238491
rect 345770 238479 345776 238491
rect 481168 238479 481174 238491
rect 345770 238451 481174 238479
rect 345770 238439 345776 238451
rect 481168 238439 481174 238451
rect 481226 238439 481232 238491
rect 42352 238365 42358 238417
rect 42410 238405 42416 238417
rect 42562 238405 42590 238439
rect 42410 238377 42590 238405
rect 42410 238365 42416 238377
rect 286864 238365 286870 238417
rect 286922 238405 286928 238417
rect 340912 238405 340918 238417
rect 286922 238377 340918 238405
rect 286922 238365 286928 238377
rect 340912 238365 340918 238377
rect 340970 238365 340976 238417
rect 341008 238365 341014 238417
rect 341066 238405 341072 238417
rect 362128 238405 362134 238417
rect 341066 238377 362134 238405
rect 341066 238365 341072 238377
rect 362128 238365 362134 238377
rect 362186 238365 362192 238417
rect 390160 238365 390166 238417
rect 390218 238405 390224 238417
rect 407824 238405 407830 238417
rect 390218 238377 407830 238405
rect 390218 238365 390224 238377
rect 407824 238365 407830 238377
rect 407882 238365 407888 238417
rect 408016 238365 408022 238417
rect 408074 238405 408080 238417
rect 410992 238405 410998 238417
rect 408074 238377 410998 238405
rect 408074 238365 408080 238377
rect 410992 238365 410998 238377
rect 411050 238365 411056 238417
rect 411280 238365 411286 238417
rect 411338 238405 411344 238417
rect 541456 238405 541462 238417
rect 411338 238377 541462 238405
rect 411338 238365 411344 238377
rect 541456 238365 541462 238377
rect 541514 238365 541520 238417
rect 286768 238291 286774 238343
rect 286826 238331 286832 238343
rect 387280 238331 387286 238343
rect 286826 238303 387286 238331
rect 286826 238291 286832 238303
rect 387280 238291 387286 238303
rect 387338 238291 387344 238343
rect 392848 238291 392854 238343
rect 392906 238331 392912 238343
rect 405904 238331 405910 238343
rect 392906 238303 405910 238331
rect 392906 238291 392912 238303
rect 405904 238291 405910 238303
rect 405962 238291 405968 238343
rect 406096 238291 406102 238343
rect 406154 238331 406160 238343
rect 532912 238331 532918 238343
rect 406154 238303 532918 238331
rect 406154 238291 406160 238303
rect 532912 238291 532918 238303
rect 532970 238291 532976 238343
rect 286000 238217 286006 238269
rect 286058 238257 286064 238269
rect 339088 238257 339094 238269
rect 286058 238229 339094 238257
rect 286058 238217 286064 238229
rect 339088 238217 339094 238229
rect 339146 238217 339152 238269
rect 344944 238217 344950 238269
rect 345002 238257 345008 238269
rect 469456 238257 469462 238269
rect 345002 238229 469462 238257
rect 345002 238217 345008 238229
rect 469456 238217 469462 238229
rect 469514 238217 469520 238269
rect 285232 238143 285238 238195
rect 285290 238183 285296 238195
rect 345616 238183 345622 238195
rect 285290 238155 345622 238183
rect 285290 238143 285296 238155
rect 345616 238143 345622 238155
rect 345674 238143 345680 238195
rect 402640 238143 402646 238195
rect 402698 238183 402704 238195
rect 403120 238183 403126 238195
rect 402698 238155 403126 238183
rect 402698 238143 402704 238155
rect 403120 238143 403126 238155
rect 403178 238143 403184 238195
rect 403216 238143 403222 238195
rect 403274 238183 403280 238195
rect 527248 238183 527254 238195
rect 403274 238155 527254 238183
rect 403274 238143 403280 238155
rect 527248 238143 527254 238155
rect 527306 238143 527312 238195
rect 305314 238081 325406 238109
rect 305104 237995 305110 238047
rect 305162 238035 305168 238047
rect 305314 238035 305342 238081
rect 305162 238007 305342 238035
rect 325378 238035 325406 238081
rect 337168 238069 337174 238121
rect 337226 238109 337232 238121
rect 341104 238109 341110 238121
rect 337226 238081 341110 238109
rect 337226 238069 337232 238081
rect 341104 238069 341110 238081
rect 341162 238069 341168 238121
rect 344656 238069 344662 238121
rect 344714 238109 344720 238121
rect 463696 238109 463702 238121
rect 344714 238081 345758 238109
rect 344714 238069 344720 238081
rect 345520 238035 345526 238047
rect 325378 238007 345526 238035
rect 305162 237995 305168 238007
rect 345520 237995 345526 238007
rect 345578 237995 345584 238047
rect 345730 238035 345758 238081
rect 345922 238081 463702 238109
rect 345922 238035 345950 238081
rect 463696 238069 463702 238081
rect 463754 238069 463760 238121
rect 345730 238007 345950 238035
rect 365680 237995 365686 238047
rect 365738 238035 365744 238047
rect 390160 238035 390166 238047
rect 365738 238007 390166 238035
rect 365738 237995 365744 238007
rect 390160 237995 390166 238007
rect 390218 237995 390224 238047
rect 393904 237995 393910 238047
rect 393962 238035 393968 238047
rect 504016 238035 504022 238047
rect 393962 238007 504022 238035
rect 393962 237995 393968 238007
rect 504016 237995 504022 238007
rect 504074 237995 504080 238047
rect 288016 237921 288022 237973
rect 288074 237961 288080 237973
rect 350704 237961 350710 237973
rect 288074 237933 350710 237961
rect 288074 237921 288080 237933
rect 350704 237921 350710 237933
rect 350762 237921 350768 237973
rect 350800 237921 350806 237973
rect 350858 237961 350864 237973
rect 361456 237961 361462 237973
rect 350858 237933 361462 237961
rect 350858 237921 350864 237933
rect 361456 237921 361462 237933
rect 361514 237921 361520 237973
rect 366352 237921 366358 237973
rect 366410 237961 366416 237973
rect 485488 237961 485494 237973
rect 366410 237933 485494 237961
rect 366410 237921 366416 237933
rect 485488 237921 485494 237933
rect 485546 237921 485552 237973
rect 288304 237847 288310 237899
rect 288362 237887 288368 237899
rect 325552 237887 325558 237899
rect 288362 237859 325558 237887
rect 288362 237847 288368 237859
rect 325552 237847 325558 237859
rect 325610 237847 325616 237899
rect 325936 237847 325942 237899
rect 325994 237887 326000 237899
rect 398896 237887 398902 237899
rect 325994 237859 398902 237887
rect 325994 237847 326000 237859
rect 398896 237847 398902 237859
rect 398954 237847 398960 237899
rect 406000 237887 406006 237899
rect 399010 237859 406006 237887
rect 282544 237773 282550 237825
rect 282602 237813 282608 237825
rect 399010 237813 399038 237859
rect 406000 237847 406006 237859
rect 406058 237847 406064 237899
rect 408976 237847 408982 237899
rect 409034 237887 409040 237899
rect 430576 237887 430582 237899
rect 409034 237859 430582 237887
rect 409034 237847 409040 237859
rect 430576 237847 430582 237859
rect 430634 237847 430640 237899
rect 435088 237847 435094 237899
rect 435146 237887 435152 237899
rect 533008 237887 533014 237899
rect 435146 237859 533014 237887
rect 435146 237847 435152 237859
rect 533008 237847 533014 237859
rect 533066 237847 533072 237899
rect 282602 237785 399038 237813
rect 282602 237773 282608 237785
rect 399472 237773 399478 237825
rect 399530 237813 399536 237825
rect 419056 237813 419062 237825
rect 399530 237785 419062 237813
rect 399530 237773 399536 237785
rect 419056 237773 419062 237785
rect 419114 237773 419120 237825
rect 436816 237773 436822 237825
rect 436874 237813 436880 237825
rect 541552 237813 541558 237825
rect 436874 237785 541558 237813
rect 436874 237773 436880 237785
rect 541552 237773 541558 237785
rect 541610 237773 541616 237825
rect 42160 237699 42166 237751
rect 42218 237739 42224 237751
rect 50416 237739 50422 237751
rect 42218 237711 50422 237739
rect 42218 237699 42224 237711
rect 50416 237699 50422 237711
rect 50474 237699 50480 237751
rect 287920 237699 287926 237751
rect 287978 237739 287984 237751
rect 350800 237739 350806 237751
rect 287978 237711 350806 237739
rect 287978 237699 287984 237711
rect 350800 237699 350806 237711
rect 350858 237699 350864 237751
rect 350896 237699 350902 237751
rect 350954 237739 350960 237751
rect 477808 237739 477814 237751
rect 350954 237711 477814 237739
rect 350954 237699 350960 237711
rect 477808 237699 477814 237711
rect 477866 237699 477872 237751
rect 350128 237625 350134 237677
rect 350186 237665 350192 237677
rect 477424 237665 477430 237677
rect 350186 237637 477430 237665
rect 350186 237625 350192 237637
rect 477424 237625 477430 237637
rect 477482 237625 477488 237677
rect 140848 237551 140854 237603
rect 140906 237591 140912 237603
rect 140906 237563 140990 237591
rect 140906 237551 140912 237563
rect 140962 237381 140990 237563
rect 287344 237551 287350 237603
rect 287402 237591 287408 237603
rect 287402 237563 328190 237591
rect 287402 237551 287408 237563
rect 328162 237443 328190 237563
rect 331408 237551 331414 237603
rect 331466 237591 331472 237603
rect 338512 237591 338518 237603
rect 331466 237563 338518 237591
rect 331466 237551 331472 237563
rect 338512 237551 338518 237563
rect 338570 237551 338576 237603
rect 351568 237551 351574 237603
rect 351626 237591 351632 237603
rect 478192 237591 478198 237603
rect 351626 237563 478198 237591
rect 351626 237551 351632 237563
rect 478192 237551 478198 237563
rect 478250 237551 478256 237603
rect 334672 237477 334678 237529
rect 334730 237517 334736 237529
rect 449392 237517 449398 237529
rect 334730 237489 449398 237517
rect 334730 237477 334736 237489
rect 449392 237477 449398 237489
rect 449450 237477 449456 237529
rect 328162 237415 328478 237443
rect 140944 237329 140950 237381
rect 141002 237329 141008 237381
rect 328450 237073 328478 237415
rect 332080 237403 332086 237455
rect 332138 237443 332144 237455
rect 446800 237443 446806 237455
rect 332138 237415 446806 237443
rect 332138 237403 332144 237415
rect 446800 237403 446806 237415
rect 446858 237403 446864 237455
rect 332464 237329 332470 237381
rect 332522 237369 332528 237381
rect 447280 237369 447286 237381
rect 332522 237341 447286 237369
rect 332522 237329 332528 237341
rect 447280 237329 447286 237341
rect 447338 237329 447344 237381
rect 335440 237255 335446 237307
rect 335498 237295 335504 237307
rect 450256 237295 450262 237307
rect 335498 237267 450262 237295
rect 335498 237255 335504 237267
rect 450256 237255 450262 237267
rect 450314 237255 450320 237307
rect 336112 237181 336118 237233
rect 336170 237221 336176 237233
rect 450832 237221 450838 237233
rect 336170 237193 450838 237221
rect 336170 237181 336176 237193
rect 450832 237181 450838 237193
rect 450890 237181 450896 237233
rect 333232 237107 333238 237159
rect 333290 237147 333296 237159
rect 448048 237147 448054 237159
rect 333290 237119 448054 237147
rect 333290 237107 333296 237119
rect 448048 237107 448054 237119
rect 448106 237107 448112 237159
rect 356272 237073 356278 237085
rect 328450 237045 356278 237073
rect 356272 237033 356278 237045
rect 356330 237033 356336 237085
rect 358480 237033 358486 237085
rect 358538 237073 358544 237085
rect 451792 237073 451798 237085
rect 358538 237045 451798 237073
rect 358538 237033 358544 237045
rect 451792 237033 451798 237045
rect 451850 237033 451856 237085
rect 287632 236959 287638 237011
rect 287690 236999 287696 237011
rect 364720 236999 364726 237011
rect 287690 236971 364726 236999
rect 287690 236959 287696 236971
rect 364720 236959 364726 236971
rect 364778 236959 364784 237011
rect 398128 236959 398134 237011
rect 398186 236999 398192 237011
rect 460816 236999 460822 237011
rect 398186 236971 460822 236999
rect 398186 236959 398192 236971
rect 460816 236959 460822 236971
rect 460874 236959 460880 237011
rect 285808 236885 285814 236937
rect 285866 236925 285872 236937
rect 365296 236925 365302 236937
rect 285866 236897 365302 236925
rect 285866 236885 285872 236897
rect 365296 236885 365302 236897
rect 365354 236885 365360 236937
rect 397264 236885 397270 236937
rect 397322 236925 397328 236937
rect 453808 236925 453814 236937
rect 397322 236897 453814 236925
rect 397322 236885 397328 236897
rect 453808 236885 453814 236897
rect 453866 236885 453872 236937
rect 284848 236811 284854 236863
rect 284906 236851 284912 236863
rect 358096 236851 358102 236863
rect 284906 236823 358102 236851
rect 284906 236811 284912 236823
rect 358096 236811 358102 236823
rect 358154 236811 358160 236863
rect 398800 236811 398806 236863
rect 398858 236851 398864 236863
rect 418960 236851 418966 236863
rect 398858 236823 418966 236851
rect 398858 236811 398864 236823
rect 418960 236811 418966 236823
rect 419018 236811 419024 236863
rect 419056 236811 419062 236863
rect 419114 236851 419120 236863
rect 454960 236851 454966 236863
rect 419114 236823 454966 236851
rect 419114 236811 419120 236823
rect 454960 236811 454966 236823
rect 455018 236811 455024 236863
rect 285136 236737 285142 236789
rect 285194 236777 285200 236789
rect 341008 236777 341014 236789
rect 285194 236749 341014 236777
rect 285194 236737 285200 236749
rect 341008 236737 341014 236749
rect 341066 236737 341072 236789
rect 341104 236737 341110 236789
rect 341162 236777 341168 236789
rect 341162 236749 352094 236777
rect 341162 236737 341168 236749
rect 42160 236663 42166 236715
rect 42218 236703 42224 236715
rect 43120 236703 43126 236715
rect 42218 236675 43126 236703
rect 42218 236663 42224 236675
rect 43120 236663 43126 236675
rect 43178 236663 43184 236715
rect 351952 236703 351958 236715
rect 338242 236675 351958 236703
rect 287728 236589 287734 236641
rect 287786 236629 287792 236641
rect 338242 236629 338270 236675
rect 351952 236663 351958 236675
rect 352010 236663 352016 236715
rect 352066 236703 352094 236749
rect 354736 236737 354742 236789
rect 354794 236777 354800 236789
rect 455440 236777 455446 236789
rect 354794 236749 455446 236777
rect 354794 236737 354800 236749
rect 455440 236737 455446 236749
rect 455498 236737 455504 236789
rect 355504 236703 355510 236715
rect 352066 236675 355510 236703
rect 355504 236663 355510 236675
rect 355562 236663 355568 236715
rect 398896 236663 398902 236715
rect 398954 236703 398960 236715
rect 409072 236703 409078 236715
rect 398954 236675 409078 236703
rect 398954 236663 398960 236675
rect 409072 236663 409078 236675
rect 409130 236663 409136 236715
rect 409168 236663 409174 236715
rect 409226 236703 409232 236715
rect 413872 236703 413878 236715
rect 409226 236675 413878 236703
rect 409226 236663 409232 236675
rect 413872 236663 413878 236675
rect 413930 236663 413936 236715
rect 430288 236703 430294 236715
rect 414082 236675 430294 236703
rect 360592 236629 360598 236641
rect 287786 236601 338270 236629
rect 338338 236601 360598 236629
rect 287786 236589 287792 236601
rect 144016 236515 144022 236567
rect 144074 236555 144080 236567
rect 148816 236555 148822 236567
rect 144074 236527 148822 236555
rect 144074 236515 144080 236527
rect 148816 236515 148822 236527
rect 148874 236515 148880 236567
rect 287824 236515 287830 236567
rect 287882 236555 287888 236567
rect 338338 236555 338366 236601
rect 360592 236589 360598 236601
rect 360650 236589 360656 236641
rect 398992 236589 398998 236641
rect 399050 236629 399056 236641
rect 414082 236629 414110 236675
rect 430288 236663 430294 236675
rect 430346 236663 430352 236715
rect 433264 236663 433270 236715
rect 433322 236703 433328 236715
rect 440176 236703 440182 236715
rect 433322 236675 440182 236703
rect 433322 236663 433328 236675
rect 440176 236663 440182 236675
rect 440234 236663 440240 236715
rect 399050 236601 414110 236629
rect 399050 236589 399056 236601
rect 418960 236589 418966 236641
rect 419018 236629 419024 236641
rect 453424 236629 453430 236641
rect 419018 236601 453430 236629
rect 419018 236589 419024 236601
rect 453424 236589 453430 236601
rect 453482 236589 453488 236641
rect 287882 236527 338366 236555
rect 287882 236515 287888 236527
rect 338416 236515 338422 236567
rect 338474 236555 338480 236567
rect 359248 236555 359254 236567
rect 338474 236527 359254 236555
rect 338474 236515 338480 236527
rect 359248 236515 359254 236527
rect 359306 236515 359312 236567
rect 389200 236515 389206 236567
rect 389258 236555 389264 236567
rect 399184 236555 399190 236567
rect 389258 236527 399190 236555
rect 389258 236515 389264 236527
rect 399184 236515 399190 236527
rect 399242 236515 399248 236567
rect 400336 236515 400342 236567
rect 400394 236555 400400 236567
rect 479632 236555 479638 236567
rect 400394 236527 479638 236555
rect 400394 236515 400400 236527
rect 479632 236515 479638 236527
rect 479690 236515 479696 236567
rect 287248 236441 287254 236493
rect 287306 236481 287312 236493
rect 357424 236481 357430 236493
rect 287306 236453 357430 236481
rect 287306 236441 287312 236453
rect 357424 236441 357430 236453
rect 357482 236441 357488 236493
rect 397840 236441 397846 236493
rect 397898 236481 397904 236493
rect 399952 236481 399958 236493
rect 397898 236453 399958 236481
rect 397898 236441 397904 236453
rect 399952 236441 399958 236453
rect 400010 236441 400016 236493
rect 400048 236441 400054 236493
rect 400106 236481 400112 236493
rect 479248 236481 479254 236493
rect 400106 236453 479254 236481
rect 400106 236441 400112 236453
rect 479248 236441 479254 236453
rect 479306 236441 479312 236493
rect 287536 236367 287542 236419
rect 287594 236407 287600 236419
rect 338224 236407 338230 236419
rect 287594 236379 338230 236407
rect 287594 236367 287600 236379
rect 338224 236367 338230 236379
rect 338282 236367 338288 236419
rect 338320 236367 338326 236419
rect 338378 236407 338384 236419
rect 359632 236407 359638 236419
rect 338378 236379 359638 236407
rect 338378 236367 338384 236379
rect 359632 236367 359638 236379
rect 359690 236367 359696 236419
rect 360112 236367 360118 236419
rect 360170 236407 360176 236419
rect 377296 236407 377302 236419
rect 360170 236379 377302 236407
rect 360170 236367 360176 236379
rect 377296 236367 377302 236379
rect 377354 236367 377360 236419
rect 398704 236367 398710 236419
rect 398762 236407 398768 236419
rect 478864 236407 478870 236419
rect 398762 236379 478870 236407
rect 398762 236367 398768 236379
rect 478864 236367 478870 236379
rect 478922 236367 478928 236419
rect 296560 236293 296566 236345
rect 296618 236333 296624 236345
rect 296618 236305 345662 236333
rect 296618 236293 296624 236305
rect 345634 236271 345662 236305
rect 351952 236293 351958 236345
rect 352010 236333 352016 236345
rect 352010 236305 356126 236333
rect 352010 236293 352016 236305
rect 287440 236219 287446 236271
rect 287498 236259 287504 236271
rect 338320 236259 338326 236271
rect 287498 236231 338326 236259
rect 287498 236219 287504 236231
rect 338320 236219 338326 236231
rect 338378 236219 338384 236271
rect 345616 236219 345622 236271
rect 345674 236219 345680 236271
rect 356098 236259 356126 236305
rect 357040 236293 357046 236345
rect 357098 236333 357104 236345
rect 396496 236333 396502 236345
rect 357098 236305 396502 236333
rect 357098 236293 357104 236305
rect 396496 236293 396502 236305
rect 396554 236293 396560 236345
rect 398896 236293 398902 236345
rect 398954 236333 398960 236345
rect 478480 236333 478486 236345
rect 398954 236305 478486 236333
rect 398954 236293 398960 236305
rect 478480 236293 478486 236305
rect 478538 236293 478544 236345
rect 360304 236259 360310 236271
rect 356098 236231 360310 236259
rect 360304 236219 360310 236231
rect 360362 236219 360368 236271
rect 360400 236219 360406 236271
rect 360458 236259 360464 236271
rect 377104 236259 377110 236271
rect 360458 236231 377110 236259
rect 360458 236219 360464 236231
rect 377104 236219 377110 236231
rect 377162 236219 377168 236271
rect 397744 236219 397750 236271
rect 397802 236259 397808 236271
rect 482608 236259 482614 236271
rect 397802 236231 482614 236259
rect 397802 236219 397808 236231
rect 482608 236219 482614 236231
rect 482666 236219 482672 236271
rect 140176 236145 140182 236197
rect 140234 236185 140240 236197
rect 141232 236185 141238 236197
rect 140234 236157 141238 236185
rect 140234 236145 140240 236157
rect 141232 236145 141238 236157
rect 141290 236145 141296 236197
rect 287152 236145 287158 236197
rect 287210 236185 287216 236197
rect 355216 236185 355222 236197
rect 287210 236157 355222 236185
rect 287210 236145 287216 236157
rect 355216 236145 355222 236157
rect 355274 236145 355280 236197
rect 390160 236145 390166 236197
rect 390218 236185 390224 236197
rect 399472 236185 399478 236197
rect 390218 236157 399478 236185
rect 390218 236145 390224 236157
rect 399472 236145 399478 236157
rect 399530 236145 399536 236197
rect 399952 236145 399958 236197
rect 400010 236185 400016 236197
rect 400010 236157 400190 236185
rect 400010 236145 400016 236157
rect 218800 236071 218806 236123
rect 218858 236111 218864 236123
rect 298192 236111 298198 236123
rect 218858 236083 298198 236111
rect 218858 236071 218864 236083
rect 298192 236071 298198 236083
rect 298250 236071 298256 236123
rect 327280 236071 327286 236123
rect 327338 236111 327344 236123
rect 353584 236111 353590 236123
rect 327338 236083 353590 236111
rect 327338 236071 327344 236083
rect 353584 236071 353590 236083
rect 353642 236071 353648 236123
rect 353776 236071 353782 236123
rect 353834 236111 353840 236123
rect 400048 236111 400054 236123
rect 353834 236083 400054 236111
rect 353834 236071 353840 236083
rect 400048 236071 400054 236083
rect 400106 236071 400112 236123
rect 400162 236111 400190 236157
rect 400240 236145 400246 236197
rect 400298 236185 400304 236197
rect 482896 236185 482902 236197
rect 400298 236157 482902 236185
rect 400298 236145 400304 236157
rect 482896 236145 482902 236157
rect 482954 236145 482960 236197
rect 404464 236111 404470 236123
rect 400162 236083 404470 236111
rect 404464 236071 404470 236083
rect 404522 236071 404528 236123
rect 404560 236071 404566 236123
rect 404618 236111 404624 236123
rect 451984 236111 451990 236123
rect 404618 236083 451990 236111
rect 404618 236071 404624 236083
rect 451984 236071 451990 236083
rect 452042 236071 452048 236123
rect 452176 236071 452182 236123
rect 452234 236111 452240 236123
rect 453520 236111 453526 236123
rect 452234 236083 453526 236111
rect 452234 236071 452240 236083
rect 453520 236071 453526 236083
rect 453578 236071 453584 236123
rect 453904 236071 453910 236123
rect 453962 236111 453968 236123
rect 501136 236111 501142 236123
rect 453962 236083 501142 236111
rect 453962 236071 453968 236083
rect 501136 236071 501142 236083
rect 501194 236071 501200 236123
rect 204304 235997 204310 236049
rect 204362 236037 204368 236049
rect 290128 236037 290134 236049
rect 204362 236009 290134 236037
rect 204362 235997 204368 236009
rect 290128 235997 290134 236009
rect 290186 235997 290192 236049
rect 324400 235997 324406 236049
rect 324458 236037 324464 236049
rect 338224 236037 338230 236049
rect 324458 236009 338230 236037
rect 324458 235997 324464 236009
rect 338224 235997 338230 236009
rect 338282 235997 338288 236049
rect 338320 235997 338326 236049
rect 338378 236037 338384 236049
rect 348880 236037 348886 236049
rect 338378 236009 348886 236037
rect 338378 235997 338384 236009
rect 348880 235997 348886 236009
rect 348938 235997 348944 236049
rect 354640 235997 354646 236049
rect 354698 236037 354704 236049
rect 400336 236037 400342 236049
rect 354698 236009 400342 236037
rect 354698 235997 354704 236009
rect 400336 235997 400342 236009
rect 400394 235997 400400 236049
rect 401680 235997 401686 236049
rect 401738 236037 401744 236049
rect 403792 236037 403798 236049
rect 401738 236009 403798 236037
rect 401738 235997 401744 236009
rect 403792 235997 403798 236009
rect 403850 235997 403856 236049
rect 403888 235997 403894 236049
rect 403946 236037 403952 236049
rect 414832 236037 414838 236049
rect 403946 236009 414838 236037
rect 403946 235997 403952 236009
rect 414832 235997 414838 236009
rect 414890 235997 414896 236049
rect 414928 235997 414934 236049
rect 414986 236037 414992 236049
rect 420304 236037 420310 236049
rect 414986 236009 420310 236037
rect 414986 235997 414992 236009
rect 420304 235997 420310 236009
rect 420362 235997 420368 236049
rect 420784 235997 420790 236049
rect 420842 236037 420848 236049
rect 430672 236037 430678 236049
rect 420842 236009 430678 236037
rect 420842 235997 420848 236009
rect 430672 235997 430678 236009
rect 430730 235997 430736 236049
rect 434416 235997 434422 236049
rect 434474 236037 434480 236049
rect 443632 236037 443638 236049
rect 434474 236009 443638 236037
rect 434474 235997 434480 236009
rect 443632 235997 443638 236009
rect 443690 235997 443696 236049
rect 444688 235997 444694 236049
rect 444746 236037 444752 236049
rect 494992 236037 494998 236049
rect 444746 236009 494998 236037
rect 444746 235997 444752 236009
rect 494992 235997 494998 236009
rect 495050 235997 495056 236049
rect 209968 235923 209974 235975
rect 210026 235963 210032 235975
rect 294160 235963 294166 235975
rect 210026 235935 294166 235963
rect 210026 235923 210032 235935
rect 294160 235923 294166 235935
rect 294218 235923 294224 235975
rect 325072 235923 325078 235975
rect 325130 235963 325136 235975
rect 374992 235963 374998 235975
rect 325130 235935 374998 235963
rect 325130 235923 325136 235935
rect 374992 235923 374998 235935
rect 375050 235923 375056 235975
rect 375088 235923 375094 235975
rect 375146 235963 375152 235975
rect 391504 235963 391510 235975
rect 375146 235935 391510 235963
rect 375146 235923 375152 235935
rect 391504 235923 391510 235935
rect 391562 235923 391568 235975
rect 398416 235923 398422 235975
rect 398474 235963 398480 235975
rect 400240 235963 400246 235975
rect 398474 235935 400246 235963
rect 398474 235923 398480 235935
rect 400240 235923 400246 235935
rect 400298 235923 400304 235975
rect 400528 235923 400534 235975
rect 400586 235963 400592 235975
rect 408784 235963 408790 235975
rect 400586 235935 408790 235963
rect 400586 235923 400592 235935
rect 408784 235923 408790 235935
rect 408842 235923 408848 235975
rect 408880 235923 408886 235975
rect 408938 235963 408944 235975
rect 413008 235963 413014 235975
rect 408938 235935 413014 235963
rect 408938 235923 408944 235935
rect 413008 235923 413014 235935
rect 413066 235923 413072 235975
rect 413104 235923 413110 235975
rect 413162 235963 413168 235975
rect 418480 235963 418486 235975
rect 413162 235935 418486 235963
rect 413162 235923 413168 235935
rect 418480 235923 418486 235935
rect 418538 235923 418544 235975
rect 418576 235923 418582 235975
rect 418634 235963 418640 235975
rect 420400 235963 420406 235975
rect 418634 235935 420406 235963
rect 418634 235923 418640 235935
rect 420400 235923 420406 235935
rect 420458 235923 420464 235975
rect 425104 235923 425110 235975
rect 425162 235963 425168 235975
rect 446320 235963 446326 235975
rect 425162 235935 446326 235963
rect 425162 235923 425168 235935
rect 446320 235923 446326 235935
rect 446378 235923 446384 235975
rect 446896 235923 446902 235975
rect 446954 235963 446960 235975
rect 497872 235963 497878 235975
rect 446954 235935 497878 235963
rect 446954 235923 446960 235935
rect 497872 235923 497878 235935
rect 497930 235923 497936 235975
rect 285424 235849 285430 235901
rect 285482 235889 285488 235901
rect 374320 235889 374326 235901
rect 285482 235861 374326 235889
rect 285482 235849 285488 235861
rect 374320 235849 374326 235861
rect 374378 235849 374384 235901
rect 374416 235849 374422 235901
rect 374474 235889 374480 235901
rect 377200 235889 377206 235901
rect 374474 235861 377206 235889
rect 374474 235849 374480 235861
rect 377200 235849 377206 235861
rect 377258 235849 377264 235901
rect 395728 235849 395734 235901
rect 395786 235889 395792 235901
rect 405424 235889 405430 235901
rect 395786 235861 405430 235889
rect 395786 235849 395792 235861
rect 405424 235849 405430 235861
rect 405482 235849 405488 235901
rect 409456 235889 409462 235901
rect 406018 235861 409462 235889
rect 285520 235775 285526 235827
rect 285578 235815 285584 235827
rect 378832 235815 378838 235827
rect 285578 235787 378838 235815
rect 285578 235775 285584 235787
rect 378832 235775 378838 235787
rect 378890 235775 378896 235827
rect 389104 235775 389110 235827
rect 389162 235815 389168 235827
rect 389162 235787 399038 235815
rect 389162 235775 389168 235787
rect 140080 235701 140086 235753
rect 140138 235741 140144 235753
rect 141520 235741 141526 235753
rect 140138 235713 141526 235741
rect 140138 235701 140144 235713
rect 141520 235701 141526 235713
rect 141578 235701 141584 235753
rect 224560 235701 224566 235753
rect 224618 235741 224624 235753
rect 302224 235741 302230 235753
rect 224618 235713 302230 235741
rect 224618 235701 224624 235713
rect 302224 235701 302230 235713
rect 302282 235701 302288 235753
rect 334288 235701 334294 235753
rect 334346 235741 334352 235753
rect 334346 235713 398942 235741
rect 334346 235701 334352 235713
rect 284368 235627 284374 235679
rect 284426 235667 284432 235679
rect 375088 235667 375094 235679
rect 284426 235639 375094 235667
rect 284426 235627 284432 235639
rect 375088 235627 375094 235639
rect 375146 235627 375152 235679
rect 375280 235627 375286 235679
rect 375338 235667 375344 235679
rect 398800 235667 398806 235679
rect 375338 235639 398806 235667
rect 375338 235627 375344 235639
rect 398800 235627 398806 235639
rect 398858 235627 398864 235679
rect 338224 235553 338230 235605
rect 338282 235593 338288 235605
rect 338704 235593 338710 235605
rect 338282 235565 338710 235593
rect 338282 235553 338288 235565
rect 338704 235553 338710 235565
rect 338762 235553 338768 235605
rect 338992 235553 338998 235605
rect 339050 235593 339056 235605
rect 346768 235593 346774 235605
rect 339050 235565 346774 235593
rect 339050 235553 339056 235565
rect 346768 235553 346774 235565
rect 346826 235553 346832 235605
rect 357040 235553 357046 235605
rect 357098 235593 357104 235605
rect 390160 235593 390166 235605
rect 357098 235565 390166 235593
rect 357098 235553 357104 235565
rect 390160 235553 390166 235565
rect 390218 235553 390224 235605
rect 398914 235593 398942 235713
rect 399010 235667 399038 235787
rect 399280 235775 399286 235827
rect 399338 235815 399344 235827
rect 406018 235815 406046 235861
rect 409456 235849 409462 235861
rect 409514 235849 409520 235901
rect 411760 235849 411766 235901
rect 411818 235889 411824 235901
rect 420496 235889 420502 235901
rect 411818 235861 420502 235889
rect 411818 235849 411824 235861
rect 420496 235849 420502 235861
rect 420554 235849 420560 235901
rect 420592 235849 420598 235901
rect 420650 235889 420656 235901
rect 441520 235889 441526 235901
rect 420650 235861 441526 235889
rect 420650 235849 420656 235861
rect 441520 235849 441526 235861
rect 441578 235849 441584 235901
rect 443248 235849 443254 235901
rect 443306 235889 443312 235901
rect 493744 235889 493750 235901
rect 443306 235861 493750 235889
rect 443306 235849 443312 235861
rect 493744 235849 493750 235861
rect 493802 235849 493808 235901
rect 399338 235787 406046 235815
rect 399338 235775 399344 235787
rect 406096 235775 406102 235827
rect 406154 235815 406160 235827
rect 435568 235815 435574 235827
rect 406154 235787 435574 235815
rect 406154 235775 406160 235787
rect 435568 235775 435574 235787
rect 435626 235775 435632 235827
rect 441808 235775 441814 235827
rect 441866 235815 441872 235827
rect 493552 235815 493558 235827
rect 441866 235787 493558 235815
rect 441866 235775 441872 235787
rect 493552 235775 493558 235787
rect 493610 235775 493616 235827
rect 399184 235701 399190 235753
rect 399242 235741 399248 235753
rect 420592 235741 420598 235753
rect 399242 235713 420598 235741
rect 399242 235701 399248 235713
rect 420592 235701 420598 235713
rect 420650 235701 420656 235753
rect 420784 235701 420790 235753
rect 420842 235741 420848 235753
rect 436432 235741 436438 235753
rect 420842 235713 436438 235741
rect 420842 235701 420848 235713
rect 436432 235701 436438 235713
rect 436490 235701 436496 235753
rect 440272 235701 440278 235753
rect 440330 235741 440336 235753
rect 494800 235741 494806 235753
rect 440330 235713 494806 235741
rect 440330 235701 440336 235713
rect 494800 235701 494806 235713
rect 494858 235701 494864 235753
rect 412624 235667 412630 235679
rect 399010 235639 412630 235667
rect 412624 235627 412630 235639
rect 412682 235627 412688 235679
rect 412720 235627 412726 235679
rect 412778 235667 412784 235679
rect 414640 235667 414646 235679
rect 412778 235639 414646 235667
rect 412778 235627 412784 235639
rect 414640 235627 414646 235639
rect 414698 235627 414704 235679
rect 414832 235627 414838 235679
rect 414890 235667 414896 235679
rect 420112 235667 420118 235679
rect 414890 235639 420118 235667
rect 414890 235627 414896 235639
rect 420112 235627 420118 235639
rect 420170 235627 420176 235679
rect 420880 235627 420886 235679
rect 420938 235667 420944 235679
rect 437776 235667 437782 235679
rect 420938 235639 437782 235667
rect 420938 235627 420944 235639
rect 437776 235627 437782 235639
rect 437834 235627 437840 235679
rect 438832 235627 438838 235679
rect 438890 235667 438896 235679
rect 494416 235667 494422 235679
rect 438890 235639 494422 235667
rect 438890 235627 438896 235639
rect 494416 235627 494422 235639
rect 494474 235627 494480 235679
rect 399184 235593 399190 235605
rect 398914 235565 399190 235593
rect 399184 235553 399190 235565
rect 399242 235553 399248 235605
rect 399472 235553 399478 235605
rect 399530 235593 399536 235605
rect 417616 235593 417622 235605
rect 399530 235565 417622 235593
rect 399530 235553 399536 235565
rect 417616 235553 417622 235565
rect 417674 235553 417680 235605
rect 424432 235553 424438 235605
rect 424490 235593 424496 235605
rect 431344 235593 431350 235605
rect 424490 235565 431350 235593
rect 424490 235553 424496 235565
rect 431344 235553 431350 235565
rect 431402 235553 431408 235605
rect 439120 235553 439126 235605
rect 439178 235593 439184 235605
rect 449776 235593 449782 235605
rect 439178 235565 449782 235593
rect 439178 235553 439184 235565
rect 449776 235553 449782 235565
rect 449834 235553 449840 235605
rect 449872 235553 449878 235605
rect 449930 235593 449936 235605
rect 506896 235593 506902 235605
rect 449930 235565 506902 235593
rect 449930 235553 449936 235565
rect 506896 235553 506902 235565
rect 506954 235553 506960 235605
rect 312976 235479 312982 235531
rect 313034 235519 313040 235531
rect 338320 235519 338326 235531
rect 313034 235491 338326 235519
rect 313034 235479 313040 235491
rect 338320 235479 338326 235491
rect 338378 235479 338384 235531
rect 353584 235479 353590 235531
rect 353642 235519 353648 235531
rect 360112 235519 360118 235531
rect 353642 235491 360118 235519
rect 353642 235479 353648 235491
rect 360112 235479 360118 235491
rect 360170 235479 360176 235531
rect 375280 235519 375286 235531
rect 360226 235491 375286 235519
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 43024 235445 43030 235457
rect 42218 235417 43030 235445
rect 42218 235405 42224 235417
rect 43024 235405 43030 235417
rect 43082 235405 43088 235457
rect 311536 235405 311542 235457
rect 311594 235445 311600 235457
rect 338608 235445 338614 235457
rect 311594 235417 338614 235445
rect 311594 235405 311600 235417
rect 338608 235405 338614 235417
rect 338666 235405 338672 235457
rect 338800 235405 338806 235457
rect 338858 235445 338864 235457
rect 360226 235445 360254 235491
rect 375280 235479 375286 235491
rect 375338 235479 375344 235531
rect 491728 235519 491734 235531
rect 378658 235491 491734 235519
rect 338858 235417 360254 235445
rect 338858 235405 338864 235417
rect 377008 235405 377014 235457
rect 377066 235445 377072 235457
rect 378658 235445 378686 235491
rect 491728 235479 491734 235491
rect 491786 235479 491792 235531
rect 377066 235417 378686 235445
rect 377066 235405 377072 235417
rect 382864 235405 382870 235457
rect 382922 235445 382928 235457
rect 497680 235445 497686 235457
rect 382922 235417 497686 235445
rect 382922 235405 382928 235417
rect 497680 235405 497686 235417
rect 497738 235405 497744 235457
rect 309328 235331 309334 235383
rect 309386 235371 309392 235383
rect 352144 235371 352150 235383
rect 309386 235343 352150 235371
rect 309386 235331 309392 235343
rect 352144 235331 352150 235343
rect 352202 235331 352208 235383
rect 356368 235331 356374 235383
rect 356426 235371 356432 235383
rect 360112 235371 360118 235383
rect 356426 235343 360118 235371
rect 356426 235331 356432 235343
rect 360112 235331 360118 235343
rect 360170 235331 360176 235383
rect 360400 235331 360406 235383
rect 360458 235371 360464 235383
rect 360688 235371 360694 235383
rect 360458 235343 360694 235371
rect 360458 235331 360464 235343
rect 360688 235331 360694 235343
rect 360746 235331 360752 235383
rect 379504 235371 379510 235383
rect 372610 235343 379510 235371
rect 328432 235257 328438 235309
rect 328490 235297 328496 235309
rect 338128 235297 338134 235309
rect 328490 235269 338134 235297
rect 328490 235257 328496 235269
rect 338128 235257 338134 235269
rect 338186 235257 338192 235309
rect 338512 235257 338518 235309
rect 338570 235297 338576 235309
rect 354832 235297 354838 235309
rect 338570 235269 354838 235297
rect 338570 235257 338576 235269
rect 354832 235257 354838 235269
rect 354890 235257 354896 235309
rect 355696 235257 355702 235309
rect 355754 235297 355760 235309
rect 372610 235297 372638 235343
rect 379504 235331 379510 235343
rect 379562 235331 379568 235383
rect 379984 235331 379990 235383
rect 380042 235371 380048 235383
rect 494704 235371 494710 235383
rect 380042 235343 494710 235371
rect 380042 235331 380048 235343
rect 494704 235331 494710 235343
rect 494762 235331 494768 235383
rect 379888 235297 379894 235309
rect 355754 235269 372638 235297
rect 372706 235269 379894 235297
rect 355754 235257 355760 235269
rect 317008 235183 317014 235235
rect 317066 235223 317072 235235
rect 317066 235195 344606 235223
rect 317066 235183 317072 235195
rect 140176 235109 140182 235161
rect 140234 235149 140240 235161
rect 141904 235149 141910 235161
rect 140234 235121 141910 235149
rect 140234 235109 140240 235121
rect 141904 235109 141910 235121
rect 141962 235109 141968 235161
rect 314032 235109 314038 235161
rect 314090 235149 314096 235161
rect 338320 235149 338326 235161
rect 314090 235121 338326 235149
rect 314090 235109 314096 235121
rect 338320 235109 338326 235121
rect 338378 235109 338384 235161
rect 338416 235109 338422 235161
rect 338474 235149 338480 235161
rect 344464 235149 344470 235161
rect 338474 235121 344470 235149
rect 338474 235109 338480 235121
rect 344464 235109 344470 235121
rect 344522 235109 344528 235161
rect 344578 235149 344606 235195
rect 354928 235183 354934 235235
rect 354986 235223 354992 235235
rect 372706 235223 372734 235269
rect 379888 235257 379894 235269
rect 379946 235257 379952 235309
rect 382192 235257 382198 235309
rect 382250 235297 382256 235309
rect 496912 235297 496918 235309
rect 382250 235269 496918 235297
rect 382250 235257 382256 235269
rect 496912 235257 496918 235269
rect 496970 235257 496976 235309
rect 376816 235223 376822 235235
rect 354986 235195 372734 235223
rect 372802 235195 376822 235223
rect 354986 235183 354992 235195
rect 360688 235149 360694 235161
rect 344578 235121 360694 235149
rect 360688 235109 360694 235121
rect 360746 235109 360752 235161
rect 360784 235109 360790 235161
rect 360842 235149 360848 235161
rect 372802 235149 372830 235195
rect 376816 235183 376822 235195
rect 376874 235183 376880 235235
rect 379216 235183 379222 235235
rect 379274 235223 379280 235235
rect 494032 235223 494038 235235
rect 379274 235195 494038 235223
rect 379274 235183 379280 235195
rect 494032 235183 494038 235195
rect 494090 235183 494096 235235
rect 360842 235121 372830 235149
rect 360842 235109 360848 235121
rect 376240 235109 376246 235161
rect 376298 235149 376304 235161
rect 491056 235149 491062 235161
rect 376298 235121 491062 235149
rect 376298 235109 376304 235121
rect 491056 235109 491062 235121
rect 491114 235109 491120 235161
rect 311152 235035 311158 235087
rect 311210 235075 311216 235087
rect 355024 235075 355030 235087
rect 311210 235047 355030 235075
rect 311210 235035 311216 235047
rect 355024 235035 355030 235047
rect 355082 235035 355088 235087
rect 357904 235035 357910 235087
rect 357962 235075 357968 235087
rect 372784 235075 372790 235087
rect 357962 235047 372790 235075
rect 357962 235035 357968 235047
rect 372784 235035 372790 235047
rect 372842 235035 372848 235087
rect 372976 235035 372982 235087
rect 373034 235075 373040 235087
rect 488848 235075 488854 235087
rect 373034 235047 488854 235075
rect 373034 235035 373040 235047
rect 488848 235035 488854 235047
rect 488906 235035 488912 235087
rect 318832 234961 318838 235013
rect 318890 235001 318896 235013
rect 356848 235001 356854 235013
rect 318890 234973 356854 235001
rect 318890 234961 318896 234973
rect 356848 234961 356854 234973
rect 356906 234961 356912 235013
rect 357136 234961 357142 235013
rect 357194 235001 357200 235013
rect 375376 235001 375382 235013
rect 357194 234973 375382 235001
rect 357194 234961 357200 234973
rect 375376 234961 375382 234973
rect 375434 234961 375440 235013
rect 377680 235001 377686 235013
rect 375490 234973 377686 235001
rect 321040 234887 321046 234939
rect 321098 234927 321104 234939
rect 357712 234927 357718 234939
rect 321098 234899 357718 234927
rect 321098 234887 321104 234899
rect 357712 234887 357718 234899
rect 357770 234887 357776 234939
rect 359344 234887 359350 234939
rect 359402 234927 359408 234939
rect 375490 234927 375518 234973
rect 377680 234961 377686 234973
rect 377738 234961 377744 235013
rect 378448 234961 378454 235013
rect 378506 235001 378512 235013
rect 493264 235001 493270 235013
rect 378506 234973 493270 235001
rect 378506 234961 378512 234973
rect 493264 234961 493270 234973
rect 493322 234961 493328 235013
rect 359402 234899 375518 234927
rect 359402 234887 359408 234899
rect 375568 234887 375574 234939
rect 375626 234927 375632 234939
rect 375626 234899 381374 234927
rect 375626 234887 375632 234899
rect 310000 234813 310006 234865
rect 310058 234853 310064 234865
rect 338224 234853 338230 234865
rect 310058 234825 338230 234853
rect 310058 234813 310064 234825
rect 338224 234813 338230 234825
rect 338282 234813 338288 234865
rect 338320 234813 338326 234865
rect 338378 234853 338384 234865
rect 359824 234853 359830 234865
rect 338378 234825 359830 234853
rect 338378 234813 338384 234825
rect 359824 234813 359830 234825
rect 359882 234813 359888 234865
rect 361168 234813 361174 234865
rect 361226 234853 361232 234865
rect 378736 234853 378742 234865
rect 361226 234825 378742 234853
rect 361226 234813 361232 234825
rect 378736 234813 378742 234825
rect 378794 234813 378800 234865
rect 381346 234853 381374 234899
rect 381424 234887 381430 234939
rect 381482 234927 381488 234939
rect 496144 234927 496150 234939
rect 381482 234899 496150 234927
rect 381482 234887 381488 234899
rect 496144 234887 496150 234899
rect 496202 234887 496208 234939
rect 490288 234853 490294 234865
rect 381346 234825 490294 234853
rect 490288 234813 490294 234825
rect 490346 234813 490352 234865
rect 318160 234739 318166 234791
rect 318218 234779 318224 234791
rect 356080 234779 356086 234791
rect 318218 234751 356086 234779
rect 318218 234739 318224 234751
rect 356080 234739 356086 234751
rect 356138 234739 356144 234791
rect 358576 234739 358582 234791
rect 358634 234779 358640 234791
rect 378064 234779 378070 234791
rect 358634 234751 378070 234779
rect 358634 234739 358640 234751
rect 378064 234739 378070 234751
rect 378122 234739 378128 234791
rect 380656 234739 380662 234791
rect 380714 234779 380720 234791
rect 495472 234779 495478 234791
rect 380714 234751 495478 234779
rect 380714 234739 380720 234751
rect 495472 234739 495478 234751
rect 495530 234739 495536 234791
rect 42352 234665 42358 234717
rect 42410 234705 42416 234717
rect 43504 234705 43510 234717
rect 42410 234677 43510 234705
rect 42410 234665 42416 234677
rect 43504 234665 43510 234677
rect 43562 234665 43568 234717
rect 317392 234665 317398 234717
rect 317450 234705 317456 234717
rect 355888 234705 355894 234717
rect 317450 234677 355894 234705
rect 317450 234665 317456 234677
rect 355888 234665 355894 234677
rect 355946 234665 355952 234717
rect 377776 234665 377782 234717
rect 377834 234705 377840 234717
rect 492496 234705 492502 234717
rect 377834 234677 492502 234705
rect 377834 234665 377840 234677
rect 492496 234665 492502 234677
rect 492554 234665 492560 234717
rect 328258 234603 328382 234631
rect 311824 234443 311830 234495
rect 311882 234483 311888 234495
rect 328258 234483 328286 234603
rect 328354 234557 328382 234603
rect 329872 234591 329878 234643
rect 329930 234631 329936 234643
rect 329930 234603 344414 234631
rect 329930 234591 329936 234603
rect 344272 234557 344278 234569
rect 328354 234529 344278 234557
rect 344272 234517 344278 234529
rect 344330 234517 344336 234569
rect 344386 234557 344414 234603
rect 344464 234591 344470 234643
rect 344522 234631 344528 234643
rect 378640 234631 378646 234643
rect 344522 234603 378646 234631
rect 344522 234591 344528 234603
rect 378640 234591 378646 234603
rect 378698 234591 378704 234643
rect 378832 234591 378838 234643
rect 378890 234631 378896 234643
rect 390544 234631 390550 234643
rect 378890 234603 390550 234631
rect 378890 234591 378896 234603
rect 390544 234591 390550 234603
rect 390602 234591 390608 234643
rect 395728 234591 395734 234643
rect 395786 234631 395792 234643
rect 408688 234631 408694 234643
rect 395786 234603 408694 234631
rect 395786 234591 395792 234603
rect 408688 234591 408694 234603
rect 408746 234591 408752 234643
rect 414736 234591 414742 234643
rect 414794 234631 414800 234643
rect 415984 234631 415990 234643
rect 414794 234603 415990 234631
rect 414794 234591 414800 234603
rect 415984 234591 415990 234603
rect 416042 234591 416048 234643
rect 417712 234591 417718 234643
rect 417770 234631 417776 234643
rect 419920 234631 419926 234643
rect 417770 234603 419926 234631
rect 417770 234591 417776 234603
rect 419920 234591 419926 234603
rect 419978 234591 419984 234643
rect 420016 234591 420022 234643
rect 420074 234631 420080 234643
rect 443536 234631 443542 234643
rect 420074 234603 443542 234631
rect 420074 234591 420080 234603
rect 443536 234591 443542 234603
rect 443594 234591 443600 234643
rect 443632 234591 443638 234643
rect 443690 234631 443696 234643
rect 446416 234631 446422 234643
rect 443690 234603 446422 234631
rect 443690 234591 443696 234603
rect 446416 234591 446422 234603
rect 446474 234591 446480 234643
rect 448432 234591 448438 234643
rect 448490 234631 448496 234643
rect 498064 234631 498070 234643
rect 448490 234603 498070 234631
rect 448490 234591 448496 234603
rect 498064 234591 498070 234603
rect 498122 234591 498128 234643
rect 375952 234557 375958 234569
rect 344386 234529 375958 234557
rect 375952 234517 375958 234529
rect 376010 234517 376016 234569
rect 396496 234517 396502 234569
rect 396554 234557 396560 234569
rect 405040 234557 405046 234569
rect 396554 234529 405046 234557
rect 396554 234517 396560 234529
rect 405040 234517 405046 234529
rect 405098 234517 405104 234569
rect 408304 234517 408310 234569
rect 408362 234557 408368 234569
rect 439120 234557 439126 234569
rect 408362 234529 439126 234557
rect 408362 234517 408368 234529
rect 439120 234517 439126 234529
rect 439178 234517 439184 234569
rect 442480 234517 442486 234569
rect 442538 234557 442544 234569
rect 447472 234557 447478 234569
rect 442538 234529 447478 234557
rect 442538 234517 442544 234529
rect 447472 234517 447478 234529
rect 447530 234517 447536 234569
rect 451312 234517 451318 234569
rect 451370 234557 451376 234569
rect 499696 234557 499702 234569
rect 451370 234529 499702 234557
rect 451370 234517 451376 234529
rect 499696 234517 499702 234529
rect 499754 234517 499760 234569
rect 311882 234455 328286 234483
rect 311882 234443 311888 234455
rect 329488 234443 329494 234495
rect 329546 234483 329552 234495
rect 338992 234483 338998 234495
rect 329546 234455 338998 234483
rect 329546 234443 329552 234455
rect 338992 234443 338998 234455
rect 339050 234443 339056 234495
rect 342736 234443 342742 234495
rect 342794 234483 342800 234495
rect 398128 234483 398134 234495
rect 342794 234455 398134 234483
rect 342794 234443 342800 234455
rect 398128 234443 398134 234455
rect 398186 234443 398192 234495
rect 399184 234443 399190 234495
rect 399242 234483 399248 234495
rect 408784 234483 408790 234495
rect 399242 234455 408790 234483
rect 399242 234443 399248 234455
rect 408784 234443 408790 234455
rect 408842 234443 408848 234495
rect 408976 234443 408982 234495
rect 409034 234483 409040 234495
rect 417424 234483 417430 234495
rect 409034 234455 417430 234483
rect 409034 234443 409040 234455
rect 417424 234443 417430 234455
rect 417482 234443 417488 234495
rect 417808 234443 417814 234495
rect 417866 234483 417872 234495
rect 425872 234483 425878 234495
rect 417866 234455 425878 234483
rect 417866 234443 417872 234455
rect 425872 234443 425878 234455
rect 425930 234443 425936 234495
rect 426160 234443 426166 234495
rect 426218 234483 426224 234495
rect 446128 234483 446134 234495
rect 426218 234455 446134 234483
rect 426218 234443 426224 234455
rect 446128 234443 446134 234455
rect 446186 234443 446192 234495
rect 446224 234443 446230 234495
rect 446282 234483 446288 234495
rect 493936 234483 493942 234495
rect 446282 234455 493942 234483
rect 446282 234443 446288 234455
rect 493936 234443 493942 234455
rect 493994 234443 494000 234495
rect 312208 234369 312214 234421
rect 312266 234409 312272 234421
rect 354736 234409 354742 234421
rect 312266 234381 354742 234409
rect 312266 234369 312272 234381
rect 354736 234369 354742 234381
rect 354794 234369 354800 234421
rect 360976 234409 360982 234421
rect 355810 234381 360982 234409
rect 310768 234295 310774 234347
rect 310826 234335 310832 234347
rect 351664 234335 351670 234347
rect 310826 234307 351670 234335
rect 310826 234295 310832 234307
rect 351664 234295 351670 234307
rect 351722 234295 351728 234347
rect 353488 234295 353494 234347
rect 353546 234335 353552 234347
rect 355810 234335 355838 234381
rect 360976 234369 360982 234381
rect 361034 234369 361040 234421
rect 361936 234369 361942 234421
rect 361994 234409 362000 234421
rect 393424 234409 393430 234421
rect 361994 234381 393430 234409
rect 361994 234369 362000 234381
rect 393424 234369 393430 234381
rect 393482 234369 393488 234421
rect 393520 234369 393526 234421
rect 393578 234409 393584 234421
rect 400240 234409 400246 234421
rect 393578 234381 400246 234409
rect 393578 234369 393584 234381
rect 400240 234369 400246 234381
rect 400298 234369 400304 234421
rect 400336 234369 400342 234421
rect 400394 234409 400400 234421
rect 408016 234409 408022 234421
rect 400394 234381 408022 234409
rect 400394 234369 400400 234381
rect 408016 234369 408022 234381
rect 408074 234369 408080 234421
rect 408112 234369 408118 234421
rect 408170 234409 408176 234421
rect 418864 234409 418870 234421
rect 408170 234381 418870 234409
rect 408170 234369 408176 234381
rect 418864 234369 418870 234381
rect 418922 234369 418928 234421
rect 424240 234409 424246 234421
rect 418978 234381 424246 234409
rect 353546 234307 355838 234335
rect 353546 234295 353552 234307
rect 355888 234295 355894 234347
rect 355946 234335 355952 234347
rect 363472 234335 363478 234347
rect 355946 234307 363478 234335
rect 355946 234295 355952 234307
rect 363472 234295 363478 234307
rect 363530 234295 363536 234347
rect 365968 234295 365974 234347
rect 366026 234335 366032 234347
rect 367984 234335 367990 234347
rect 366026 234307 367990 234335
rect 366026 234295 366032 234307
rect 367984 234295 367990 234307
rect 368042 234295 368048 234347
rect 368656 234295 368662 234347
rect 368714 234335 368720 234347
rect 376240 234335 376246 234347
rect 368714 234307 376246 234335
rect 368714 234295 368720 234307
rect 376240 234295 376246 234307
rect 376298 234295 376304 234347
rect 388048 234295 388054 234347
rect 388106 234335 388112 234347
rect 408400 234335 408406 234347
rect 388106 234307 408406 234335
rect 388106 234295 388112 234307
rect 408400 234295 408406 234307
rect 408458 234295 408464 234347
rect 418978 234335 419006 234381
rect 424240 234369 424246 234381
rect 424298 234369 424304 234421
rect 431920 234369 431926 234421
rect 431978 234409 431984 234421
rect 452176 234409 452182 234421
rect 431978 234381 452182 234409
rect 431978 234369 431984 234381
rect 452176 234369 452182 234381
rect 452234 234369 452240 234421
rect 452848 234369 452854 234421
rect 452906 234409 452912 234421
rect 499600 234409 499606 234421
rect 452906 234381 499606 234409
rect 452906 234369 452912 234381
rect 499600 234369 499606 234381
rect 499658 234369 499664 234421
rect 428080 234335 428086 234347
rect 408514 234307 419006 234335
rect 419074 234307 428086 234335
rect 320368 234221 320374 234273
rect 320426 234261 320432 234273
rect 359920 234261 359926 234273
rect 320426 234233 359926 234261
rect 320426 234221 320432 234233
rect 359920 234221 359926 234233
rect 359978 234221 359984 234273
rect 361552 234221 361558 234273
rect 361610 234261 361616 234273
rect 376528 234261 376534 234273
rect 361610 234233 376534 234261
rect 361610 234221 361616 234233
rect 376528 234221 376534 234233
rect 376586 234221 376592 234273
rect 377200 234221 377206 234273
rect 377258 234261 377264 234273
rect 397360 234261 397366 234273
rect 377258 234233 397366 234261
rect 377258 234221 377264 234233
rect 397360 234221 397366 234233
rect 397418 234221 397424 234273
rect 399280 234261 399286 234273
rect 397474 234233 399286 234261
rect 42448 234187 42454 234199
rect 42082 234159 42454 234187
rect 42082 234051 42110 234159
rect 42448 234147 42454 234159
rect 42506 234147 42512 234199
rect 323632 234147 323638 234199
rect 323690 234187 323696 234199
rect 338512 234187 338518 234199
rect 323690 234159 338518 234187
rect 323690 234147 323696 234159
rect 338512 234147 338518 234159
rect 338570 234147 338576 234199
rect 338608 234147 338614 234199
rect 338666 234187 338672 234199
rect 355120 234187 355126 234199
rect 338666 234159 355126 234187
rect 338666 234147 338672 234159
rect 355120 234147 355126 234159
rect 355178 234147 355184 234199
rect 362320 234147 362326 234199
rect 362378 234187 362384 234199
rect 368656 234187 368662 234199
rect 362378 234159 368662 234187
rect 362378 234147 362384 234159
rect 368656 234147 368662 234159
rect 368714 234147 368720 234199
rect 374992 234147 374998 234199
rect 375050 234187 375056 234199
rect 394576 234187 394582 234199
rect 375050 234159 394582 234187
rect 375050 234147 375056 234159
rect 394576 234147 394582 234159
rect 394634 234147 394640 234199
rect 397264 234147 397270 234199
rect 397322 234187 397328 234199
rect 397474 234187 397502 234233
rect 399280 234221 399286 234233
rect 399338 234221 399344 234273
rect 399472 234221 399478 234273
rect 399530 234261 399536 234273
rect 399530 234233 405758 234261
rect 399530 234221 399536 234233
rect 397322 234159 397502 234187
rect 397322 234147 397328 234159
rect 397552 234147 397558 234199
rect 397610 234187 397616 234199
rect 404656 234187 404662 234199
rect 397610 234159 404662 234187
rect 397610 234147 397616 234159
rect 404656 234147 404662 234159
rect 404714 234147 404720 234199
rect 313744 234073 313750 234125
rect 313802 234113 313808 234125
rect 327184 234113 327190 234125
rect 313802 234085 327190 234113
rect 313802 234073 313808 234085
rect 327184 234073 327190 234085
rect 327242 234073 327248 234125
rect 328720 234073 328726 234125
rect 328778 234113 328784 234125
rect 346672 234113 346678 234125
rect 328778 234085 346678 234113
rect 328778 234073 328784 234085
rect 346672 234073 346678 234085
rect 346730 234073 346736 234125
rect 346768 234073 346774 234125
rect 346826 234113 346832 234125
rect 352624 234113 352630 234125
rect 346826 234085 352630 234113
rect 346826 234073 346832 234085
rect 352624 234073 352630 234085
rect 352682 234073 352688 234125
rect 352720 234073 352726 234125
rect 352778 234113 352784 234125
rect 362800 234113 362806 234125
rect 352778 234085 362806 234113
rect 352778 234073 352784 234085
rect 362800 234073 362806 234085
rect 362858 234073 362864 234125
rect 375952 234073 375958 234125
rect 376010 234113 376016 234125
rect 395152 234113 395158 234125
rect 376010 234085 395158 234113
rect 376010 234073 376016 234085
rect 395152 234073 395158 234085
rect 395210 234073 395216 234125
rect 396880 234073 396886 234125
rect 396938 234113 396944 234125
rect 405136 234113 405142 234125
rect 396938 234085 405142 234113
rect 396938 234073 396944 234085
rect 405136 234073 405142 234085
rect 405194 234073 405200 234125
rect 405730 234113 405758 234233
rect 407056 234221 407062 234273
rect 407114 234261 407120 234273
rect 408514 234261 408542 234307
rect 407114 234233 408542 234261
rect 407114 234221 407120 234233
rect 410032 234221 410038 234273
rect 410090 234261 410096 234273
rect 416752 234261 416758 234273
rect 410090 234233 416758 234261
rect 410090 234221 410096 234233
rect 416752 234221 416758 234233
rect 416810 234221 416816 234273
rect 418480 234221 418486 234273
rect 418538 234261 418544 234273
rect 419074 234261 419102 234307
rect 428080 234295 428086 234307
rect 428138 234295 428144 234347
rect 431440 234295 431446 234347
rect 431498 234335 431504 234347
rect 475600 234335 475606 234347
rect 431498 234307 475606 234335
rect 431498 234295 431504 234307
rect 475600 234295 475606 234307
rect 475658 234295 475664 234347
rect 418538 234233 419102 234261
rect 418538 234221 418544 234233
rect 422992 234221 422998 234273
rect 423050 234261 423056 234273
rect 450544 234261 450550 234273
rect 423050 234233 450550 234261
rect 423050 234221 423056 234233
rect 450544 234221 450550 234233
rect 450602 234221 450608 234273
rect 450640 234221 450646 234273
rect 450698 234261 450704 234273
rect 451888 234261 451894 234273
rect 450698 234233 451894 234261
rect 450698 234221 450704 234233
rect 451888 234221 451894 234233
rect 451946 234221 451952 234273
rect 405904 234147 405910 234199
rect 405962 234187 405968 234199
rect 415312 234187 415318 234199
rect 405962 234159 415318 234187
rect 405962 234147 405968 234159
rect 415312 234147 415318 234159
rect 415370 234147 415376 234199
rect 415504 234147 415510 234199
rect 415562 234187 415568 234199
rect 425392 234187 425398 234199
rect 415562 234159 425398 234187
rect 415562 234147 415568 234159
rect 425392 234147 425398 234159
rect 425450 234147 425456 234199
rect 425968 234147 425974 234199
rect 426026 234187 426032 234199
rect 470032 234187 470038 234199
rect 426026 234159 470038 234187
rect 426026 234147 426032 234159
rect 470032 234147 470038 234159
rect 470090 234147 470096 234199
rect 405730 234085 408734 234113
rect 42064 233999 42070 234051
rect 42122 233999 42128 234051
rect 42448 233999 42454 234051
rect 42506 234039 42512 234051
rect 43120 234039 43126 234051
rect 42506 234011 43126 234039
rect 42506 233999 42512 234011
rect 43120 233999 43126 234011
rect 43178 233999 43184 234051
rect 314416 233999 314422 234051
rect 314474 234039 314480 234051
rect 327088 234039 327094 234051
rect 314474 234011 327094 234039
rect 314474 233999 314480 234011
rect 327088 233999 327094 234011
rect 327146 233999 327152 234051
rect 338320 233999 338326 234051
rect 338378 234039 338384 234051
rect 351472 234039 351478 234051
rect 338378 234011 351478 234039
rect 338378 233999 338384 234011
rect 351472 233999 351478 234011
rect 351530 233999 351536 234051
rect 352336 233999 352342 234051
rect 352394 234039 352400 234051
rect 398896 234039 398902 234051
rect 352394 234011 398902 234039
rect 352394 233999 352400 234011
rect 398896 233999 398902 234011
rect 398954 233999 398960 234051
rect 400144 233999 400150 234051
rect 400202 234039 400208 234051
rect 408592 234039 408598 234051
rect 400202 234011 408598 234039
rect 400202 233999 400208 234011
rect 408592 233999 408598 234011
rect 408650 233999 408656 234051
rect 408706 234039 408734 234085
rect 408880 234073 408886 234125
rect 408938 234113 408944 234125
rect 410800 234113 410806 234125
rect 408938 234085 410806 234113
rect 408938 234073 408944 234085
rect 410800 234073 410806 234085
rect 410858 234073 410864 234125
rect 410896 234073 410902 234125
rect 410954 234113 410960 234125
rect 426256 234113 426262 234125
rect 410954 234085 426262 234113
rect 410954 234073 410960 234085
rect 426256 234073 426262 234085
rect 426314 234073 426320 234125
rect 427408 234073 427414 234125
rect 427466 234113 427472 234125
rect 471568 234113 471574 234125
rect 427466 234085 471574 234113
rect 427466 234073 427472 234085
rect 471568 234073 471574 234085
rect 471626 234073 471632 234125
rect 410128 234039 410134 234051
rect 408706 234011 410134 234039
rect 410128 233999 410134 234011
rect 410186 233999 410192 234051
rect 410416 233999 410422 234051
rect 410474 234039 410480 234051
rect 415216 234039 415222 234051
rect 410474 234011 415222 234039
rect 410474 233999 410480 234011
rect 415216 233999 415222 234011
rect 415274 233999 415280 234051
rect 416368 233999 416374 234051
rect 416426 234039 416432 234051
rect 428464 234039 428470 234051
rect 416426 234011 428470 234039
rect 416426 233999 416432 234011
rect 428464 233999 428470 234011
rect 428522 233999 428528 234051
rect 428848 233999 428854 234051
rect 428906 234039 428912 234051
rect 470608 234039 470614 234051
rect 428906 234011 470614 234039
rect 428906 233999 428912 234011
rect 470608 233999 470614 234011
rect 470666 233999 470672 234051
rect 322192 233925 322198 233977
rect 322250 233965 322256 233977
rect 338416 233965 338422 233977
rect 322250 233937 338422 233965
rect 322250 233925 322256 233937
rect 338416 233925 338422 233937
rect 338474 233925 338480 233977
rect 338704 233925 338710 233977
rect 338762 233965 338768 233977
rect 349168 233965 349174 233977
rect 338762 233937 349174 233965
rect 338762 233925 338768 233937
rect 349168 233925 349174 233937
rect 349226 233925 349232 233977
rect 356080 233925 356086 233977
rect 356138 233965 356144 233977
rect 363568 233965 363574 233977
rect 356138 233937 363574 233965
rect 356138 233925 356144 233937
rect 363568 233925 363574 233937
rect 363626 233925 363632 233977
rect 375088 233965 375094 233977
rect 368770 233937 375094 233965
rect 319600 233851 319606 233903
rect 319658 233891 319664 233903
rect 354448 233891 354454 233903
rect 319658 233863 354454 233891
rect 319658 233851 319664 233863
rect 354448 233851 354454 233863
rect 354506 233851 354512 233903
rect 364528 233851 364534 233903
rect 364586 233891 364592 233903
rect 368770 233891 368798 233937
rect 375088 233925 375094 233937
rect 375146 233925 375152 233977
rect 378640 233925 378646 233977
rect 378698 233965 378704 233977
rect 395248 233965 395254 233977
rect 378698 233937 395254 233965
rect 378698 233925 378704 233937
rect 395248 233925 395254 233937
rect 395306 233925 395312 233977
rect 400624 233925 400630 233977
rect 400682 233965 400688 233977
rect 407920 233965 407926 233977
rect 400682 233937 407926 233965
rect 400682 233925 400688 233937
rect 407920 233925 407926 233937
rect 407978 233925 407984 233977
rect 411760 233925 411766 233977
rect 411818 233965 411824 233977
rect 429904 233965 429910 233977
rect 411818 233937 429910 233965
rect 411818 233925 411824 233937
rect 429904 233925 429910 233937
rect 429962 233925 429968 233977
rect 430768 233925 430774 233977
rect 430826 233965 430832 233977
rect 474832 233965 474838 233977
rect 430826 233937 474838 233965
rect 430826 233925 430832 233937
rect 474832 233925 474838 233937
rect 474890 233925 474896 233977
rect 364586 233863 368798 233891
rect 364586 233851 364592 233863
rect 374320 233851 374326 233903
rect 374378 233891 374384 233903
rect 388336 233891 388342 233903
rect 374378 233863 388342 233891
rect 374378 233851 374384 233863
rect 388336 233851 388342 233863
rect 388394 233851 388400 233903
rect 394768 233851 394774 233903
rect 394826 233891 394832 233903
rect 400528 233891 400534 233903
rect 394826 233863 400534 233891
rect 394826 233851 394832 233863
rect 400528 233851 400534 233863
rect 400586 233851 400592 233903
rect 400912 233851 400918 233903
rect 400970 233891 400976 233903
rect 407152 233891 407158 233903
rect 400970 233863 407158 233891
rect 400970 233851 400976 233863
rect 407152 233851 407158 233863
rect 407210 233851 407216 233903
rect 407248 233851 407254 233903
rect 407306 233891 407312 233903
rect 410032 233891 410038 233903
rect 407306 233863 410038 233891
rect 407306 233851 407312 233863
rect 410032 233851 410038 233863
rect 410090 233851 410096 233903
rect 413776 233891 413782 233903
rect 410146 233863 413782 233891
rect 319984 233777 319990 233829
rect 320042 233817 320048 233829
rect 354256 233817 354262 233829
rect 320042 233789 354262 233817
rect 320042 233777 320048 233789
rect 354256 233777 354262 233789
rect 354314 233777 354320 233829
rect 357712 233777 357718 233829
rect 357770 233817 357776 233829
rect 357770 233789 359774 233817
rect 357770 233777 357776 233789
rect 320656 233703 320662 233755
rect 320714 233743 320720 233755
rect 320714 233715 327038 233743
rect 320714 233703 320720 233715
rect 308944 233629 308950 233681
rect 309002 233669 309008 233681
rect 326896 233669 326902 233681
rect 309002 233641 326902 233669
rect 309002 233629 309008 233641
rect 326896 233629 326902 233641
rect 326954 233629 326960 233681
rect 321424 233555 321430 233607
rect 321482 233595 321488 233607
rect 327010 233595 327038 233715
rect 327088 233703 327094 233755
rect 327146 233743 327152 233755
rect 327146 233715 338366 233743
rect 327146 233703 327152 233715
rect 327184 233629 327190 233681
rect 327242 233669 327248 233681
rect 328720 233669 328726 233681
rect 327242 233641 328726 233669
rect 327242 233629 327248 233641
rect 328720 233629 328726 233641
rect 328778 233629 328784 233681
rect 328816 233629 328822 233681
rect 328874 233669 328880 233681
rect 330448 233669 330454 233681
rect 328874 233641 330454 233669
rect 328874 233629 328880 233641
rect 330448 233629 330454 233641
rect 330506 233629 330512 233681
rect 338338 233669 338366 233715
rect 338416 233703 338422 233755
rect 338474 233743 338480 233755
rect 359536 233743 359542 233755
rect 338474 233715 359542 233743
rect 338474 233703 338480 233715
rect 359536 233703 359542 233715
rect 359594 233703 359600 233755
rect 359746 233743 359774 233789
rect 360976 233777 360982 233829
rect 361034 233817 361040 233829
rect 365104 233817 365110 233829
rect 361034 233789 365110 233817
rect 361034 233777 361040 233789
rect 365104 233777 365110 233789
rect 365162 233777 365168 233829
rect 365200 233777 365206 233829
rect 365258 233817 365264 233829
rect 368656 233817 368662 233829
rect 365258 233789 368662 233817
rect 365258 233777 365264 233789
rect 368656 233777 368662 233789
rect 368714 233777 368720 233829
rect 387664 233817 387670 233829
rect 373282 233789 387670 233817
rect 366640 233743 366646 233755
rect 359746 233715 366646 233743
rect 366640 233703 366646 233715
rect 366698 233703 366704 233755
rect 373282 233743 373310 233789
rect 387664 233777 387670 233789
rect 387722 233777 387728 233829
rect 393424 233777 393430 233829
rect 393482 233817 393488 233829
rect 398896 233817 398902 233829
rect 393482 233789 398902 233817
rect 393482 233777 393488 233789
rect 398896 233777 398902 233789
rect 398954 233777 398960 233829
rect 399856 233777 399862 233829
rect 399914 233817 399920 233829
rect 404560 233817 404566 233829
rect 399914 233789 404566 233817
rect 399914 233777 399920 233789
rect 404560 233777 404566 233789
rect 404618 233777 404624 233829
rect 404656 233777 404662 233829
rect 404714 233817 404720 233829
rect 410146 233817 410174 233863
rect 413776 233851 413782 233863
rect 413834 233851 413840 233903
rect 413872 233851 413878 233903
rect 413930 233891 413936 233903
rect 425104 233891 425110 233903
rect 413930 233863 425110 233891
rect 413930 233851 413936 233863
rect 425104 233851 425110 233863
rect 425162 233851 425168 233903
rect 425200 233851 425206 233903
rect 425258 233891 425264 233903
rect 469360 233891 469366 233903
rect 425258 233863 469366 233891
rect 425258 233851 425264 233863
rect 469360 233851 469366 233863
rect 469418 233851 469424 233903
rect 404714 233789 410174 233817
rect 404714 233777 404720 233789
rect 410512 233777 410518 233829
rect 410570 233817 410576 233829
rect 428368 233817 428374 233829
rect 410570 233789 428374 233817
rect 410570 233777 410576 233789
rect 428368 233777 428374 233789
rect 428426 233777 428432 233829
rect 428464 233777 428470 233829
rect 428522 233817 428528 233829
rect 456112 233817 456118 233829
rect 428522 233789 456118 233817
rect 428522 233777 428528 233789
rect 456112 233777 456118 233789
rect 456170 233777 456176 233829
rect 372994 233715 373310 233743
rect 348496 233669 348502 233681
rect 338338 233641 348502 233669
rect 348496 233629 348502 233641
rect 348554 233629 348560 233681
rect 352624 233629 352630 233681
rect 352682 233669 352688 233681
rect 367120 233669 367126 233681
rect 352682 233641 367126 233669
rect 352682 233629 352688 233641
rect 367120 233629 367126 233641
rect 367178 233629 367184 233681
rect 371152 233629 371158 233681
rect 371210 233669 371216 233681
rect 371920 233669 371926 233681
rect 371210 233641 371926 233669
rect 371210 233629 371216 233641
rect 371920 233629 371926 233641
rect 371978 233629 371984 233681
rect 372304 233629 372310 233681
rect 372362 233669 372368 233681
rect 372994 233669 373022 233715
rect 376912 233703 376918 233755
rect 376970 233743 376976 233755
rect 386896 233743 386902 233755
rect 376970 233715 386902 233743
rect 376970 233703 376976 233715
rect 386896 233703 386902 233715
rect 386954 233703 386960 233755
rect 396112 233703 396118 233755
rect 396170 233743 396176 233755
rect 401872 233743 401878 233755
rect 396170 233715 401878 233743
rect 396170 233703 396176 233715
rect 401872 233703 401878 233715
rect 401930 233703 401936 233755
rect 401968 233703 401974 233755
rect 402026 233743 402032 233755
rect 404944 233743 404950 233755
rect 402026 233715 404950 233743
rect 402026 233703 402032 233715
rect 404944 233703 404950 233715
rect 405002 233703 405008 233755
rect 405040 233703 405046 233755
rect 405098 233743 405104 233755
rect 414736 233743 414742 233755
rect 405098 233715 414742 233743
rect 405098 233703 405104 233715
rect 414736 233703 414742 233715
rect 414794 233703 414800 233755
rect 429424 233743 429430 233755
rect 418978 233715 429430 233743
rect 372362 233641 373022 233669
rect 372362 233629 372368 233641
rect 392464 233629 392470 233681
rect 392522 233669 392528 233681
rect 401200 233669 401206 233681
rect 392522 233641 401206 233669
rect 392522 233629 392528 233641
rect 401200 233629 401206 233641
rect 401258 233629 401264 233681
rect 401296 233629 401302 233681
rect 401354 233669 401360 233681
rect 404080 233669 404086 233681
rect 401354 233641 404086 233669
rect 401354 233629 401360 233641
rect 404080 233629 404086 233641
rect 404138 233629 404144 233681
rect 405232 233629 405238 233681
rect 405290 233669 405296 233681
rect 415504 233669 415510 233681
rect 405290 233641 415510 233669
rect 405290 233629 405296 233641
rect 415504 233629 415510 233641
rect 415562 233629 415568 233681
rect 415600 233629 415606 233681
rect 415658 233669 415664 233681
rect 417520 233669 417526 233681
rect 415658 233641 417526 233669
rect 415658 233629 415664 233641
rect 417520 233629 417526 233641
rect 417578 233629 417584 233681
rect 351376 233595 351382 233607
rect 321482 233567 326942 233595
rect 327010 233567 351382 233595
rect 321482 233555 321488 233567
rect 308560 233481 308566 233533
rect 308618 233521 308624 233533
rect 326800 233521 326806 233533
rect 308618 233493 326806 233521
rect 308618 233481 308624 233493
rect 326800 233481 326806 233493
rect 326858 233481 326864 233533
rect 326914 233521 326942 233567
rect 351376 233555 351382 233567
rect 351434 233555 351440 233607
rect 353104 233555 353110 233607
rect 353162 233595 353168 233607
rect 398704 233595 398710 233607
rect 353162 233567 398710 233595
rect 353162 233555 353168 233567
rect 398704 233555 398710 233567
rect 398762 233555 398768 233607
rect 401680 233555 401686 233607
rect 401738 233595 401744 233607
rect 405712 233595 405718 233607
rect 401738 233567 405718 233595
rect 401738 233555 401744 233567
rect 405712 233555 405718 233567
rect 405770 233555 405776 233607
rect 411760 233555 411766 233607
rect 411818 233595 411824 233607
rect 418978 233595 419006 233715
rect 429424 233703 429430 233715
rect 429482 233703 429488 233755
rect 437392 233703 437398 233755
rect 437450 233743 437456 233755
rect 475120 233743 475126 233755
rect 437450 233715 475126 233743
rect 437450 233703 437456 233715
rect 475120 233703 475126 233715
rect 475178 233703 475184 233755
rect 419920 233629 419926 233681
rect 419978 233669 419984 233681
rect 426160 233669 426166 233681
rect 419978 233641 426166 233669
rect 419978 233629 419984 233641
rect 426160 233629 426166 233641
rect 426218 233629 426224 233681
rect 426256 233629 426262 233681
rect 426314 233669 426320 233681
rect 428272 233669 428278 233681
rect 426314 233641 428278 233669
rect 426314 233629 426320 233641
rect 428272 233629 428278 233641
rect 428330 233629 428336 233681
rect 436624 233629 436630 233681
rect 436682 233669 436688 233681
rect 466576 233669 466582 233681
rect 436682 233641 466582 233669
rect 436682 233629 436688 233641
rect 466576 233629 466582 233641
rect 466634 233629 466640 233681
rect 411818 233567 419006 233595
rect 411818 233555 411824 233567
rect 427792 233555 427798 233607
rect 427850 233595 427856 233607
rect 428464 233595 428470 233607
rect 427850 233567 428470 233595
rect 427850 233555 427856 233567
rect 428464 233555 428470 233567
rect 428522 233555 428528 233607
rect 435184 233555 435190 233607
rect 435242 233595 435248 233607
rect 437680 233595 437686 233607
rect 435242 233567 437686 233595
rect 435242 233555 435248 233567
rect 437680 233555 437686 233567
rect 437738 233555 437744 233607
rect 438064 233555 438070 233607
rect 438122 233595 438128 233607
rect 440560 233595 440566 233607
rect 438122 233567 440566 233595
rect 438122 233555 438128 233567
rect 440560 233555 440566 233567
rect 440618 233555 440624 233607
rect 443536 233555 443542 233607
rect 443594 233595 443600 233607
rect 446320 233595 446326 233607
rect 443594 233567 446326 233595
rect 443594 233555 443600 233567
rect 446320 233555 446326 233567
rect 446378 233555 446384 233607
rect 446512 233555 446518 233607
rect 446570 233595 446576 233607
rect 446896 233595 446902 233607
rect 446570 233567 446902 233595
rect 446570 233555 446576 233567
rect 446896 233555 446902 233567
rect 446954 233555 446960 233607
rect 450544 233555 450550 233607
rect 450602 233595 450608 233607
rect 467152 233595 467158 233607
rect 450602 233567 467158 233595
rect 450602 233555 450608 233567
rect 467152 233555 467158 233567
rect 467210 233555 467216 233607
rect 338320 233521 338326 233533
rect 326914 233493 338326 233521
rect 338320 233481 338326 233493
rect 338378 233481 338384 233533
rect 338512 233481 338518 233533
rect 338570 233521 338576 233533
rect 362704 233521 362710 233533
rect 338570 233493 362710 233521
rect 338570 233481 338576 233493
rect 362704 233481 362710 233493
rect 362762 233481 362768 233533
rect 362800 233481 362806 233533
rect 362858 233521 362864 233533
rect 367600 233521 367606 233533
rect 362858 233493 367606 233521
rect 362858 233481 362864 233493
rect 367600 233481 367606 233493
rect 367658 233481 367664 233533
rect 368656 233481 368662 233533
rect 368714 233521 368720 233533
rect 374704 233521 374710 233533
rect 368714 233493 374710 233521
rect 368714 233481 368720 233493
rect 374704 233481 374710 233493
rect 374762 233481 374768 233533
rect 378736 233481 378742 233533
rect 378794 233521 378800 233533
rect 398416 233521 398422 233533
rect 378794 233493 398422 233521
rect 378794 233481 378800 233493
rect 398416 233481 398422 233493
rect 398474 233481 398480 233533
rect 402064 233481 402070 233533
rect 402122 233521 402128 233533
rect 402928 233521 402934 233533
rect 402122 233493 402934 233521
rect 402122 233481 402128 233493
rect 402928 233481 402934 233493
rect 402986 233481 402992 233533
rect 410416 233521 410422 233533
rect 403234 233493 410422 233521
rect 322864 233407 322870 233459
rect 322922 233447 322928 233459
rect 348592 233447 348598 233459
rect 322922 233419 348598 233447
rect 322922 233407 322928 233419
rect 348592 233407 348598 233419
rect 348650 233407 348656 233459
rect 356848 233407 356854 233459
rect 356906 233447 356912 233459
rect 365104 233447 365110 233459
rect 356906 233419 365110 233447
rect 356906 233407 356912 233419
rect 365104 233407 365110 233419
rect 365162 233407 365168 233459
rect 365200 233407 365206 233459
rect 365258 233447 365264 233459
rect 366448 233447 366454 233459
rect 365258 233419 366454 233447
rect 365258 233407 365264 233419
rect 366448 233407 366454 233419
rect 366506 233407 366512 233459
rect 376912 233447 376918 233459
rect 372418 233419 376918 233447
rect 144016 233333 144022 233385
rect 144074 233373 144080 233385
rect 149200 233373 149206 233385
rect 144074 233345 149206 233373
rect 144074 233333 144080 233345
rect 149200 233333 149206 233345
rect 149258 233333 149264 233385
rect 286192 233333 286198 233385
rect 286250 233373 286256 233385
rect 368560 233373 368566 233385
rect 286250 233345 368566 233373
rect 286250 233333 286256 233345
rect 368560 233333 368566 233345
rect 368618 233333 368624 233385
rect 368656 233333 368662 233385
rect 368714 233373 368720 233385
rect 372418 233373 372446 233419
rect 376912 233407 376918 233419
rect 376970 233407 376976 233459
rect 377104 233407 377110 233459
rect 377162 233447 377168 233459
rect 397744 233447 397750 233459
rect 377162 233419 397750 233447
rect 377162 233407 377168 233419
rect 397744 233407 397750 233419
rect 397802 233407 397808 233459
rect 368714 233345 372446 233373
rect 368714 233333 368720 233345
rect 397072 233333 397078 233385
rect 397130 233373 397136 233385
rect 403234 233373 403262 233493
rect 410416 233481 410422 233493
rect 410474 233481 410480 233533
rect 413776 233481 413782 233533
rect 413834 233521 413840 233533
rect 432496 233521 432502 233533
rect 413834 233493 432502 233521
rect 413834 233481 413840 233493
rect 432496 233481 432502 233493
rect 432554 233481 432560 233533
rect 436240 233481 436246 233533
rect 436298 233521 436304 233533
rect 453616 233521 453622 233533
rect 436298 233493 453622 233521
rect 436298 233481 436304 233493
rect 453616 233481 453622 233493
rect 453674 233481 453680 233533
rect 403504 233407 403510 233459
rect 403562 233447 403568 233459
rect 481840 233447 481846 233459
rect 403562 233419 481846 233447
rect 403562 233407 403568 233419
rect 481840 233407 481846 233419
rect 481898 233407 481904 233459
rect 397130 233345 403262 233373
rect 397130 233333 397136 233345
rect 404464 233333 404470 233385
rect 404522 233373 404528 233385
rect 482224 233373 482230 233385
rect 404522 233345 482230 233373
rect 404522 233333 404528 233345
rect 482224 233333 482230 233345
rect 482282 233333 482288 233385
rect 142480 233259 142486 233311
rect 142538 233299 142544 233311
rect 142538 233271 144062 233299
rect 142538 233259 142544 233271
rect 144034 233225 144062 233271
rect 144112 233259 144118 233311
rect 144170 233299 144176 233311
rect 168400 233299 168406 233311
rect 144170 233271 168406 233299
rect 144170 233259 144176 233271
rect 168400 233259 168406 233271
rect 168458 233259 168464 233311
rect 283120 233259 283126 233311
rect 283178 233299 283184 233311
rect 372304 233299 372310 233311
rect 283178 233271 372310 233299
rect 283178 233259 283184 233271
rect 372304 233259 372310 233271
rect 372362 233259 372368 233311
rect 402640 233259 402646 233311
rect 402698 233299 402704 233311
rect 402928 233299 402934 233311
rect 402698 233271 402934 233299
rect 402698 233259 402704 233271
rect 402928 233259 402934 233271
rect 402986 233259 402992 233311
rect 403024 233259 403030 233311
rect 403082 233299 403088 233311
rect 403216 233299 403222 233311
rect 403082 233271 403222 233299
rect 403082 233259 403088 233271
rect 403216 233259 403222 233271
rect 403274 233259 403280 233311
rect 409360 233299 409366 233311
rect 406066 233271 409366 233299
rect 147184 233225 147190 233237
rect 144034 233197 147190 233225
rect 147184 233185 147190 233197
rect 147242 233185 147248 233237
rect 283504 233185 283510 233237
rect 283562 233225 283568 233237
rect 388720 233225 388726 233237
rect 283562 233197 388726 233225
rect 283562 233185 283568 233197
rect 388720 233185 388726 233197
rect 388778 233185 388784 233237
rect 399760 233185 399766 233237
rect 399818 233225 399824 233237
rect 406066 233225 406094 233271
rect 409360 233259 409366 233271
rect 409418 233259 409424 233311
rect 409456 233259 409462 233311
rect 409514 233299 409520 233311
rect 411856 233299 411862 233311
rect 409514 233271 411862 233299
rect 409514 233259 409520 233271
rect 411856 233259 411862 233271
rect 411914 233259 411920 233311
rect 411952 233259 411958 233311
rect 412010 233299 412016 233311
rect 415408 233299 415414 233311
rect 412010 233271 415414 233299
rect 412010 233259 412016 233271
rect 415408 233259 415414 233271
rect 415466 233259 415472 233311
rect 415504 233259 415510 233311
rect 415562 233299 415568 233311
rect 443536 233299 443542 233311
rect 415562 233271 443542 233299
rect 415562 233259 415568 233271
rect 443536 233259 443542 233271
rect 443594 233259 443600 233311
rect 444112 233259 444118 233311
rect 444170 233299 444176 233311
rect 481456 233299 481462 233311
rect 444170 233271 481462 233299
rect 444170 233259 444176 233271
rect 481456 233259 481462 233271
rect 481514 233259 481520 233311
rect 456400 233225 456406 233237
rect 399818 233197 406094 233225
rect 406210 233197 443870 233225
rect 399818 233185 399824 233197
rect 283216 233111 283222 233163
rect 283274 233151 283280 233163
rect 386512 233151 386518 233163
rect 283274 233123 386518 233151
rect 283274 233111 283280 233123
rect 386512 233111 386518 233123
rect 386570 233111 386576 233163
rect 402352 233111 402358 233163
rect 402410 233151 402416 233163
rect 406210 233151 406238 233197
rect 402410 233123 406238 233151
rect 402410 233111 402416 233123
rect 406672 233111 406678 233163
rect 406730 233151 406736 233163
rect 407536 233151 407542 233163
rect 406730 233123 407542 233151
rect 406730 233111 406736 233123
rect 407536 233111 407542 233123
rect 407594 233111 407600 233163
rect 410224 233111 410230 233163
rect 410282 233151 410288 233163
rect 421648 233151 421654 233163
rect 410282 233123 421654 233151
rect 410282 233111 410288 233123
rect 421648 233111 421654 233123
rect 421706 233111 421712 233163
rect 424144 233111 424150 233163
rect 424202 233151 424208 233163
rect 440272 233151 440278 233163
rect 424202 233123 440278 233151
rect 424202 233111 424208 233123
rect 440272 233111 440278 233123
rect 440330 233111 440336 233163
rect 443842 233151 443870 233197
rect 456034 233197 456406 233225
rect 456034 233151 456062 233197
rect 456400 233185 456406 233197
rect 456458 233185 456464 233237
rect 443842 233123 456062 233151
rect 456112 233111 456118 233163
rect 456170 233151 456176 233163
rect 463408 233151 463414 233163
rect 456170 233123 463414 233151
rect 456170 233111 456176 233123
rect 463408 233111 463414 233123
rect 463466 233111 463472 233163
rect 286384 233037 286390 233089
rect 286442 233077 286448 233089
rect 386128 233077 386134 233089
rect 286442 233049 386134 233077
rect 286442 233037 286448 233049
rect 386128 233037 386134 233049
rect 386186 233037 386192 233089
rect 401008 233037 401014 233089
rect 401066 233077 401072 233089
rect 407056 233077 407062 233089
rect 401066 233049 407062 233077
rect 401066 233037 401072 233049
rect 407056 233037 407062 233049
rect 407114 233037 407120 233089
rect 407152 233037 407158 233089
rect 407210 233077 407216 233089
rect 413968 233077 413974 233089
rect 407210 233049 413974 233077
rect 407210 233037 407216 233049
rect 413968 233037 413974 233049
rect 414026 233037 414032 233089
rect 414160 233037 414166 233089
rect 414218 233077 414224 233089
rect 414218 233049 418814 233077
rect 414218 233037 414224 233049
rect 349072 232963 349078 233015
rect 349130 233003 349136 233015
rect 414544 233003 414550 233015
rect 349130 232975 414550 233003
rect 349130 232963 349136 232975
rect 414544 232963 414550 232975
rect 414602 232963 414608 233015
rect 415024 232963 415030 233015
rect 415082 233003 415088 233015
rect 417904 233003 417910 233015
rect 415082 232975 417910 233003
rect 415082 232963 415088 232975
rect 417904 232963 417910 232975
rect 417962 232963 417968 233015
rect 418786 233003 418814 233049
rect 418960 233037 418966 233089
rect 419018 233077 419024 233089
rect 443536 233077 443542 233089
rect 419018 233049 443542 233077
rect 419018 233037 419024 233049
rect 443536 233037 443542 233049
rect 443594 233037 443600 233089
rect 462352 233077 462358 233089
rect 443650 233049 462358 233077
rect 443650 233003 443678 233049
rect 462352 233037 462358 233049
rect 462410 233037 462416 233089
rect 470608 233037 470614 233089
rect 470666 233077 470672 233089
rect 473008 233077 473014 233089
rect 470666 233049 473014 233077
rect 470666 233037 470672 233049
rect 473008 233037 473014 233049
rect 473066 233037 473072 233089
rect 418786 232975 443678 233003
rect 443824 232963 443830 233015
rect 443882 233003 443888 233015
rect 454576 233003 454582 233015
rect 443882 232975 454582 233003
rect 443882 232963 443888 232975
rect 454576 232963 454582 232975
rect 454634 232963 454640 233015
rect 336496 232889 336502 232941
rect 336554 232929 336560 232941
rect 398704 232929 398710 232941
rect 336554 232901 398710 232929
rect 336554 232889 336560 232901
rect 398704 232889 398710 232901
rect 398762 232889 398768 232941
rect 398800 232889 398806 232941
rect 398858 232929 398864 232941
rect 418960 232929 418966 232941
rect 398858 232901 418966 232929
rect 398858 232889 398864 232901
rect 418960 232889 418966 232901
rect 419018 232889 419024 232941
rect 419152 232889 419158 232941
rect 419210 232929 419216 232941
rect 424528 232929 424534 232941
rect 419210 232901 424534 232929
rect 419210 232889 419216 232901
rect 424528 232889 424534 232901
rect 424586 232889 424592 232941
rect 424816 232889 424822 232941
rect 424874 232929 424880 232941
rect 468976 232929 468982 232941
rect 424874 232901 468982 232929
rect 424874 232889 424880 232901
rect 468976 232889 468982 232901
rect 469034 232889 469040 232941
rect 348688 232815 348694 232867
rect 348746 232855 348752 232867
rect 414640 232855 414646 232867
rect 348746 232827 414646 232855
rect 348746 232815 348752 232827
rect 414640 232815 414646 232827
rect 414698 232815 414704 232867
rect 414736 232815 414742 232867
rect 414794 232855 414800 232867
rect 443632 232855 443638 232867
rect 414794 232827 443638 232855
rect 414794 232815 414800 232827
rect 443632 232815 443638 232827
rect 443690 232815 443696 232867
rect 443728 232815 443734 232867
rect 443786 232815 443792 232867
rect 443824 232815 443830 232867
rect 443882 232855 443888 232867
rect 455344 232855 455350 232867
rect 443882 232827 455350 232855
rect 443882 232815 443888 232827
rect 455344 232815 455350 232827
rect 455402 232815 455408 232867
rect 283408 232741 283414 232793
rect 283466 232781 283472 232793
rect 363376 232781 363382 232793
rect 283466 232753 363382 232781
rect 283466 232741 283472 232753
rect 363376 232741 363382 232753
rect 363434 232741 363440 232793
rect 364816 232741 364822 232793
rect 364874 232781 364880 232793
rect 374320 232781 374326 232793
rect 364874 232753 374326 232781
rect 364874 232741 364880 232753
rect 374320 232741 374326 232753
rect 374378 232741 374384 232793
rect 398704 232741 398710 232793
rect 398762 232781 398768 232793
rect 413584 232781 413590 232793
rect 398762 232753 413590 232781
rect 398762 232741 398768 232753
rect 413584 232741 413590 232753
rect 413642 232741 413648 232793
rect 443536 232781 443542 232793
rect 414082 232753 443542 232781
rect 321808 232667 321814 232719
rect 321866 232707 321872 232719
rect 409648 232707 409654 232719
rect 321866 232679 409654 232707
rect 321866 232667 321872 232679
rect 409648 232667 409654 232679
rect 409706 232667 409712 232719
rect 409744 232667 409750 232719
rect 409802 232707 409808 232719
rect 413968 232707 413974 232719
rect 409802 232679 413974 232707
rect 409802 232667 409808 232679
rect 413968 232667 413974 232679
rect 414026 232667 414032 232719
rect 141136 232593 141142 232645
rect 141194 232633 141200 232645
rect 141712 232633 141718 232645
rect 141194 232605 141718 232633
rect 141194 232593 141200 232605
rect 141712 232593 141718 232605
rect 141770 232593 141776 232645
rect 326992 232593 326998 232645
rect 327050 232633 327056 232645
rect 399952 232633 399958 232645
rect 327050 232605 399958 232633
rect 327050 232593 327056 232605
rect 399952 232593 399958 232605
rect 400010 232593 400016 232645
rect 400048 232593 400054 232645
rect 400106 232633 400112 232645
rect 414082 232633 414110 232753
rect 443536 232741 443542 232753
rect 443594 232741 443600 232793
rect 443746 232781 443774 232815
rect 461584 232781 461590 232793
rect 443746 232753 461590 232781
rect 461584 232741 461590 232753
rect 461642 232741 461648 232793
rect 414256 232667 414262 232719
rect 414314 232707 414320 232719
rect 415024 232707 415030 232719
rect 414314 232679 415030 232707
rect 414314 232667 414320 232679
rect 415024 232667 415030 232679
rect 415082 232667 415088 232719
rect 415408 232667 415414 232719
rect 415466 232707 415472 232719
rect 415466 232679 424478 232707
rect 415466 232667 415472 232679
rect 400106 232605 414110 232633
rect 400106 232593 400112 232605
rect 417136 232593 417142 232645
rect 417194 232633 417200 232645
rect 424450 232633 424478 232679
rect 424528 232667 424534 232719
rect 424586 232707 424592 232719
rect 443632 232707 443638 232719
rect 424586 232679 443638 232707
rect 424586 232667 424592 232679
rect 443632 232667 443638 232679
rect 443690 232667 443696 232719
rect 461200 232707 461206 232719
rect 443746 232679 461206 232707
rect 443746 232633 443774 232679
rect 461200 232667 461206 232679
rect 461258 232667 461264 232719
rect 417194 232605 423134 232633
rect 424450 232605 443774 232633
rect 417194 232593 417200 232605
rect 326224 232519 326230 232571
rect 326282 232559 326288 232571
rect 417808 232559 417814 232571
rect 326282 232531 417814 232559
rect 326282 232519 326288 232531
rect 417808 232519 417814 232531
rect 417866 232519 417872 232571
rect 417904 232519 417910 232571
rect 417962 232559 417968 232571
rect 421168 232559 421174 232571
rect 417962 232531 421174 232559
rect 417962 232519 417968 232531
rect 421168 232519 421174 232531
rect 421226 232519 421232 232571
rect 327664 232445 327670 232497
rect 327722 232485 327728 232497
rect 391120 232485 391126 232497
rect 327722 232457 391126 232485
rect 327722 232445 327728 232457
rect 391120 232445 391126 232457
rect 391178 232445 391184 232497
rect 418000 232485 418006 232497
rect 391330 232457 418006 232485
rect 341584 232371 341590 232423
rect 341642 232411 341648 232423
rect 391330 232411 391358 232457
rect 418000 232445 418006 232457
rect 418058 232445 418064 232497
rect 418288 232445 418294 232497
rect 418346 232485 418352 232497
rect 423106 232485 423134 232605
rect 423472 232519 423478 232571
rect 423530 232559 423536 232571
rect 443824 232559 443830 232571
rect 423530 232531 443830 232559
rect 423530 232519 423536 232531
rect 443824 232519 443830 232531
rect 443882 232519 443888 232571
rect 443938 232531 444158 232559
rect 443938 232485 443966 232531
rect 418346 232457 423038 232485
rect 423106 232457 443966 232485
rect 444130 232485 444158 232531
rect 453712 232519 453718 232571
rect 453770 232559 453776 232571
rect 467344 232559 467350 232571
rect 453770 232531 467350 232559
rect 453770 232519 453776 232531
rect 467344 232519 467350 232531
rect 467402 232519 467408 232571
rect 463792 232485 463798 232497
rect 444130 232457 463798 232485
rect 418346 232445 418352 232457
rect 341642 232383 391358 232411
rect 341642 232371 341648 232383
rect 391408 232371 391414 232423
rect 391466 232411 391472 232423
rect 418384 232411 418390 232423
rect 391466 232383 418390 232411
rect 391466 232371 391472 232383
rect 418384 232371 418390 232383
rect 418442 232371 418448 232423
rect 423010 232411 423038 232457
rect 463792 232445 463798 232457
rect 463850 232445 463856 232497
rect 423472 232411 423478 232423
rect 423010 232383 423478 232411
rect 423472 232371 423478 232383
rect 423530 232371 423536 232423
rect 423760 232371 423766 232423
rect 423818 232411 423824 232423
rect 443536 232411 443542 232423
rect 423818 232383 443542 232411
rect 423818 232371 423824 232383
rect 443536 232371 443542 232383
rect 443594 232371 443600 232423
rect 444400 232371 444406 232423
rect 444458 232411 444464 232423
rect 453328 232411 453334 232423
rect 444458 232383 453334 232411
rect 444458 232371 444464 232383
rect 453328 232371 453334 232383
rect 453386 232371 453392 232423
rect 453424 232371 453430 232423
rect 453482 232411 453488 232423
rect 467824 232411 467830 232423
rect 453482 232383 467830 232411
rect 453482 232371 453488 232383
rect 467824 232371 467830 232383
rect 467882 232371 467888 232423
rect 337648 232297 337654 232349
rect 337706 232337 337712 232349
rect 428752 232337 428758 232349
rect 337706 232309 428758 232337
rect 337706 232297 337712 232309
rect 428752 232297 428758 232309
rect 428810 232297 428816 232349
rect 429232 232297 429238 232349
rect 429290 232337 429296 232349
rect 473392 232337 473398 232349
rect 429290 232309 473398 232337
rect 429290 232297 429296 232309
rect 473392 232297 473398 232309
rect 473450 232297 473456 232349
rect 335824 232223 335830 232275
rect 335882 232263 335888 232275
rect 426256 232263 426262 232275
rect 335882 232235 426262 232263
rect 335882 232223 335888 232235
rect 426256 232223 426262 232235
rect 426314 232223 426320 232275
rect 426640 232223 426646 232275
rect 426698 232263 426704 232275
rect 470800 232263 470806 232275
rect 426698 232235 470806 232263
rect 426698 232223 426704 232235
rect 470800 232223 470806 232235
rect 470858 232223 470864 232275
rect 324784 232149 324790 232201
rect 324842 232189 324848 232201
rect 391216 232189 391222 232201
rect 324842 232161 391222 232189
rect 324842 232149 324848 232161
rect 391216 232149 391222 232161
rect 391274 232149 391280 232201
rect 417232 232189 417238 232201
rect 391330 232161 417238 232189
rect 324016 232075 324022 232127
rect 324074 232115 324080 232127
rect 391330 232115 391358 232161
rect 417232 232149 417238 232161
rect 417290 232149 417296 232201
rect 420304 232149 420310 232201
rect 420362 232189 420368 232201
rect 462736 232189 462742 232201
rect 420362 232161 462742 232189
rect 420362 232149 420368 232161
rect 462736 232149 462742 232161
rect 462794 232149 462800 232201
rect 324074 232087 391358 232115
rect 324074 232075 324080 232087
rect 398800 232075 398806 232127
rect 398858 232115 398864 232127
rect 419632 232115 419638 232127
rect 398858 232087 419638 232115
rect 398858 232075 398864 232087
rect 419632 232075 419638 232087
rect 419690 232075 419696 232127
rect 421168 232075 421174 232127
rect 421226 232115 421232 232127
rect 421840 232115 421846 232127
rect 421226 232087 421846 232115
rect 421226 232075 421232 232087
rect 421840 232075 421846 232087
rect 421898 232075 421904 232127
rect 422608 232075 422614 232127
rect 422666 232115 422672 232127
rect 466768 232115 466774 232127
rect 422666 232087 466774 232115
rect 422666 232075 422672 232087
rect 466768 232075 466774 232087
rect 466826 232075 466832 232127
rect 323248 232001 323254 232053
rect 323306 232041 323312 232053
rect 419248 232041 419254 232053
rect 323306 232013 419254 232041
rect 323306 232001 323312 232013
rect 419248 232001 419254 232013
rect 419306 232001 419312 232053
rect 420400 232001 420406 232053
rect 420458 232041 420464 232053
rect 464560 232041 464566 232053
rect 420458 232013 464566 232041
rect 420458 232001 420464 232013
rect 464560 232001 464566 232013
rect 464618 232001 464624 232053
rect 475120 232001 475126 232053
rect 475178 232041 475184 232053
rect 505744 232041 505750 232053
rect 475178 232013 505750 232041
rect 475178 232001 475184 232013
rect 505744 232001 505750 232013
rect 505802 232001 505808 232053
rect 335056 231927 335062 231979
rect 335114 231967 335120 231979
rect 431824 231967 431830 231979
rect 335114 231939 431830 231967
rect 335114 231927 335120 231939
rect 431824 231927 431830 231939
rect 431882 231927 431888 231979
rect 432208 231927 432214 231979
rect 432266 231967 432272 231979
rect 476272 231967 476278 231979
rect 432266 231939 476278 231967
rect 432266 231927 432272 231939
rect 476272 231927 476278 231939
rect 476330 231927 476336 231979
rect 322480 231853 322486 231905
rect 322538 231893 322544 231905
rect 398800 231893 398806 231905
rect 322538 231865 398806 231893
rect 322538 231853 322544 231865
rect 398800 231853 398806 231865
rect 398858 231853 398864 231905
rect 399952 231853 399958 231905
rect 400010 231893 400016 231905
rect 408880 231893 408886 231905
rect 400010 231865 408886 231893
rect 400010 231853 400016 231865
rect 408880 231853 408886 231865
rect 408938 231853 408944 231905
rect 411184 231853 411190 231905
rect 411242 231893 411248 231905
rect 419152 231893 419158 231905
rect 411242 231865 419158 231893
rect 411242 231853 411248 231865
rect 419152 231853 419158 231865
rect 419210 231853 419216 231905
rect 419344 231853 419350 231905
rect 419402 231893 419408 231905
rect 464944 231893 464950 231905
rect 419402 231865 464950 231893
rect 419402 231853 419408 231865
rect 464944 231853 464950 231865
rect 465002 231853 465008 231905
rect 466576 231853 466582 231905
rect 466634 231893 466640 231905
rect 504976 231893 504982 231905
rect 466634 231865 504982 231893
rect 466634 231853 466640 231865
rect 504976 231853 504982 231865
rect 505034 231853 505040 231905
rect 333616 231779 333622 231831
rect 333674 231819 333680 231831
rect 436048 231819 436054 231831
rect 333674 231791 436054 231819
rect 333674 231779 333680 231791
rect 436048 231779 436054 231791
rect 436106 231779 436112 231831
rect 437680 231779 437686 231831
rect 437738 231819 437744 231831
rect 503536 231819 503542 231831
rect 437738 231791 503542 231819
rect 437738 231779 437744 231791
rect 503536 231779 503542 231791
rect 503594 231779 503600 231831
rect 285904 231705 285910 231757
rect 285962 231745 285968 231757
rect 363664 231745 363670 231757
rect 285962 231717 363670 231745
rect 285962 231705 285968 231717
rect 363664 231705 363670 231717
rect 363722 231705 363728 231757
rect 397936 231705 397942 231757
rect 397994 231745 398000 231757
rect 403888 231745 403894 231757
rect 397994 231717 403894 231745
rect 397994 231705 398000 231717
rect 403888 231705 403894 231717
rect 403946 231705 403952 231757
rect 403984 231705 403990 231757
rect 404042 231745 404048 231757
rect 405232 231745 405238 231757
rect 404042 231717 405238 231745
rect 404042 231705 404048 231717
rect 405232 231705 405238 231717
rect 405290 231705 405296 231757
rect 406192 231705 406198 231757
rect 406250 231745 406256 231757
rect 406250 231717 419006 231745
rect 406250 231705 406256 231717
rect 286096 231631 286102 231683
rect 286154 231671 286160 231683
rect 361168 231671 361174 231683
rect 286154 231643 361174 231671
rect 286154 231631 286160 231643
rect 361168 231631 361174 231643
rect 361226 231631 361232 231683
rect 394672 231631 394678 231683
rect 394730 231671 394736 231683
rect 394730 231643 406718 231671
rect 394730 231631 394736 231643
rect 336880 231557 336886 231609
rect 336938 231597 336944 231609
rect 404272 231597 404278 231609
rect 336938 231569 404278 231597
rect 336938 231557 336944 231569
rect 404272 231557 404278 231569
rect 404330 231557 404336 231609
rect 406690 231597 406718 231643
rect 406768 231631 406774 231683
rect 406826 231671 406832 231683
rect 406826 231643 410078 231671
rect 406826 231631 406832 231643
rect 406960 231597 406966 231609
rect 406690 231569 406966 231597
rect 406960 231557 406966 231569
rect 407018 231557 407024 231609
rect 410050 231597 410078 231643
rect 410128 231631 410134 231683
rect 410186 231671 410192 231683
rect 418096 231671 418102 231683
rect 410186 231643 418102 231671
rect 410186 231631 410192 231643
rect 418096 231631 418102 231643
rect 418154 231631 418160 231683
rect 418978 231671 419006 231717
rect 419056 231705 419062 231757
rect 419114 231745 419120 231757
rect 454192 231745 454198 231757
rect 419114 231717 454198 231745
rect 419114 231705 419120 231717
rect 454192 231705 454198 231717
rect 454250 231705 454256 231757
rect 458320 231671 458326 231683
rect 418978 231643 458326 231671
rect 458320 231631 458326 231643
rect 458378 231631 458384 231683
rect 420496 231597 420502 231609
rect 410050 231569 420502 231597
rect 420496 231557 420502 231569
rect 420554 231557 420560 231609
rect 422032 231557 422038 231609
rect 422090 231597 422096 231609
rect 428560 231597 428566 231609
rect 422090 231569 428566 231597
rect 422090 231557 422096 231569
rect 428560 231557 428566 231569
rect 428618 231557 428624 231609
rect 430672 231557 430678 231609
rect 430730 231597 430736 231609
rect 439504 231597 439510 231609
rect 430730 231569 439510 231597
rect 430730 231557 430736 231569
rect 439504 231557 439510 231569
rect 439562 231557 439568 231609
rect 439600 231557 439606 231609
rect 439658 231597 439664 231609
rect 458608 231597 458614 231609
rect 439658 231569 458614 231597
rect 439658 231557 439664 231569
rect 458608 231557 458614 231569
rect 458666 231557 458672 231609
rect 286672 231483 286678 231535
rect 286730 231523 286736 231535
rect 362608 231523 362614 231535
rect 286730 231495 362614 231523
rect 286730 231483 286736 231495
rect 362608 231483 362614 231495
rect 362666 231483 362672 231535
rect 363760 231483 363766 231535
rect 363818 231523 363824 231535
rect 375472 231523 375478 231535
rect 363818 231495 375478 231523
rect 363818 231483 363824 231495
rect 375472 231483 375478 231495
rect 375530 231483 375536 231535
rect 386512 231483 386518 231535
rect 386570 231523 386576 231535
rect 411760 231523 411766 231535
rect 386570 231495 411766 231523
rect 386570 231483 386576 231495
rect 411760 231483 411766 231495
rect 411818 231483 411824 231535
rect 413488 231483 413494 231535
rect 413546 231523 413552 231535
rect 421168 231523 421174 231535
rect 413546 231495 421174 231523
rect 413546 231483 413552 231495
rect 421168 231483 421174 231495
rect 421226 231483 421232 231535
rect 421648 231483 421654 231535
rect 421706 231523 421712 231535
rect 427600 231523 427606 231535
rect 421706 231495 427606 231523
rect 421706 231483 421712 231495
rect 427600 231483 427606 231495
rect 427658 231483 427664 231535
rect 460144 231523 460150 231535
rect 427714 231495 460150 231523
rect 284560 231409 284566 231461
rect 284618 231449 284624 231461
rect 353392 231449 353398 231461
rect 284618 231421 353398 231449
rect 284618 231409 284624 231421
rect 353392 231409 353398 231421
rect 353450 231409 353456 231461
rect 362992 231409 362998 231461
rect 363050 231449 363056 231461
rect 375856 231449 375862 231461
rect 363050 231421 375862 231449
rect 363050 231409 363056 231421
rect 375856 231409 375862 231421
rect 375914 231409 375920 231461
rect 391408 231409 391414 231461
rect 391466 231449 391472 231461
rect 403600 231449 403606 231461
rect 391466 231421 403606 231449
rect 391466 231409 391472 231421
rect 403600 231409 403606 231421
rect 403658 231409 403664 231461
rect 403696 231409 403702 231461
rect 403754 231449 403760 231461
rect 423376 231449 423382 231461
rect 403754 231421 423382 231449
rect 403754 231409 403760 231421
rect 423376 231409 423382 231421
rect 423434 231409 423440 231461
rect 426352 231409 426358 231461
rect 426410 231449 426416 231461
rect 427714 231449 427742 231495
rect 460144 231483 460150 231495
rect 460202 231483 460208 231535
rect 426410 231421 427742 231449
rect 426410 231409 426416 231421
rect 431344 231409 431350 231461
rect 431402 231449 431408 231461
rect 468592 231449 468598 231461
rect 431402 231421 468598 231449
rect 431402 231409 431408 231421
rect 468592 231409 468598 231421
rect 468650 231409 468656 231461
rect 351280 231335 351286 231387
rect 351338 231375 351344 231387
rect 372688 231375 372694 231387
rect 351338 231347 372694 231375
rect 351338 231335 351344 231347
rect 372688 231335 372694 231347
rect 372746 231335 372752 231387
rect 391600 231335 391606 231387
rect 391658 231375 391664 231387
rect 413776 231375 413782 231387
rect 391658 231347 413782 231375
rect 391658 231335 391664 231347
rect 413776 231335 413782 231347
rect 413834 231335 413840 231387
rect 413968 231335 413974 231387
rect 414026 231375 414032 231387
rect 414026 231347 422174 231375
rect 414026 231335 414032 231347
rect 338032 231261 338038 231313
rect 338090 231301 338096 231313
rect 391216 231301 391222 231313
rect 338090 231273 391222 231301
rect 338090 231261 338096 231273
rect 391216 231261 391222 231273
rect 391274 231261 391280 231313
rect 414448 231301 414454 231313
rect 391330 231273 414454 231301
rect 349744 231187 349750 231239
rect 349802 231227 349808 231239
rect 373744 231227 373750 231239
rect 349802 231199 373750 231227
rect 349802 231187 349808 231199
rect 373744 231187 373750 231199
rect 373802 231187 373808 231239
rect 384784 231187 384790 231239
rect 384842 231227 384848 231239
rect 391330 231227 391358 231273
rect 414448 231261 414454 231273
rect 414506 231261 414512 231313
rect 417616 231261 417622 231313
rect 417674 231301 417680 231313
rect 420208 231301 420214 231313
rect 417674 231273 420214 231301
rect 417674 231261 417680 231273
rect 420208 231261 420214 231273
rect 420266 231261 420272 231313
rect 422032 231301 422038 231313
rect 420322 231273 422038 231301
rect 417040 231227 417046 231239
rect 384842 231199 391358 231227
rect 391426 231199 417046 231227
rect 384842 231187 384848 231199
rect 282640 231113 282646 231165
rect 282698 231153 282704 231165
rect 362992 231153 362998 231165
rect 282698 231125 362998 231153
rect 282698 231113 282704 231125
rect 362992 231113 362998 231125
rect 363050 231113 363056 231165
rect 391120 231113 391126 231165
rect 391178 231153 391184 231165
rect 391426 231153 391454 231199
rect 417040 231187 417046 231199
rect 417098 231187 417104 231239
rect 417712 231187 417718 231239
rect 417770 231227 417776 231239
rect 420322 231227 420350 231273
rect 422032 231261 422038 231273
rect 422090 231261 422096 231313
rect 422146 231301 422174 231347
rect 422224 231335 422230 231387
rect 422282 231375 422288 231387
rect 426448 231375 426454 231387
rect 422282 231347 426454 231375
rect 422282 231335 422288 231347
rect 426448 231335 426454 231347
rect 426506 231335 426512 231387
rect 428176 231335 428182 231387
rect 428234 231375 428240 231387
rect 472240 231375 472246 231387
rect 428234 231347 472246 231375
rect 428234 231335 428240 231347
rect 472240 231335 472246 231347
rect 472298 231335 472304 231387
rect 426352 231301 426358 231313
rect 422146 231273 426358 231301
rect 426352 231261 426358 231273
rect 426410 231261 426416 231313
rect 426640 231261 426646 231313
rect 426698 231301 426704 231313
rect 470416 231301 470422 231313
rect 426698 231273 470422 231301
rect 426698 231261 426704 231273
rect 470416 231261 470422 231273
rect 470474 231261 470480 231313
rect 417770 231199 420350 231227
rect 417770 231187 417776 231199
rect 420592 231187 420598 231239
rect 420650 231227 420656 231239
rect 439408 231227 439414 231239
rect 420650 231199 439414 231227
rect 420650 231187 420656 231199
rect 439408 231187 439414 231199
rect 439466 231187 439472 231239
rect 439504 231187 439510 231239
rect 439562 231227 439568 231239
rect 465616 231227 465622 231239
rect 439562 231199 465622 231227
rect 439562 231187 439568 231199
rect 465616 231187 465622 231199
rect 465674 231187 465680 231239
rect 391178 231125 391454 231153
rect 391178 231113 391184 231125
rect 393040 231113 393046 231165
rect 393098 231153 393104 231165
rect 431920 231153 431926 231165
rect 393098 231125 431926 231153
rect 393098 231113 393104 231125
rect 431920 231113 431926 231125
rect 431978 231113 431984 231165
rect 432016 231113 432022 231165
rect 432074 231153 432080 231165
rect 439216 231153 439222 231165
rect 432074 231125 439222 231153
rect 432074 231113 432080 231125
rect 439216 231113 439222 231125
rect 439274 231113 439280 231165
rect 473776 231153 473782 231165
rect 439330 231125 473782 231153
rect 286960 231039 286966 231091
rect 287018 231079 287024 231091
rect 364048 231079 364054 231091
rect 287018 231051 364054 231079
rect 287018 231039 287024 231051
rect 364048 231039 364054 231051
rect 364106 231039 364112 231091
rect 390928 231039 390934 231091
rect 390986 231079 390992 231091
rect 403696 231079 403702 231091
rect 390986 231051 403702 231079
rect 390986 231039 390992 231051
rect 403696 231039 403702 231051
rect 403754 231039 403760 231091
rect 403888 231039 403894 231091
rect 403946 231079 403952 231091
rect 419056 231079 419062 231091
rect 403946 231051 419062 231079
rect 403946 231039 403952 231051
rect 419056 231039 419062 231051
rect 419114 231039 419120 231091
rect 421552 231039 421558 231091
rect 421610 231079 421616 231091
rect 421610 231051 427934 231079
rect 421610 231039 421616 231051
rect 345616 230965 345622 231017
rect 345674 231005 345680 231017
rect 355984 231005 355990 231017
rect 345674 230977 355990 231005
rect 345674 230965 345680 230977
rect 355984 230965 355990 230977
rect 356042 230965 356048 231017
rect 356752 230965 356758 231017
rect 356810 231005 356816 231017
rect 427312 231005 427318 231017
rect 356810 230977 427318 231005
rect 356810 230965 356816 230977
rect 427312 230965 427318 230977
rect 427370 230965 427376 231017
rect 353200 230891 353206 230943
rect 353258 230931 353264 230943
rect 365488 230931 365494 230943
rect 353258 230903 365494 230931
rect 353258 230891 353264 230903
rect 365488 230891 365494 230903
rect 365546 230891 365552 230943
rect 389872 230891 389878 230943
rect 389930 230931 389936 230943
rect 389930 230903 409118 230931
rect 389930 230891 389936 230903
rect 345904 230817 345910 230869
rect 345962 230857 345968 230869
rect 364432 230857 364438 230869
rect 345962 230829 364438 230857
rect 345962 230817 345968 230829
rect 364432 230817 364438 230829
rect 364490 230817 364496 230869
rect 392080 230817 392086 230869
rect 392138 230857 392144 230869
rect 403696 230857 403702 230869
rect 392138 230829 403702 230857
rect 392138 230817 392144 230829
rect 403696 230817 403702 230829
rect 403754 230817 403760 230869
rect 409090 230857 409118 230903
rect 409168 230891 409174 230943
rect 409226 230931 409232 230943
rect 427792 230931 427798 230943
rect 409226 230903 427798 230931
rect 409226 230891 409232 230903
rect 427792 230891 427798 230903
rect 427850 230891 427856 230943
rect 427906 230931 427934 231051
rect 427984 231039 427990 231091
rect 428042 231079 428048 231091
rect 428944 231079 428950 231091
rect 428042 231051 428950 231079
rect 428042 231039 428048 231051
rect 428944 231039 428950 231051
rect 429002 231039 429008 231091
rect 429616 231039 429622 231091
rect 429674 231079 429680 231091
rect 439330 231079 439358 231125
rect 473776 231113 473782 231125
rect 473834 231113 473840 231165
rect 466000 231079 466006 231091
rect 429674 231051 439358 231079
rect 439618 231051 466006 231079
rect 429674 231039 429680 231051
rect 428560 230965 428566 231017
rect 428618 231005 428624 231017
rect 439504 231005 439510 231017
rect 428618 230977 439510 231005
rect 428618 230965 428624 230977
rect 439504 230965 439510 230977
rect 439562 230965 439568 231017
rect 439618 230931 439646 231051
rect 466000 231039 466006 231051
rect 466058 231039 466064 231091
rect 440272 230965 440278 231017
rect 440330 231005 440336 231017
rect 468208 231005 468214 231017
rect 440330 230977 468214 231005
rect 440330 230965 440336 230977
rect 468208 230965 468214 230977
rect 468266 230965 468272 231017
rect 427906 230903 439646 230931
rect 439696 230891 439702 230943
rect 439754 230931 439760 230943
rect 474064 230931 474070 230943
rect 439754 230903 474070 230931
rect 439754 230891 439760 230903
rect 474064 230891 474070 230903
rect 474122 230891 474128 230943
rect 426064 230857 426070 230869
rect 409090 230829 426070 230857
rect 426064 230817 426070 230829
rect 426122 230817 426128 230869
rect 430000 230817 430006 230869
rect 430058 230857 430064 230869
rect 431920 230857 431926 230869
rect 430058 230829 431926 230857
rect 430058 230817 430064 230829
rect 431920 230817 431926 230829
rect 431978 230817 431984 230869
rect 432592 230817 432598 230869
rect 432650 230857 432656 230869
rect 476656 230857 476662 230869
rect 432650 230829 476662 230857
rect 432650 230817 432656 230829
rect 476656 230817 476662 230829
rect 476714 230817 476720 230869
rect 389488 230743 389494 230795
rect 389546 230783 389552 230795
rect 403600 230783 403606 230795
rect 389546 230755 403606 230783
rect 389546 230743 389552 230755
rect 403600 230743 403606 230755
rect 403658 230743 403664 230795
rect 409072 230783 409078 230795
rect 403714 230755 409078 230783
rect 387664 230669 387670 230721
rect 387722 230709 387728 230721
rect 403312 230709 403318 230721
rect 387722 230681 403318 230709
rect 387722 230669 387728 230681
rect 403312 230669 403318 230681
rect 403370 230669 403376 230721
rect 403714 230709 403742 230755
rect 409072 230743 409078 230755
rect 409130 230743 409136 230795
rect 426160 230783 426166 230795
rect 409186 230755 426166 230783
rect 403522 230681 403742 230709
rect 155344 230595 155350 230647
rect 155402 230635 155408 230647
rect 156880 230635 156886 230647
rect 155402 230607 156886 230635
rect 155402 230595 155408 230607
rect 156880 230595 156886 230607
rect 156938 230595 156944 230647
rect 391696 230595 391702 230647
rect 391754 230635 391760 230647
rect 403522 230635 403550 230681
rect 403888 230669 403894 230721
rect 403946 230709 403952 230721
rect 409186 230709 409214 230755
rect 426160 230743 426166 230755
rect 426218 230743 426224 230795
rect 426448 230743 426454 230795
rect 426506 230783 426512 230795
rect 466384 230783 466390 230795
rect 426506 230755 466390 230783
rect 426506 230743 426512 230755
rect 466384 230743 466390 230755
rect 466442 230743 466448 230795
rect 403946 230681 409214 230709
rect 403946 230669 403952 230681
rect 409744 230669 409750 230721
rect 409802 230709 409808 230721
rect 414064 230709 414070 230721
rect 409802 230681 414070 230709
rect 409802 230669 409808 230681
rect 414064 230669 414070 230681
rect 414122 230669 414128 230721
rect 415312 230669 415318 230721
rect 415370 230709 415376 230721
rect 419344 230709 419350 230721
rect 415370 230681 419350 230709
rect 415370 230669 415376 230681
rect 419344 230669 419350 230681
rect 419402 230669 419408 230721
rect 427024 230669 427030 230721
rect 427082 230709 427088 230721
rect 471184 230709 471190 230721
rect 427082 230681 471190 230709
rect 427082 230669 427088 230681
rect 471184 230669 471190 230681
rect 471242 230669 471248 230721
rect 391754 230607 403550 230635
rect 391754 230595 391760 230607
rect 403600 230595 403606 230647
rect 403658 230635 403664 230647
rect 423952 230635 423958 230647
rect 403658 230607 423958 230635
rect 403658 230595 403664 230607
rect 423952 230595 423958 230607
rect 424010 230595 424016 230647
rect 456112 230635 456118 230647
rect 426178 230607 456118 230635
rect 383632 230521 383638 230573
rect 383690 230561 383696 230573
rect 425776 230561 425782 230573
rect 383690 230533 425782 230561
rect 383690 230521 383696 230533
rect 425776 230521 425782 230533
rect 425834 230521 425840 230573
rect 426178 230561 426206 230607
rect 456112 230595 456118 230607
rect 456170 230595 456176 230647
rect 425986 230533 426206 230561
rect 144016 230447 144022 230499
rect 144074 230487 144080 230499
rect 194320 230487 194326 230499
rect 144074 230459 194326 230487
rect 144074 230447 144080 230459
rect 194320 230447 194326 230459
rect 194378 230447 194384 230499
rect 360304 230447 360310 230499
rect 360362 230487 360368 230499
rect 379120 230487 379126 230499
rect 360362 230459 379126 230487
rect 360362 230447 360368 230459
rect 379120 230447 379126 230459
rect 379178 230447 379184 230499
rect 402658 230459 403646 230487
rect 140272 230373 140278 230425
rect 140330 230413 140336 230425
rect 141040 230413 141046 230425
rect 140330 230385 141046 230413
rect 140330 230373 140336 230385
rect 141040 230373 141046 230385
rect 141098 230373 141104 230425
rect 147184 230373 147190 230425
rect 147242 230413 147248 230425
rect 207856 230413 207862 230425
rect 147242 230385 207862 230413
rect 147242 230373 147248 230385
rect 207856 230373 207862 230385
rect 207914 230373 207920 230425
rect 285712 230373 285718 230425
rect 285770 230413 285776 230425
rect 369520 230413 369526 230425
rect 285770 230385 369526 230413
rect 285770 230373 285776 230385
rect 369520 230373 369526 230385
rect 369578 230373 369584 230425
rect 371056 230373 371062 230425
rect 371114 230413 371120 230425
rect 372592 230413 372598 230425
rect 371114 230385 372598 230413
rect 371114 230373 371120 230385
rect 372592 230373 372598 230385
rect 372650 230373 372656 230425
rect 395344 230373 395350 230425
rect 395402 230413 395408 230425
rect 402658 230413 402686 230459
rect 395402 230385 402686 230413
rect 395402 230373 395408 230385
rect 402736 230373 402742 230425
rect 402794 230413 402800 230425
rect 403504 230413 403510 230425
rect 402794 230385 403510 230413
rect 402794 230373 402800 230385
rect 403504 230373 403510 230385
rect 403562 230373 403568 230425
rect 403618 230413 403646 230459
rect 403696 230447 403702 230499
rect 403754 230487 403760 230499
rect 409168 230487 409174 230499
rect 403754 230459 409174 230487
rect 403754 230447 403760 230459
rect 409168 230447 409174 230459
rect 409226 230447 409232 230499
rect 409360 230447 409366 230499
rect 409418 230487 409424 230499
rect 417424 230487 417430 230499
rect 409418 230459 417430 230487
rect 409418 230447 409424 230459
rect 417424 230447 417430 230459
rect 417482 230447 417488 230499
rect 417520 230447 417526 230499
rect 417578 230487 417584 230499
rect 425986 230487 426014 230533
rect 427600 230521 427606 230573
rect 427658 230561 427664 230573
rect 457936 230561 457942 230573
rect 427658 230533 457942 230561
rect 427658 230521 427664 230533
rect 457936 230521 457942 230533
rect 457994 230521 458000 230573
rect 417578 230459 426014 230487
rect 417578 230447 417584 230459
rect 430576 230447 430582 230499
rect 430634 230487 430640 230499
rect 440752 230487 440758 230499
rect 430634 230459 440758 230487
rect 430634 230447 430640 230459
rect 440752 230447 440758 230459
rect 440810 230447 440816 230499
rect 442978 230459 443198 230487
rect 410128 230413 410134 230425
rect 403618 230385 410134 230413
rect 410128 230373 410134 230385
rect 410186 230373 410192 230425
rect 411856 230373 411862 230425
rect 411914 230413 411920 230425
rect 428080 230413 428086 230425
rect 411914 230385 428086 230413
rect 411914 230373 411920 230385
rect 428080 230373 428086 230385
rect 428138 230373 428144 230425
rect 428464 230373 428470 230425
rect 428522 230413 428528 230425
rect 439216 230413 439222 230425
rect 428522 230385 439222 230413
rect 428522 230373 428528 230385
rect 439216 230373 439222 230385
rect 439274 230373 439280 230425
rect 439504 230373 439510 230425
rect 439562 230413 439568 230425
rect 442768 230413 442774 230425
rect 439562 230385 442774 230413
rect 439562 230373 439568 230385
rect 442768 230373 442774 230385
rect 442826 230373 442832 230425
rect 149776 230299 149782 230351
rect 149834 230339 149840 230351
rect 207760 230339 207766 230351
rect 149834 230311 207766 230339
rect 149834 230299 149840 230311
rect 207760 230299 207766 230311
rect 207818 230299 207824 230351
rect 283984 230299 283990 230351
rect 284042 230339 284048 230351
rect 357808 230339 357814 230351
rect 284042 230311 357814 230339
rect 284042 230299 284048 230311
rect 357808 230299 357814 230311
rect 357866 230299 357872 230351
rect 367408 230339 367414 230351
rect 357922 230311 367414 230339
rect 152080 230225 152086 230277
rect 152138 230265 152144 230277
rect 208144 230265 208150 230277
rect 152138 230237 208150 230265
rect 152138 230225 152144 230237
rect 208144 230225 208150 230237
rect 208202 230225 208208 230277
rect 283312 230225 283318 230277
rect 283370 230265 283376 230277
rect 357922 230265 357950 230311
rect 367408 230299 367414 230311
rect 367466 230299 367472 230351
rect 367600 230299 367606 230351
rect 367658 230339 367664 230351
rect 370288 230339 370294 230351
rect 367658 230311 370294 230339
rect 367658 230299 367664 230311
rect 370288 230299 370294 230311
rect 370346 230299 370352 230351
rect 370384 230299 370390 230351
rect 370442 230339 370448 230351
rect 372208 230339 372214 230351
rect 370442 230311 372214 230339
rect 370442 230299 370448 230311
rect 372208 230299 372214 230311
rect 372266 230299 372272 230351
rect 393520 230299 393526 230351
rect 393578 230339 393584 230351
rect 402256 230339 402262 230351
rect 393578 230311 402262 230339
rect 393578 230299 393584 230311
rect 402256 230299 402262 230311
rect 402314 230299 402320 230351
rect 402352 230299 402358 230351
rect 402410 230339 402416 230351
rect 404176 230339 404182 230351
rect 402410 230311 404182 230339
rect 402410 230299 402416 230311
rect 404176 230299 404182 230311
rect 404234 230299 404240 230351
rect 404272 230299 404278 230351
rect 404330 230339 404336 230351
rect 442978 230339 443006 230459
rect 404330 230311 443006 230339
rect 443170 230339 443198 230459
rect 446320 230447 446326 230499
rect 446378 230487 446384 230499
rect 465232 230487 465238 230499
rect 446378 230459 465238 230487
rect 446378 230447 446384 230459
rect 465232 230447 465238 230459
rect 465290 230447 465296 230499
rect 443248 230373 443254 230425
rect 443306 230413 443312 230425
rect 495184 230413 495190 230425
rect 443306 230385 495190 230413
rect 443306 230373 443312 230385
rect 495184 230373 495190 230385
rect 495242 230373 495248 230425
rect 495280 230373 495286 230425
rect 495338 230413 495344 230425
rect 500944 230413 500950 230425
rect 495338 230385 500950 230413
rect 495338 230373 495344 230385
rect 500944 230373 500950 230385
rect 501002 230373 501008 230425
rect 451696 230339 451702 230351
rect 443170 230311 451702 230339
rect 404330 230299 404336 230311
rect 451696 230299 451702 230311
rect 451754 230299 451760 230351
rect 451888 230299 451894 230351
rect 451946 230339 451952 230351
rect 463120 230339 463126 230351
rect 451946 230311 463126 230339
rect 451946 230299 451952 230311
rect 463120 230299 463126 230311
rect 463178 230299 463184 230351
rect 368848 230265 368854 230277
rect 283370 230237 357950 230265
rect 358498 230237 368854 230265
rect 283370 230225 283376 230237
rect 166960 230151 166966 230203
rect 167018 230191 167024 230203
rect 212464 230191 212470 230203
rect 167018 230163 212470 230191
rect 167018 230151 167024 230163
rect 212464 230151 212470 230163
rect 212522 230151 212528 230203
rect 285328 230151 285334 230203
rect 285386 230191 285392 230203
rect 358498 230191 358526 230237
rect 368848 230225 368854 230237
rect 368906 230225 368912 230277
rect 370768 230225 370774 230277
rect 370826 230265 370832 230277
rect 373264 230265 373270 230277
rect 370826 230237 373270 230265
rect 370826 230225 370832 230237
rect 373264 230225 373270 230237
rect 373322 230225 373328 230277
rect 373648 230225 373654 230277
rect 373706 230265 373712 230277
rect 382864 230265 382870 230277
rect 373706 230237 382870 230265
rect 373706 230225 373712 230237
rect 382864 230225 382870 230237
rect 382922 230225 382928 230277
rect 387280 230225 387286 230277
rect 387338 230265 387344 230277
rect 398512 230265 398518 230277
rect 387338 230237 398518 230265
rect 387338 230225 387344 230237
rect 398512 230225 398518 230237
rect 398570 230225 398576 230277
rect 399088 230225 399094 230277
rect 399146 230265 399152 230277
rect 404944 230265 404950 230277
rect 399146 230237 404950 230265
rect 399146 230225 399152 230237
rect 404944 230225 404950 230237
rect 405002 230225 405008 230277
rect 413488 230265 413494 230277
rect 405058 230237 413494 230265
rect 285386 230163 358526 230191
rect 285386 230151 285392 230163
rect 367504 230151 367510 230203
rect 367562 230191 367568 230203
rect 369424 230191 369430 230203
rect 367562 230163 369430 230191
rect 367562 230151 367568 230163
rect 369424 230151 369430 230163
rect 369482 230151 369488 230203
rect 369616 230151 369622 230203
rect 369674 230191 369680 230203
rect 372496 230191 372502 230203
rect 369674 230163 372502 230191
rect 369674 230151 369680 230163
rect 372496 230151 372502 230163
rect 372554 230151 372560 230203
rect 373744 230151 373750 230203
rect 373802 230191 373808 230203
rect 382480 230191 382486 230203
rect 373802 230163 382486 230191
rect 373802 230151 373808 230163
rect 382480 230151 382486 230163
rect 382538 230151 382544 230203
rect 398704 230151 398710 230203
rect 398762 230191 398768 230203
rect 400240 230191 400246 230203
rect 398762 230163 400246 230191
rect 398762 230151 398768 230163
rect 400240 230151 400246 230163
rect 400298 230151 400304 230203
rect 400432 230151 400438 230203
rect 400490 230191 400496 230203
rect 404176 230191 404182 230203
rect 400490 230163 404182 230191
rect 400490 230151 400496 230163
rect 404176 230151 404182 230163
rect 404234 230151 404240 230203
rect 404368 230151 404374 230203
rect 404426 230191 404432 230203
rect 405058 230191 405086 230237
rect 413488 230225 413494 230237
rect 413546 230225 413552 230277
rect 413584 230225 413590 230277
rect 413642 230265 413648 230277
rect 427984 230265 427990 230277
rect 413642 230237 427990 230265
rect 413642 230225 413648 230237
rect 427984 230225 427990 230237
rect 428042 230225 428048 230277
rect 428752 230225 428758 230277
rect 428810 230265 428816 230277
rect 429328 230265 429334 230277
rect 428810 230237 429334 230265
rect 428810 230225 428816 230237
rect 429328 230225 429334 230237
rect 429386 230225 429392 230277
rect 431056 230225 431062 230277
rect 431114 230265 431120 230277
rect 436912 230265 436918 230277
rect 431114 230237 436918 230265
rect 431114 230225 431120 230237
rect 436912 230225 436918 230237
rect 436970 230225 436976 230277
rect 437008 230225 437014 230277
rect 437066 230265 437072 230277
rect 443056 230265 443062 230277
rect 437066 230237 443062 230265
rect 437066 230225 437072 230237
rect 443056 230225 443062 230237
rect 443114 230225 443120 230277
rect 501712 230265 501718 230277
rect 443170 230237 501718 230265
rect 404426 230163 405086 230191
rect 404426 230151 404432 230163
rect 405232 230151 405238 230203
rect 405290 230191 405296 230203
rect 419152 230191 419158 230203
rect 405290 230163 419158 230191
rect 405290 230151 405296 230163
rect 419152 230151 419158 230163
rect 419210 230151 419216 230203
rect 425584 230151 425590 230203
rect 425642 230191 425648 230203
rect 439120 230191 439126 230203
rect 425642 230163 439126 230191
rect 425642 230151 425648 230163
rect 439120 230151 439126 230163
rect 439178 230151 439184 230203
rect 439234 230163 439838 230191
rect 161200 230077 161206 230129
rect 161258 230117 161264 230129
rect 212080 230117 212086 230129
rect 161258 230089 212086 230117
rect 161258 230077 161264 230089
rect 212080 230077 212086 230089
rect 212138 230077 212144 230129
rect 352336 230077 352342 230129
rect 352394 230117 352400 230129
rect 352394 230089 433214 230117
rect 352394 230077 352400 230089
rect 152560 230003 152566 230055
rect 152618 230043 152624 230055
rect 211696 230043 211702 230055
rect 152618 230015 211702 230043
rect 152618 230003 152624 230015
rect 211696 230003 211702 230015
rect 211754 230003 211760 230055
rect 351952 230003 351958 230055
rect 352010 230043 352016 230055
rect 352010 230015 433118 230043
rect 352010 230003 352016 230015
rect 146512 229929 146518 229981
rect 146570 229969 146576 229981
rect 211024 229969 211030 229981
rect 146570 229941 211030 229969
rect 146570 229929 146576 229941
rect 211024 229929 211030 229941
rect 211082 229929 211088 229981
rect 350128 229929 350134 229981
rect 350186 229969 350192 229981
rect 350186 229941 433022 229969
rect 350186 229929 350192 229941
rect 140752 229855 140758 229907
rect 140810 229895 140816 229907
rect 209488 229895 209494 229907
rect 140810 229867 209494 229895
rect 140810 229855 140816 229867
rect 209488 229855 209494 229867
rect 209546 229855 209552 229907
rect 349744 229855 349750 229907
rect 349802 229895 349808 229907
rect 349802 229867 432926 229895
rect 349802 229855 349808 229867
rect 140656 229781 140662 229833
rect 140714 229821 140720 229833
rect 209872 229821 209878 229833
rect 140714 229793 209878 229821
rect 140714 229781 140720 229793
rect 209872 229781 209878 229793
rect 209930 229781 209936 229833
rect 348976 229781 348982 229833
rect 349034 229821 349040 229833
rect 349034 229793 432830 229821
rect 349034 229781 349040 229793
rect 140944 229707 140950 229759
rect 141002 229747 141008 229759
rect 208816 229747 208822 229759
rect 141002 229719 208822 229747
rect 141002 229707 141008 229719
rect 208816 229707 208822 229719
rect 208874 229707 208880 229759
rect 348688 229707 348694 229759
rect 348746 229747 348752 229759
rect 348746 229719 432734 229747
rect 348746 229707 348752 229719
rect 140464 229633 140470 229685
rect 140522 229673 140528 229685
rect 209104 229673 209110 229685
rect 140522 229645 209110 229673
rect 140522 229633 140528 229645
rect 209104 229633 209110 229645
rect 209162 229633 209168 229685
rect 348304 229633 348310 229685
rect 348362 229673 348368 229685
rect 432592 229673 432598 229685
rect 348362 229645 432598 229673
rect 348362 229633 348368 229645
rect 432592 229633 432598 229645
rect 432650 229633 432656 229685
rect 210640 229599 210646 229611
rect 141058 229571 210646 229599
rect 140368 229485 140374 229537
rect 140426 229525 140432 229537
rect 141058 229525 141086 229571
rect 210640 229559 210646 229571
rect 210698 229559 210704 229611
rect 347920 229559 347926 229611
rect 347978 229599 347984 229611
rect 368080 229599 368086 229611
rect 347978 229571 368086 229599
rect 347978 229559 347984 229571
rect 368080 229559 368086 229571
rect 368138 229559 368144 229611
rect 368176 229559 368182 229611
rect 368234 229599 368240 229611
rect 373264 229599 373270 229611
rect 368234 229571 373270 229599
rect 368234 229559 368240 229571
rect 373264 229559 373270 229571
rect 373322 229559 373328 229611
rect 373360 229559 373366 229611
rect 373418 229599 373424 229611
rect 432400 229599 432406 229611
rect 373418 229571 432406 229599
rect 373418 229559 373424 229571
rect 432400 229559 432406 229571
rect 432458 229559 432464 229611
rect 140426 229497 141086 229525
rect 140426 229485 140432 229497
rect 141136 229485 141142 229537
rect 141194 229525 141200 229537
rect 210256 229525 210262 229537
rect 141194 229497 210262 229525
rect 141194 229485 141200 229497
rect 210256 229485 210262 229497
rect 210314 229485 210320 229537
rect 350512 229485 350518 229537
rect 350570 229525 350576 229537
rect 354064 229525 354070 229537
rect 350570 229497 354070 229525
rect 350570 229485 350576 229497
rect 354064 229485 354070 229497
rect 354122 229485 354128 229537
rect 354160 229485 354166 229537
rect 354218 229525 354224 229537
rect 358384 229525 358390 229537
rect 354218 229497 358390 229525
rect 354218 229485 354224 229497
rect 358384 229485 358390 229497
rect 358442 229485 358448 229537
rect 358480 229485 358486 229537
rect 358538 229525 358544 229537
rect 432304 229525 432310 229537
rect 358538 229497 432310 229525
rect 358538 229485 358544 229497
rect 432304 229485 432310 229497
rect 432362 229485 432368 229537
rect 432706 229525 432734 229719
rect 432802 229599 432830 229793
rect 432898 229673 432926 229867
rect 432994 229821 433022 229941
rect 433090 229895 433118 230015
rect 433186 229969 433214 230089
rect 434800 230077 434806 230129
rect 434858 230117 434864 230129
rect 439234 230117 439262 230163
rect 434858 230089 439262 230117
rect 439810 230117 439838 230163
rect 440176 230151 440182 230203
rect 440234 230191 440240 230203
rect 443170 230191 443198 230237
rect 501712 230225 501718 230237
rect 501770 230225 501776 230277
rect 483856 230191 483862 230203
rect 440234 230163 443198 230191
rect 453538 230163 483862 230191
rect 440234 230151 440240 230163
rect 453538 230117 453566 230163
rect 483856 230151 483862 230163
rect 483914 230151 483920 230203
rect 495184 230151 495190 230203
rect 495242 230191 495248 230203
rect 505360 230191 505366 230203
rect 495242 230163 505366 230191
rect 495242 230151 495248 230163
rect 505360 230151 505366 230163
rect 505418 230151 505424 230203
rect 439810 230089 453566 230117
rect 434858 230077 434864 230089
rect 454672 230077 454678 230129
rect 454730 230117 454736 230129
rect 501328 230117 501334 230129
rect 454730 230089 501334 230117
rect 454730 230077 454736 230089
rect 501328 230077 501334 230089
rect 501386 230077 501392 230129
rect 439792 230003 439798 230055
rect 439850 230043 439856 230055
rect 507568 230043 507574 230055
rect 439850 230015 507574 230043
rect 439850 230003 439856 230015
rect 507568 230003 507574 230015
rect 507626 230003 507632 230055
rect 438832 229969 438838 229981
rect 433186 229941 438838 229969
rect 438832 229929 438838 229941
rect 438890 229929 438896 229981
rect 439024 229929 439030 229981
rect 439082 229969 439088 229981
rect 447856 229969 447862 229981
rect 439082 229941 447862 229969
rect 439082 229929 439088 229941
rect 447856 229929 447862 229941
rect 447914 229929 447920 229981
rect 452080 229929 452086 229981
rect 452138 229969 452144 229981
rect 480400 229969 480406 229981
rect 452138 229941 480406 229969
rect 452138 229929 452144 229941
rect 480400 229929 480406 229941
rect 480458 229929 480464 229981
rect 494416 229929 494422 229981
rect 494474 229969 494480 229981
rect 507184 229969 507190 229981
rect 494474 229941 507190 229969
rect 494474 229929 494480 229941
rect 507184 229929 507190 229941
rect 507242 229929 507248 229981
rect 439888 229895 439894 229907
rect 433090 229867 439894 229895
rect 439888 229855 439894 229867
rect 439946 229855 439952 229907
rect 439984 229855 439990 229907
rect 440042 229895 440048 229907
rect 445936 229895 445942 229907
rect 440042 229867 445942 229895
rect 440042 229855 440048 229867
rect 445936 229855 445942 229867
rect 445994 229855 446000 229907
rect 446416 229855 446422 229907
rect 446474 229895 446480 229907
rect 502768 229895 502774 229907
rect 446474 229867 502774 229895
rect 446474 229855 446480 229867
rect 502768 229855 502774 229867
rect 502826 229855 502832 229907
rect 443632 229821 443638 229833
rect 432994 229793 443638 229821
rect 443632 229781 443638 229793
rect 443690 229781 443696 229833
rect 443842 229793 445502 229821
rect 436048 229707 436054 229759
rect 436106 229747 436112 229759
rect 443842 229747 443870 229793
rect 436106 229719 443870 229747
rect 445474 229747 445502 229793
rect 445552 229781 445558 229833
rect 445610 229821 445616 229833
rect 510544 229821 510550 229833
rect 445610 229793 510550 229821
rect 445610 229781 445616 229793
rect 510544 229781 510550 229793
rect 510602 229781 510608 229833
rect 448336 229747 448342 229759
rect 445474 229719 448342 229747
rect 436106 229707 436112 229719
rect 448336 229707 448342 229719
rect 448394 229707 448400 229759
rect 453616 229707 453622 229759
rect 453674 229747 453680 229759
rect 504688 229747 504694 229759
rect 453674 229719 504694 229747
rect 453674 229707 453680 229719
rect 504688 229707 504694 229719
rect 504746 229707 504752 229759
rect 444496 229673 444502 229685
rect 432898 229645 444502 229673
rect 444496 229633 444502 229645
rect 444554 229633 444560 229685
rect 447472 229633 447478 229685
rect 447530 229673 447536 229685
rect 459280 229673 459286 229685
rect 447530 229645 459286 229673
rect 447530 229633 447536 229645
rect 459280 229633 459286 229645
rect 459338 229633 459344 229685
rect 501136 229633 501142 229685
rect 501194 229673 501200 229685
rect 514576 229673 514582 229685
rect 501194 229645 514582 229673
rect 501194 229633 501200 229645
rect 514576 229633 514582 229645
rect 514634 229633 514640 229685
rect 445840 229599 445846 229611
rect 432802 229571 445846 229599
rect 445840 229559 445846 229571
rect 445898 229559 445904 229611
rect 445936 229559 445942 229611
rect 445994 229599 446000 229611
rect 445994 229571 447518 229599
rect 445994 229559 446000 229571
rect 447490 229537 447518 229571
rect 447664 229559 447670 229611
rect 447722 229599 447728 229611
rect 511600 229599 511606 229611
rect 447722 229571 511606 229599
rect 447722 229559 447728 229571
rect 511600 229559 511606 229571
rect 511658 229559 511664 229611
rect 633808 229559 633814 229611
rect 633866 229599 633872 229611
rect 649840 229599 649846 229611
rect 633866 229571 649846 229599
rect 633866 229559 633872 229571
rect 649840 229559 649846 229571
rect 649898 229559 649904 229611
rect 446896 229525 446902 229537
rect 432706 229497 446902 229525
rect 446896 229485 446902 229497
rect 446954 229485 446960 229537
rect 447472 229485 447478 229537
rect 447530 229485 447536 229537
rect 449104 229485 449110 229537
rect 449162 229525 449168 229537
rect 512368 229525 512374 229537
rect 449162 229497 512374 229525
rect 449162 229485 449168 229497
rect 512368 229485 512374 229497
rect 512426 229485 512432 229537
rect 633136 229485 633142 229537
rect 633194 229525 633200 229537
rect 649552 229525 649558 229537
rect 633194 229497 649558 229525
rect 633194 229485 633200 229497
rect 649552 229485 649558 229497
rect 649610 229485 649616 229537
rect 663952 229485 663958 229537
rect 664010 229525 664016 229537
rect 674416 229525 674422 229537
rect 664010 229497 674422 229525
rect 664010 229485 664016 229497
rect 674416 229485 674422 229497
rect 674474 229485 674480 229537
rect 139984 229411 139990 229463
rect 140042 229411 140048 229463
rect 140560 229411 140566 229463
rect 140618 229451 140624 229463
rect 215056 229451 215062 229463
rect 140618 229423 215062 229451
rect 140618 229411 140624 229423
rect 215056 229411 215062 229423
rect 215114 229411 215120 229463
rect 282832 229411 282838 229463
rect 282890 229451 282896 229463
rect 370192 229451 370198 229463
rect 282890 229423 370198 229451
rect 282890 229411 282896 229423
rect 370192 229411 370198 229423
rect 370250 229411 370256 229463
rect 370384 229411 370390 229463
rect 370442 229451 370448 229463
rect 374032 229451 374038 229463
rect 370442 229423 374038 229451
rect 370442 229411 370448 229423
rect 374032 229411 374038 229423
rect 374090 229411 374096 229463
rect 375184 229411 375190 229463
rect 375242 229451 375248 229463
rect 382768 229451 382774 229463
rect 375242 229423 382774 229451
rect 375242 229411 375248 229423
rect 382768 229411 382774 229423
rect 382826 229411 382832 229463
rect 398320 229411 398326 229463
rect 398378 229451 398384 229463
rect 405328 229451 405334 229463
rect 398378 229423 405334 229451
rect 398378 229411 398384 229423
rect 405328 229411 405334 229423
rect 405386 229411 405392 229463
rect 406384 229411 406390 229463
rect 406442 229451 406448 229463
rect 413008 229451 413014 229463
rect 406442 229423 413014 229451
rect 406442 229411 406448 229423
rect 413008 229411 413014 229423
rect 413066 229411 413072 229463
rect 413104 229411 413110 229463
rect 413162 229451 413168 229463
rect 427600 229451 427606 229463
rect 413162 229423 427606 229451
rect 413162 229411 413168 229423
rect 427600 229411 427606 229423
rect 427658 229411 427664 229463
rect 428176 229411 428182 229463
rect 428234 229451 428240 229463
rect 433072 229451 433078 229463
rect 428234 229423 433078 229451
rect 428234 229411 428240 229423
rect 433072 229411 433078 229423
rect 433130 229411 433136 229463
rect 433648 229411 433654 229463
rect 433706 229451 433712 229463
rect 479440 229451 479446 229463
rect 433706 229423 479446 229451
rect 433706 229411 433712 229423
rect 479440 229411 479446 229423
rect 479498 229411 479504 229463
rect 494800 229411 494806 229463
rect 494858 229451 494864 229463
rect 507952 229451 507958 229463
rect 494858 229423 507958 229451
rect 494858 229411 494864 229423
rect 507952 229411 507958 229423
rect 508010 229411 508016 229463
rect 632752 229411 632758 229463
rect 632810 229451 632816 229463
rect 649456 229451 649462 229463
rect 632810 229423 649462 229451
rect 632810 229411 632816 229423
rect 649456 229411 649462 229423
rect 649514 229411 649520 229463
rect 140002 229377 140030 229411
rect 211312 229377 211318 229389
rect 140002 229349 211318 229377
rect 211312 229337 211318 229349
rect 211370 229337 211376 229389
rect 347152 229337 347158 229389
rect 347210 229377 347216 229389
rect 449488 229377 449494 229389
rect 347210 229349 449494 229377
rect 347210 229337 347216 229349
rect 449488 229337 449494 229349
rect 449546 229337 449552 229389
rect 451984 229337 451990 229389
rect 452042 229377 452048 229389
rect 513808 229377 513814 229389
rect 452042 229349 513814 229377
rect 452042 229337 452048 229349
rect 513808 229337 513814 229349
rect 513866 229337 513872 229389
rect 632368 229337 632374 229389
rect 632426 229377 632432 229389
rect 650416 229377 650422 229389
rect 632426 229349 650422 229377
rect 632426 229337 632432 229349
rect 650416 229337 650422 229349
rect 650474 229337 650480 229389
rect 141232 229263 141238 229315
rect 141290 229303 141296 229315
rect 213904 229303 213910 229315
rect 141290 229275 213910 229303
rect 141290 229263 141296 229275
rect 213904 229263 213910 229275
rect 213962 229263 213968 229315
rect 347536 229263 347542 229315
rect 347594 229303 347600 229315
rect 358480 229303 358486 229315
rect 347594 229275 358486 229303
rect 347594 229263 347600 229275
rect 358480 229263 358486 229275
rect 358538 229263 358544 229315
rect 358576 229263 358582 229315
rect 358634 229303 358640 229315
rect 367888 229303 367894 229315
rect 358634 229275 367894 229303
rect 358634 229263 358640 229275
rect 367888 229263 367894 229275
rect 367946 229263 367952 229315
rect 417616 229303 417622 229315
rect 369346 229275 417622 229303
rect 139984 229189 139990 229241
rect 140042 229189 140048 229241
rect 141424 229189 141430 229241
rect 141482 229229 141488 229241
rect 214672 229229 214678 229241
rect 141482 229201 214678 229229
rect 141482 229189 141488 229201
rect 214672 229189 214678 229201
rect 214730 229189 214736 229241
rect 284176 229189 284182 229241
rect 284234 229229 284240 229241
rect 356272 229229 356278 229241
rect 284234 229201 356278 229229
rect 284234 229189 284240 229201
rect 356272 229189 356278 229201
rect 356330 229189 356336 229241
rect 366640 229229 366646 229241
rect 356386 229201 366646 229229
rect 140002 229155 140030 229189
rect 215440 229155 215446 229167
rect 140002 229127 215446 229155
rect 215440 229115 215446 229127
rect 215498 229115 215504 229167
rect 282928 229115 282934 229167
rect 282986 229155 282992 229167
rect 356386 229155 356414 229201
rect 366640 229189 366646 229201
rect 366698 229189 366704 229241
rect 358192 229155 358198 229167
rect 282986 229127 356414 229155
rect 357634 229127 358198 229155
rect 282986 229115 282992 229127
rect 144304 229041 144310 229093
rect 144362 229081 144368 229093
rect 215728 229081 215734 229093
rect 144362 229053 215734 229081
rect 144362 229041 144368 229053
rect 215728 229041 215734 229053
rect 215786 229041 215792 229093
rect 282256 229041 282262 229093
rect 282314 229081 282320 229093
rect 357634 229081 357662 229127
rect 358192 229115 358198 229127
rect 358250 229115 358256 229167
rect 358768 229115 358774 229167
rect 358826 229155 358832 229167
rect 368176 229155 368182 229167
rect 358826 229127 368182 229155
rect 358826 229115 358832 229127
rect 368176 229115 368182 229127
rect 368234 229115 368240 229167
rect 369346 229081 369374 229275
rect 417616 229263 417622 229275
rect 417674 229263 417680 229315
rect 456112 229263 456118 229315
rect 456170 229303 456176 229315
rect 463024 229303 463030 229315
rect 456170 229275 463030 229303
rect 456170 229263 456176 229275
rect 463024 229263 463030 229275
rect 463082 229263 463088 229315
rect 463120 229263 463126 229315
rect 463178 229303 463184 229315
rect 513136 229303 513142 229315
rect 463178 229275 513142 229303
rect 463178 229263 463184 229275
rect 513136 229263 513142 229275
rect 513194 229263 513200 229315
rect 631984 229263 631990 229315
rect 632042 229303 632048 229315
rect 650224 229303 650230 229315
rect 632042 229275 650230 229303
rect 632042 229263 632048 229275
rect 650224 229263 650230 229275
rect 650282 229263 650288 229315
rect 369424 229189 369430 229241
rect 369482 229229 369488 229241
rect 373648 229229 373654 229241
rect 369482 229201 373654 229229
rect 369482 229189 369488 229201
rect 373648 229189 373654 229201
rect 373706 229189 373712 229241
rect 376720 229189 376726 229241
rect 376778 229229 376784 229241
rect 376778 229201 382718 229229
rect 376778 229189 376784 229201
rect 370288 229115 370294 229167
rect 370346 229155 370352 229167
rect 381040 229155 381046 229167
rect 370346 229127 381046 229155
rect 370346 229115 370352 229127
rect 381040 229115 381046 229127
rect 381098 229115 381104 229167
rect 282314 229053 357662 229081
rect 357730 229053 369374 229081
rect 282314 229041 282320 229053
rect 148720 228967 148726 229019
rect 148778 229007 148784 229019
rect 288688 229007 288694 229019
rect 148778 228979 288694 229007
rect 148778 228967 148784 228979
rect 288688 228967 288694 228979
rect 288746 229007 288752 229019
rect 318832 229007 318838 229019
rect 288746 228979 318838 229007
rect 288746 228967 288752 228979
rect 318832 228967 318838 228979
rect 318890 228967 318896 229019
rect 346480 228967 346486 229019
rect 346538 229007 346544 229019
rect 357730 229007 357758 229053
rect 372688 229041 372694 229093
rect 372746 229081 372752 229093
rect 381712 229081 381718 229093
rect 372746 229053 381718 229081
rect 372746 229041 372752 229053
rect 381712 229041 381718 229053
rect 381770 229041 381776 229093
rect 382690 229081 382718 229201
rect 382768 229189 382774 229241
rect 382826 229229 382832 229241
rect 382826 229201 477662 229229
rect 382826 229189 382832 229201
rect 382864 229115 382870 229167
rect 382922 229155 382928 229167
rect 477520 229155 477526 229167
rect 382922 229127 477526 229155
rect 382922 229115 382928 229127
rect 477520 229115 477526 229127
rect 477578 229115 477584 229167
rect 477634 229155 477662 229201
rect 479440 229189 479446 229241
rect 479498 229229 479504 229241
rect 502096 229229 502102 229241
rect 479498 229201 502102 229229
rect 479498 229189 479504 229201
rect 502096 229189 502102 229201
rect 502154 229189 502160 229241
rect 631600 229189 631606 229241
rect 631658 229229 631664 229241
rect 650128 229229 650134 229241
rect 631658 229201 650134 229229
rect 631658 229189 631664 229201
rect 650128 229189 650134 229201
rect 650186 229189 650192 229241
rect 489904 229155 489910 229167
rect 477634 229127 489910 229155
rect 489904 229115 489910 229127
rect 489962 229115 489968 229167
rect 493552 229115 493558 229167
rect 493610 229155 493616 229167
rect 508720 229155 508726 229167
rect 493610 229127 508726 229155
rect 493610 229115 493616 229127
rect 508720 229115 508726 229127
rect 508778 229115 508784 229167
rect 631312 229115 631318 229167
rect 631370 229155 631376 229167
rect 649936 229155 649942 229167
rect 631370 229127 649942 229155
rect 631370 229115 631376 229127
rect 649936 229115 649942 229127
rect 649994 229115 650000 229167
rect 491440 229081 491446 229093
rect 382690 229053 491446 229081
rect 491440 229041 491446 229053
rect 491498 229041 491504 229093
rect 493936 229041 493942 229093
rect 493994 229081 494000 229093
rect 510928 229081 510934 229093
rect 493994 229053 510934 229081
rect 493994 229041 494000 229053
rect 510928 229041 510934 229053
rect 510986 229041 510992 229093
rect 633520 229041 633526 229093
rect 633578 229081 633584 229093
rect 649744 229081 649750 229093
rect 633578 229053 649750 229081
rect 633578 229041 633584 229053
rect 649744 229041 649750 229053
rect 649802 229041 649808 229093
rect 346538 228979 357758 229007
rect 346538 228967 346544 228979
rect 357808 228967 357814 229019
rect 357866 229007 357872 229019
rect 367792 229007 367798 229019
rect 357866 228979 367798 229007
rect 357866 228967 357872 228979
rect 367792 228967 367798 228979
rect 367850 228967 367856 229019
rect 367888 228967 367894 229019
rect 367946 229007 367952 229019
rect 380272 229007 380278 229019
rect 367946 228979 380278 229007
rect 367946 228967 367952 228979
rect 380272 228967 380278 228979
rect 380330 228967 380336 229019
rect 380560 228967 380566 229019
rect 380618 229007 380624 229019
rect 380618 228979 477470 229007
rect 380618 228967 380624 228979
rect 169840 228893 169846 228945
rect 169898 228933 169904 228945
rect 212848 228933 212854 228945
rect 169898 228905 212854 228933
rect 169898 228893 169904 228905
rect 212848 228893 212854 228905
rect 212906 228893 212912 228945
rect 284080 228893 284086 228945
rect 284138 228933 284144 228945
rect 350320 228933 350326 228945
rect 284138 228905 350326 228933
rect 284138 228893 284144 228905
rect 350320 228893 350326 228905
rect 350378 228893 350384 228945
rect 368464 228933 368470 228945
rect 350434 228905 368470 228933
rect 178480 228819 178486 228871
rect 178538 228859 178544 228871
rect 213232 228859 213238 228871
rect 178538 228831 213238 228859
rect 178538 228819 178544 228831
rect 213232 228819 213238 228831
rect 213290 228819 213296 228871
rect 286288 228819 286294 228871
rect 286346 228859 286352 228871
rect 350434 228859 350462 228905
rect 368464 228893 368470 228905
rect 368522 228893 368528 228945
rect 370192 228893 370198 228945
rect 370250 228933 370256 228945
rect 397456 228933 397462 228945
rect 370250 228905 380798 228933
rect 370250 228893 370256 228905
rect 286346 228831 350462 228859
rect 286346 228819 286352 228831
rect 350512 228819 350518 228871
rect 350570 228859 350576 228871
rect 350570 228831 366398 228859
rect 350570 228819 350576 228831
rect 184240 228745 184246 228797
rect 184298 228785 184304 228797
rect 213520 228785 213526 228797
rect 184298 228757 213526 228785
rect 184298 228745 184304 228757
rect 213520 228745 213526 228757
rect 213578 228745 213584 228797
rect 286480 228745 286486 228797
rect 286538 228785 286544 228797
rect 366256 228785 366262 228797
rect 286538 228757 366262 228785
rect 286538 228745 286544 228757
rect 366256 228745 366262 228757
rect 366314 228745 366320 228797
rect 204592 228671 204598 228723
rect 204650 228711 204656 228723
rect 205840 228711 205846 228723
rect 204650 228683 205846 228711
rect 204650 228671 204656 228683
rect 205840 228671 205846 228683
rect 205898 228671 205904 228723
rect 214288 228711 214294 228723
rect 205954 228683 214294 228711
rect 192880 228597 192886 228649
rect 192938 228637 192944 228649
rect 205954 228637 205982 228683
rect 214288 228671 214294 228683
rect 214346 228671 214352 228723
rect 285616 228671 285622 228723
rect 285674 228711 285680 228723
rect 365872 228711 365878 228723
rect 285674 228683 365878 228711
rect 285674 228671 285680 228683
rect 365872 228671 365878 228683
rect 365930 228671 365936 228723
rect 366370 228711 366398 228831
rect 366448 228819 366454 228871
rect 366506 228859 366512 228871
rect 380656 228859 380662 228871
rect 366506 228831 380662 228859
rect 366506 228819 366512 228831
rect 380656 228819 380662 228831
rect 380714 228819 380720 228871
rect 367984 228745 367990 228797
rect 368042 228785 368048 228797
rect 374416 228785 374422 228797
rect 368042 228757 374422 228785
rect 368042 228745 368048 228757
rect 374416 228745 374422 228757
rect 374474 228745 374480 228797
rect 376048 228745 376054 228797
rect 376106 228785 376112 228797
rect 380560 228785 380566 228797
rect 376106 228757 380566 228785
rect 376106 228745 376112 228757
rect 380560 228745 380566 228757
rect 380618 228745 380624 228797
rect 366370 228683 368510 228711
rect 192938 228609 205982 228637
rect 192938 228597 192944 228609
rect 349360 228597 349366 228649
rect 349418 228637 349424 228649
rect 360976 228637 360982 228649
rect 349418 228609 360982 228637
rect 349418 228597 349424 228609
rect 360976 228597 360982 228609
rect 361034 228597 361040 228649
rect 361072 228597 361078 228649
rect 361130 228637 361136 228649
rect 368368 228637 368374 228649
rect 361130 228609 368374 228637
rect 361130 228597 361136 228609
rect 368368 228597 368374 228609
rect 368426 228597 368432 228649
rect 368482 228637 368510 228683
rect 370000 228671 370006 228723
rect 370058 228711 370064 228723
rect 374800 228711 374806 228723
rect 370058 228683 374806 228711
rect 370058 228671 370064 228683
rect 374800 228671 374806 228683
rect 374858 228671 374864 228723
rect 380770 228711 380798 228905
rect 394210 228905 397462 228933
rect 384304 228819 384310 228871
rect 384362 228859 384368 228871
rect 394210 228859 394238 228905
rect 397456 228893 397462 228905
rect 397514 228893 397520 228945
rect 397648 228893 397654 228945
rect 397706 228933 397712 228945
rect 405616 228933 405622 228945
rect 397706 228905 405622 228933
rect 397706 228893 397712 228905
rect 405616 228893 405622 228905
rect 405674 228893 405680 228945
rect 410608 228893 410614 228945
rect 410666 228933 410672 228945
rect 414256 228933 414262 228945
rect 410666 228905 414262 228933
rect 410666 228893 410672 228905
rect 414256 228893 414262 228905
rect 414314 228893 414320 228945
rect 414832 228893 414838 228945
rect 414890 228933 414896 228945
rect 427888 228933 427894 228945
rect 414890 228905 427894 228933
rect 414890 228893 414896 228905
rect 427888 228893 427894 228905
rect 427946 228893 427952 228945
rect 427984 228893 427990 228945
rect 428042 228933 428048 228945
rect 451312 228933 451318 228945
rect 428042 228905 451318 228933
rect 428042 228893 428048 228905
rect 451312 228893 451318 228905
rect 451370 228893 451376 228945
rect 452272 228893 452278 228945
rect 452330 228933 452336 228945
rect 457552 228933 457558 228945
rect 452330 228905 457558 228933
rect 452330 228893 452336 228905
rect 457552 228893 457558 228905
rect 457610 228893 457616 228945
rect 477442 228933 477470 228979
rect 477520 228967 477526 229019
rect 477578 229007 477584 229019
rect 489232 229007 489238 229019
rect 477578 228979 489238 229007
rect 477578 228967 477584 228979
rect 489232 228967 489238 228979
rect 489290 228967 489296 229019
rect 497872 228967 497878 229019
rect 497930 229007 497936 229019
rect 511312 229007 511318 229019
rect 497930 228979 511318 229007
rect 497930 228967 497936 228979
rect 511312 228967 511318 228979
rect 511370 228967 511376 229019
rect 541360 228967 541366 229019
rect 541418 229007 541424 229019
rect 650896 229007 650902 229019
rect 541418 228979 650902 229007
rect 541418 228967 541424 228979
rect 650896 228967 650902 228979
rect 650954 228967 650960 229019
rect 490672 228933 490678 228945
rect 477442 228905 490678 228933
rect 490672 228893 490678 228905
rect 490730 228893 490736 228945
rect 494992 228893 494998 228945
rect 495050 228933 495056 228945
rect 510160 228933 510166 228945
rect 495050 228905 510166 228933
rect 495050 228893 495056 228905
rect 510160 228893 510166 228905
rect 510218 228893 510224 228945
rect 669520 228893 669526 228945
rect 669578 228933 669584 228945
rect 674704 228933 674710 228945
rect 669578 228905 674710 228933
rect 669578 228893 669584 228905
rect 674704 228893 674710 228905
rect 674762 228893 674768 228945
rect 384362 228831 394238 228859
rect 384362 228819 384368 228831
rect 394288 228819 394294 228871
rect 394346 228859 394352 228871
rect 394346 228831 403358 228859
rect 394346 228819 394352 228831
rect 393904 228745 393910 228797
rect 393962 228785 393968 228797
rect 403216 228785 403222 228797
rect 393962 228757 403222 228785
rect 393962 228745 393968 228757
rect 403216 228745 403222 228757
rect 403274 228745 403280 228797
rect 403330 228785 403358 228831
rect 403984 228819 403990 228871
rect 404042 228859 404048 228871
rect 404042 228831 418718 228859
rect 404042 228819 404048 228831
rect 417520 228785 417526 228797
rect 403330 228757 417526 228785
rect 417520 228745 417526 228757
rect 417578 228745 417584 228797
rect 388720 228711 388726 228723
rect 380770 228683 388726 228711
rect 388720 228671 388726 228683
rect 388778 228671 388784 228723
rect 394192 228671 394198 228723
rect 394250 228711 394256 228723
rect 398128 228711 398134 228723
rect 394250 228683 398134 228711
rect 394250 228671 394256 228683
rect 398128 228671 398134 228683
rect 398186 228671 398192 228723
rect 398320 228671 398326 228723
rect 398378 228711 398384 228723
rect 412240 228711 412246 228723
rect 398378 228683 412246 228711
rect 398378 228671 398384 228683
rect 412240 228671 412246 228683
rect 412298 228671 412304 228723
rect 413680 228671 413686 228723
rect 413738 228711 413744 228723
rect 418576 228711 418582 228723
rect 413738 228683 418582 228711
rect 413738 228671 413744 228683
rect 418576 228671 418582 228683
rect 418634 228671 418640 228723
rect 418690 228711 418718 228831
rect 418768 228819 418774 228871
rect 418826 228859 418832 228871
rect 456784 228859 456790 228871
rect 418826 228831 456790 228859
rect 418826 228819 418832 228831
rect 456784 228819 456790 228831
rect 456842 228819 456848 228871
rect 498064 228819 498070 228871
rect 498122 228859 498128 228871
rect 511984 228859 511990 228871
rect 498122 228831 511990 228859
rect 498122 228819 498128 228831
rect 511984 228819 511990 228831
rect 512042 228819 512048 228871
rect 419152 228745 419158 228797
rect 419210 228785 419216 228797
rect 456112 228785 456118 228797
rect 419210 228757 456118 228785
rect 419210 228745 419216 228757
rect 456112 228745 456118 228757
rect 456170 228745 456176 228797
rect 493744 228745 493750 228797
rect 493802 228785 493808 228797
rect 509392 228785 509398 228797
rect 493802 228757 509398 228785
rect 493802 228745 493808 228757
rect 509392 228745 509398 228757
rect 509450 228745 509456 228797
rect 453136 228711 453142 228723
rect 418690 228683 453142 228711
rect 453136 228671 453142 228683
rect 453194 228671 453200 228723
rect 432208 228637 432214 228649
rect 368482 228609 432214 228637
rect 432208 228597 432214 228609
rect 432266 228597 432272 228649
rect 432400 228597 432406 228649
rect 432458 228637 432464 228649
rect 434896 228637 434902 228649
rect 432458 228609 434902 228637
rect 432458 228597 432464 228609
rect 434896 228597 434902 228609
rect 434954 228597 434960 228649
rect 450544 228637 450550 228649
rect 438850 228609 450550 228637
rect 282736 228523 282742 228575
rect 282794 228563 282800 228575
rect 352624 228563 352630 228575
rect 282794 228535 352630 228563
rect 282794 228523 282800 228535
rect 352624 228523 352630 228535
rect 352682 228523 352688 228575
rect 356272 228523 356278 228575
rect 356330 228563 356336 228575
rect 367024 228563 367030 228575
rect 356330 228535 367030 228563
rect 356330 228523 356336 228535
rect 367024 228523 367030 228535
rect 367082 228523 367088 228575
rect 368944 228523 368950 228575
rect 369002 228563 369008 228575
rect 372880 228563 372886 228575
rect 369002 228535 372886 228563
rect 369002 228523 369008 228535
rect 372880 228523 372886 228535
rect 372938 228523 372944 228575
rect 375376 228523 375382 228575
rect 375434 228563 375440 228575
rect 378832 228563 378838 228575
rect 375434 228535 378838 228563
rect 375434 228523 375440 228535
rect 378832 228523 378838 228535
rect 378890 228523 378896 228575
rect 382864 228523 382870 228575
rect 382922 228563 382928 228575
rect 403024 228563 403030 228575
rect 382922 228535 403030 228563
rect 382922 228523 382928 228535
rect 403024 228523 403030 228535
rect 403082 228523 403088 228575
rect 403216 228523 403222 228575
rect 403274 228563 403280 228575
rect 410608 228563 410614 228575
rect 403274 228535 410614 228563
rect 403274 228523 403280 228535
rect 410608 228523 410614 228535
rect 410666 228523 410672 228575
rect 420016 228563 420022 228575
rect 411394 228535 420022 228563
rect 283600 228449 283606 228501
rect 283658 228489 283664 228501
rect 361840 228489 361846 228501
rect 283658 228461 361846 228489
rect 283658 228449 283664 228461
rect 361840 228449 361846 228461
rect 361898 228449 361904 228501
rect 372784 228449 372790 228501
rect 372842 228489 372848 228501
rect 378448 228489 378454 228501
rect 372842 228461 378454 228489
rect 372842 228449 372848 228461
rect 378448 228449 378454 228461
rect 378506 228449 378512 228501
rect 394192 228489 394198 228501
rect 378658 228461 394198 228489
rect 346096 228375 346102 228427
rect 346154 228415 346160 228427
rect 378658 228415 378686 228461
rect 394192 228449 394198 228461
rect 394250 228449 394256 228501
rect 403312 228449 403318 228501
rect 403370 228489 403376 228501
rect 411280 228489 411286 228501
rect 403370 228461 411286 228489
rect 403370 228449 403376 228461
rect 411280 228449 411286 228461
rect 411338 228449 411344 228501
rect 346154 228387 378686 228415
rect 346154 228375 346160 228387
rect 390256 228375 390262 228427
rect 390314 228415 390320 228427
rect 399376 228415 399382 228427
rect 390314 228387 399382 228415
rect 390314 228375 390320 228387
rect 399376 228375 399382 228387
rect 399434 228375 399440 228427
rect 409648 228375 409654 228427
rect 409706 228415 409712 228427
rect 411394 228415 411422 228535
rect 420016 228523 420022 228535
rect 420074 228523 420080 228575
rect 426256 228523 426262 228575
rect 426314 228563 426320 228575
rect 438850 228563 438878 228609
rect 450544 228597 450550 228609
rect 450602 228597 450608 228649
rect 499600 228597 499606 228649
rect 499658 228637 499664 228649
rect 514192 228637 514198 228649
rect 499658 228609 514198 228637
rect 499658 228597 499664 228609
rect 514192 228597 514198 228609
rect 514250 228597 514256 228649
rect 426314 228535 438878 228563
rect 426314 228523 426320 228535
rect 438928 228523 438934 228575
rect 438986 228563 438992 228575
rect 475984 228563 475990 228575
rect 438986 228535 475990 228563
rect 438986 228523 438992 228535
rect 475984 228523 475990 228535
rect 476042 228523 476048 228575
rect 411472 228449 411478 228501
rect 411530 228489 411536 228501
rect 434896 228489 434902 228501
rect 411530 228461 434902 228489
rect 411530 228449 411536 228461
rect 434896 228449 434902 228461
rect 434954 228449 434960 228501
rect 434992 228449 434998 228501
rect 435050 228489 435056 228501
rect 439024 228489 439030 228501
rect 435050 228461 439030 228489
rect 435050 228449 435056 228461
rect 439024 228449 439030 228461
rect 439082 228449 439088 228501
rect 440080 228449 440086 228501
rect 440138 228489 440144 228501
rect 452752 228489 452758 228501
rect 440138 228461 452758 228489
rect 440138 228449 440144 228461
rect 452752 228449 452758 228461
rect 452810 228449 452816 228501
rect 459280 228449 459286 228501
rect 459338 228489 459344 228501
rect 509104 228489 509110 228501
rect 459338 228461 509110 228489
rect 459338 228449 459344 228461
rect 509104 228449 509110 228461
rect 509162 228449 509168 228501
rect 409706 228387 411422 228415
rect 409706 228375 409712 228387
rect 411568 228375 411574 228427
rect 411626 228415 411632 228427
rect 416560 228415 416566 228427
rect 411626 228387 416566 228415
rect 411626 228375 411632 228387
rect 416560 228375 416566 228387
rect 416618 228375 416624 228427
rect 418576 228375 418582 228427
rect 418634 228415 418640 228427
rect 418634 228387 419198 228415
rect 418634 228375 418640 228387
rect 204688 228301 204694 228353
rect 204746 228341 204752 228353
rect 205072 228341 205078 228353
rect 204746 228313 205078 228341
rect 204746 228301 204752 228313
rect 205072 228301 205078 228313
rect 205130 228341 205136 228353
rect 206608 228341 206614 228353
rect 205130 228313 206614 228341
rect 205130 228301 205136 228313
rect 206608 228301 206614 228313
rect 206666 228301 206672 228353
rect 284272 228301 284278 228353
rect 284330 228341 284336 228353
rect 284330 228313 323966 228341
rect 284330 228301 284336 228313
rect 323938 228193 323966 228313
rect 346768 228301 346774 228353
rect 346826 228341 346832 228353
rect 358384 228341 358390 228353
rect 346826 228313 358390 228341
rect 346826 228301 346832 228313
rect 358384 228301 358390 228313
rect 358442 228301 358448 228353
rect 368080 228341 368086 228353
rect 358498 228313 368086 228341
rect 350320 228227 350326 228279
rect 350378 228267 350384 228279
rect 358498 228267 358526 228313
rect 368080 228301 368086 228313
rect 368138 228301 368144 228353
rect 368176 228301 368182 228353
rect 368234 228341 368240 228353
rect 382096 228341 382102 228353
rect 368234 228313 382102 228341
rect 368234 228301 368240 228313
rect 382096 228301 382102 228313
rect 382154 228301 382160 228353
rect 395056 228301 395062 228353
rect 395114 228341 395120 228353
rect 399088 228341 399094 228353
rect 395114 228313 399094 228341
rect 395114 228301 395120 228313
rect 399088 228301 399094 228313
rect 399146 228301 399152 228353
rect 402928 228301 402934 228353
rect 402986 228341 402992 228353
rect 418768 228341 418774 228353
rect 402986 228313 418774 228341
rect 402986 228301 402992 228313
rect 418768 228301 418774 228313
rect 418826 228301 418832 228353
rect 419170 228341 419198 228387
rect 423472 228375 423478 228427
rect 423530 228415 423536 228427
rect 435952 228415 435958 228427
rect 423530 228387 435958 228415
rect 423530 228375 423536 228387
rect 435952 228375 435958 228387
rect 436010 228375 436016 228427
rect 472624 228415 472630 228427
rect 436066 228387 472630 228415
rect 428176 228341 428182 228353
rect 419170 228313 428182 228341
rect 428176 228301 428182 228313
rect 428234 228301 428240 228353
rect 428656 228301 428662 228353
rect 428714 228341 428720 228353
rect 436066 228341 436094 228387
rect 472624 228375 472630 228387
rect 472682 228375 472688 228427
rect 428714 228313 436094 228341
rect 428714 228301 428720 228313
rect 439120 228301 439126 228353
rect 439178 228341 439184 228353
rect 469648 228341 469654 228353
rect 439178 228313 469654 228341
rect 439178 228301 439184 228313
rect 469648 228301 469654 228313
rect 469706 228301 469712 228353
rect 350378 228239 358526 228267
rect 350378 228227 350384 228239
rect 360016 228227 360022 228279
rect 360074 228267 360080 228279
rect 411376 228267 411382 228279
rect 360074 228239 411382 228267
rect 360074 228227 360080 228239
rect 411376 228227 411382 228239
rect 411434 228227 411440 228279
rect 411664 228227 411670 228279
rect 411722 228267 411728 228279
rect 423088 228267 423094 228279
rect 411722 228239 423094 228267
rect 411722 228227 411728 228239
rect 423088 228227 423094 228239
rect 423146 228227 423152 228279
rect 431728 228227 431734 228279
rect 431786 228267 431792 228279
rect 438928 228267 438934 228279
rect 431786 228239 438934 228267
rect 431786 228227 431792 228239
rect 438928 228227 438934 228239
rect 438986 228227 438992 228279
rect 439216 228227 439222 228279
rect 439274 228267 439280 228279
rect 471856 228267 471862 228279
rect 439274 228239 471862 228267
rect 439274 228227 439280 228239
rect 471856 228227 471862 228239
rect 471914 228227 471920 228279
rect 499696 228227 499702 228279
rect 499754 228267 499760 228279
rect 513520 228267 513526 228279
rect 499754 228239 513526 228267
rect 499754 228227 499760 228239
rect 513520 228227 513526 228239
rect 513578 228227 513584 228279
rect 360784 228193 360790 228205
rect 323938 228165 360790 228193
rect 360784 228153 360790 228165
rect 360842 228153 360848 228205
rect 360880 228153 360886 228205
rect 360938 228193 360944 228205
rect 431152 228193 431158 228205
rect 360938 228165 431158 228193
rect 360938 228153 360944 228165
rect 431152 228153 431158 228165
rect 431210 228153 431216 228205
rect 432592 228153 432598 228205
rect 432650 228193 432656 228205
rect 447184 228193 447190 228205
rect 432650 228165 447190 228193
rect 432650 228153 432656 228165
rect 447184 228153 447190 228165
rect 447242 228153 447248 228205
rect 447376 228153 447382 228205
rect 447434 228193 447440 228205
rect 474448 228193 474454 228205
rect 447434 228165 474454 228193
rect 447434 228153 447440 228165
rect 474448 228153 474454 228165
rect 474506 228153 474512 228205
rect 283792 228079 283798 228131
rect 283850 228119 283856 228131
rect 357808 228119 357814 228131
rect 283850 228091 357814 228119
rect 283850 228079 283856 228091
rect 357808 228079 357814 228091
rect 357866 228079 357872 228131
rect 358576 228079 358582 228131
rect 358634 228119 358640 228131
rect 434992 228119 434998 228131
rect 358634 228091 434998 228119
rect 358634 228079 358640 228091
rect 434992 228079 434998 228091
rect 435050 228079 435056 228131
rect 440752 228079 440758 228131
rect 440810 228119 440816 228131
rect 459760 228119 459766 228131
rect 440810 228091 459766 228119
rect 440810 228079 440816 228091
rect 459760 228079 459766 228091
rect 459818 228079 459824 228131
rect 354928 228005 354934 228057
rect 354986 228045 354992 228057
rect 360880 228045 360886 228057
rect 354986 228017 360886 228045
rect 354986 228005 354992 228017
rect 360880 228005 360886 228017
rect 360938 228005 360944 228057
rect 360976 228005 360982 228057
rect 361034 228045 361040 228057
rect 414832 228045 414838 228057
rect 361034 228017 414838 228045
rect 361034 228005 361040 228017
rect 414832 228005 414838 228017
rect 414890 228005 414896 228057
rect 414928 228005 414934 228057
rect 414986 228045 414992 228057
rect 423280 228045 423286 228057
rect 414986 228017 423286 228045
rect 414986 228005 414992 228017
rect 423280 228005 423286 228017
rect 423338 228005 423344 228057
rect 431824 228005 431830 228057
rect 431882 228045 431888 228057
rect 435760 228045 435766 228057
rect 431882 228017 435766 228045
rect 431882 228005 431888 228017
rect 435760 228005 435766 228017
rect 435818 228005 435824 228057
rect 435856 228005 435862 228057
rect 435914 228045 435920 228057
rect 440848 228045 440854 228057
rect 435914 228017 440854 228045
rect 435914 228005 435920 228017
rect 440848 228005 440854 228017
rect 440906 228005 440912 228057
rect 440962 228017 448862 228045
rect 352048 227931 352054 227983
rect 352106 227971 352112 227983
rect 358480 227971 358486 227983
rect 352106 227943 358486 227971
rect 352106 227931 352112 227943
rect 358480 227931 358486 227943
rect 358538 227931 358544 227983
rect 358672 227931 358678 227983
rect 358730 227971 358736 227983
rect 369232 227971 369238 227983
rect 358730 227943 369238 227971
rect 358730 227931 358736 227943
rect 369232 227931 369238 227943
rect 369290 227931 369296 227983
rect 378640 227931 378646 227983
rect 378698 227971 378704 227983
rect 435184 227971 435190 227983
rect 378698 227943 435190 227971
rect 378698 227931 378704 227943
rect 435184 227931 435190 227943
rect 435242 227931 435248 227983
rect 440560 227971 440566 227983
rect 435394 227943 440566 227971
rect 351568 227857 351574 227909
rect 351626 227897 351632 227909
rect 432112 227897 432118 227909
rect 351626 227869 432118 227897
rect 351626 227857 351632 227869
rect 432112 227857 432118 227869
rect 432170 227857 432176 227909
rect 432304 227857 432310 227909
rect 432362 227897 432368 227909
rect 435394 227897 435422 227943
rect 440560 227931 440566 227943
rect 440618 227931 440624 227983
rect 440962 227897 440990 228017
rect 448834 227971 448862 228017
rect 449776 228005 449782 228057
rect 449834 228045 449840 228057
rect 459376 228045 459382 228057
rect 449834 228017 459382 228045
rect 449834 228005 449840 228017
rect 459376 228005 459382 228017
rect 459434 228005 459440 228057
rect 477040 227971 477046 227983
rect 448834 227943 477046 227971
rect 477040 227931 477046 227943
rect 477098 227931 477104 227983
rect 432362 227869 435422 227897
rect 435682 227869 440990 227897
rect 432362 227857 432368 227869
rect 351184 227783 351190 227835
rect 351242 227823 351248 227835
rect 432880 227823 432886 227835
rect 351242 227795 432886 227823
rect 351242 227783 351248 227795
rect 432880 227783 432886 227795
rect 432938 227783 432944 227835
rect 204496 227709 204502 227761
rect 204554 227749 204560 227761
rect 206896 227749 206902 227761
rect 204554 227721 206902 227749
rect 204554 227709 204560 227721
rect 206896 227709 206902 227721
rect 206954 227709 206960 227761
rect 207760 227709 207766 227761
rect 207818 227749 207824 227761
rect 242032 227749 242038 227761
rect 207818 227721 242038 227749
rect 207818 227709 207824 227721
rect 242032 227709 242038 227721
rect 242090 227709 242096 227761
rect 350896 227709 350902 227761
rect 350954 227749 350960 227761
rect 432304 227749 432310 227761
rect 350954 227721 432310 227749
rect 350954 227709 350960 227721
rect 432304 227709 432310 227721
rect 432362 227709 432368 227761
rect 434032 227709 434038 227761
rect 434090 227749 434096 227761
rect 435568 227749 435574 227761
rect 434090 227721 435574 227749
rect 434090 227709 434096 227721
rect 435568 227709 435574 227721
rect 435626 227709 435632 227761
rect 144112 227635 144118 227687
rect 144170 227675 144176 227687
rect 149392 227675 149398 227687
rect 144170 227647 149398 227675
rect 144170 227635 144176 227647
rect 149392 227635 149398 227647
rect 149450 227635 149456 227687
rect 204976 227635 204982 227687
rect 205034 227675 205040 227687
rect 207280 227675 207286 227687
rect 205034 227647 207286 227675
rect 205034 227635 205040 227647
rect 207280 227635 207286 227647
rect 207338 227635 207344 227687
rect 207856 227635 207862 227687
rect 207914 227675 207920 227687
rect 293392 227675 293398 227687
rect 207914 227647 293398 227675
rect 207914 227635 207920 227647
rect 293392 227635 293398 227647
rect 293450 227635 293456 227687
rect 358960 227675 358966 227687
rect 343618 227647 358966 227675
rect 139984 227561 139990 227613
rect 140042 227601 140048 227613
rect 140272 227601 140278 227613
rect 140042 227573 140278 227601
rect 140042 227561 140048 227573
rect 140272 227561 140278 227573
rect 140330 227561 140336 227613
rect 144016 227561 144022 227613
rect 144074 227601 144080 227613
rect 177040 227601 177046 227613
rect 144074 227573 177046 227601
rect 144074 227561 144080 227573
rect 177040 227561 177046 227573
rect 177098 227561 177104 227613
rect 199984 227561 199990 227613
rect 200042 227601 200048 227613
rect 200042 227573 200126 227601
rect 200042 227561 200048 227573
rect 200098 227539 200126 227573
rect 204784 227561 204790 227613
rect 204842 227601 204848 227613
rect 206224 227601 206230 227613
rect 204842 227573 206230 227601
rect 204842 227561 204848 227573
rect 206224 227561 206230 227573
rect 206282 227561 206288 227613
rect 221872 227561 221878 227613
rect 221930 227601 221936 227613
rect 242032 227601 242038 227613
rect 221930 227573 242038 227601
rect 221930 227561 221936 227573
rect 242032 227561 242038 227573
rect 242090 227561 242096 227613
rect 343618 227601 343646 227647
rect 358960 227635 358966 227647
rect 359018 227635 359024 227687
rect 359152 227635 359158 227687
rect 359210 227675 359216 227687
rect 432016 227675 432022 227687
rect 359210 227647 432022 227675
rect 359210 227635 359216 227647
rect 432016 227635 432022 227647
rect 432074 227635 432080 227687
rect 432976 227635 432982 227687
rect 433034 227675 433040 227687
rect 435682 227675 435710 227869
rect 441136 227857 441142 227909
rect 441194 227897 441200 227909
rect 447376 227897 447382 227909
rect 441194 227869 447382 227897
rect 441194 227857 441200 227869
rect 447376 227857 447382 227869
rect 447434 227857 447440 227909
rect 447472 227857 447478 227909
rect 447530 227897 447536 227909
rect 475216 227897 475222 227909
rect 447530 227869 475222 227897
rect 447530 227857 447536 227869
rect 475216 227857 475222 227869
rect 475274 227857 475280 227909
rect 669616 227857 669622 227909
rect 669674 227897 669680 227909
rect 674416 227897 674422 227909
rect 669674 227869 674422 227897
rect 669674 227857 669680 227869
rect 674416 227857 674422 227869
rect 674474 227857 674480 227909
rect 435760 227783 435766 227835
rect 435818 227823 435824 227835
rect 449776 227823 449782 227835
rect 435818 227795 449782 227823
rect 435818 227783 435824 227795
rect 449776 227783 449782 227795
rect 449834 227783 449840 227835
rect 502480 227749 502486 227761
rect 437410 227721 502486 227749
rect 433034 227647 435710 227675
rect 433034 227635 433040 227647
rect 435760 227635 435766 227687
rect 435818 227675 435824 227687
rect 437410 227675 437438 227721
rect 502480 227709 502486 227721
rect 502538 227709 502544 227761
rect 435818 227647 437438 227675
rect 435818 227635 435824 227647
rect 437488 227635 437494 227687
rect 437546 227675 437552 227687
rect 506128 227675 506134 227687
rect 437546 227647 506134 227675
rect 437546 227635 437552 227647
rect 506128 227635 506134 227647
rect 506186 227635 506192 227687
rect 506896 227635 506902 227687
rect 506954 227675 506960 227687
rect 512752 227675 512758 227687
rect 506954 227647 512758 227675
rect 506954 227635 506960 227647
rect 512752 227635 512758 227647
rect 512810 227635 512816 227687
rect 283618 227573 343646 227601
rect 200080 227487 200086 227539
rect 200138 227487 200144 227539
rect 208144 227487 208150 227539
rect 208202 227527 208208 227539
rect 221776 227527 221782 227539
rect 208202 227499 221782 227527
rect 208202 227487 208208 227499
rect 221776 227487 221782 227499
rect 221834 227487 221840 227539
rect 256354 227425 282110 227453
rect 242032 227339 242038 227391
rect 242090 227379 242096 227391
rect 256354 227379 256382 227425
rect 242090 227351 256382 227379
rect 282082 227379 282110 227425
rect 283618 227379 283646 227573
rect 357520 227561 357526 227613
rect 357578 227601 357584 227613
rect 378640 227601 378646 227613
rect 357578 227573 366014 227601
rect 357578 227561 357584 227573
rect 360016 227487 360022 227539
rect 360074 227527 360080 227539
rect 360592 227527 360598 227539
rect 360074 227499 360598 227527
rect 360074 227487 360080 227499
rect 360592 227487 360598 227499
rect 360650 227487 360656 227539
rect 365986 227527 366014 227573
rect 367426 227573 378646 227601
rect 367426 227527 367454 227573
rect 378640 227561 378646 227573
rect 378698 227561 378704 227613
rect 386896 227561 386902 227613
rect 386954 227601 386960 227613
rect 398896 227601 398902 227613
rect 386954 227573 398902 227601
rect 386954 227561 386960 227573
rect 398896 227561 398902 227573
rect 398954 227561 398960 227613
rect 399088 227561 399094 227613
rect 399146 227601 399152 227613
rect 408112 227601 408118 227613
rect 399146 227573 408118 227601
rect 399146 227561 399152 227573
rect 408112 227561 408118 227573
rect 408170 227561 408176 227613
rect 415984 227561 415990 227613
rect 416042 227601 416048 227613
rect 423184 227601 423190 227613
rect 416042 227573 423190 227601
rect 416042 227561 416048 227573
rect 423184 227561 423190 227573
rect 423242 227561 423248 227613
rect 430384 227561 430390 227613
rect 430442 227601 430448 227613
rect 435856 227601 435862 227613
rect 430442 227573 435862 227601
rect 430442 227561 430448 227573
rect 435856 227561 435862 227573
rect 435914 227561 435920 227613
rect 435952 227561 435958 227613
rect 436010 227601 436016 227613
rect 461968 227601 461974 227613
rect 436010 227573 461974 227601
rect 436010 227561 436016 227573
rect 461968 227561 461974 227573
rect 462026 227561 462032 227613
rect 501040 227561 501046 227613
rect 501098 227601 501104 227613
rect 539632 227601 539638 227613
rect 501098 227573 539638 227601
rect 501098 227561 501104 227573
rect 539632 227561 539638 227573
rect 539690 227601 539696 227613
rect 541360 227601 541366 227613
rect 539690 227573 541366 227601
rect 539690 227561 539696 227573
rect 541360 227561 541366 227573
rect 541418 227561 541424 227613
rect 365986 227499 367454 227527
rect 384016 227487 384022 227539
rect 384074 227527 384080 227539
rect 391600 227527 391606 227539
rect 384074 227499 391606 227527
rect 384074 227487 384080 227499
rect 391600 227487 391606 227499
rect 391658 227487 391664 227539
rect 403216 227487 403222 227539
rect 403274 227527 403280 227539
rect 409648 227527 409654 227539
rect 403274 227499 409654 227527
rect 403274 227487 403280 227499
rect 409648 227487 409654 227499
rect 409706 227487 409712 227539
rect 418576 227527 418582 227539
rect 409762 227499 418582 227527
rect 329200 227413 329206 227465
rect 329258 227453 329264 227465
rect 348208 227453 348214 227465
rect 329258 227425 348214 227453
rect 329258 227413 329264 227425
rect 348208 227413 348214 227425
rect 348266 227413 348272 227465
rect 348496 227413 348502 227465
rect 348554 227453 348560 227465
rect 409762 227453 409790 227499
rect 418576 227487 418582 227499
rect 418634 227487 418640 227539
rect 418672 227487 418678 227539
rect 418730 227527 418736 227539
rect 432784 227527 432790 227539
rect 418730 227499 432790 227527
rect 418730 227487 418736 227499
rect 432784 227487 432790 227499
rect 432842 227487 432848 227539
rect 432880 227487 432886 227539
rect 432938 227527 432944 227539
rect 441328 227527 441334 227539
rect 432938 227499 441334 227527
rect 432938 227487 432944 227499
rect 441328 227487 441334 227499
rect 441386 227487 441392 227539
rect 441424 227487 441430 227539
rect 441482 227527 441488 227539
rect 455728 227527 455734 227539
rect 441482 227499 455734 227527
rect 441482 227487 441488 227499
rect 455728 227487 455734 227499
rect 455786 227487 455792 227539
rect 418096 227453 418102 227465
rect 348554 227425 409790 227453
rect 409858 227425 418102 227453
rect 348554 227413 348560 227425
rect 282082 227351 283646 227379
rect 242090 227339 242096 227351
rect 346672 227339 346678 227391
rect 346730 227379 346736 227391
rect 409858 227379 409886 227425
rect 418096 227413 418102 227425
rect 418154 227413 418160 227465
rect 418768 227413 418774 227465
rect 418826 227453 418832 227465
rect 431824 227453 431830 227465
rect 418826 227425 431830 227453
rect 418826 227413 418832 227425
rect 431824 227413 431830 227425
rect 431882 227413 431888 227465
rect 432112 227413 432118 227465
rect 432170 227453 432176 227465
rect 440656 227453 440662 227465
rect 432170 227425 440662 227453
rect 432170 227413 432176 227425
rect 440656 227413 440662 227425
rect 440714 227413 440720 227465
rect 346730 227351 409886 227379
rect 346730 227339 346736 227351
rect 409936 227339 409942 227391
rect 409994 227379 410000 227391
rect 422896 227379 422902 227391
rect 409994 227351 422902 227379
rect 409994 227339 410000 227351
rect 422896 227339 422902 227351
rect 422954 227339 422960 227391
rect 423376 227339 423382 227391
rect 423434 227379 423440 227391
rect 430672 227379 430678 227391
rect 423434 227351 430678 227379
rect 423434 227339 423440 227351
rect 430672 227339 430678 227351
rect 430730 227339 430736 227391
rect 432304 227339 432310 227391
rect 432362 227379 432368 227391
rect 442096 227379 442102 227391
rect 432362 227351 442102 227379
rect 432362 227339 432368 227351
rect 442096 227339 442102 227351
rect 442154 227339 442160 227391
rect 527152 227379 527158 227391
rect 442978 227351 527158 227379
rect 344272 227265 344278 227317
rect 344330 227305 344336 227317
rect 344330 227277 414782 227305
rect 344330 227265 344336 227277
rect 326800 227191 326806 227243
rect 326858 227231 326864 227243
rect 409840 227231 409846 227243
rect 326858 227203 409846 227231
rect 326858 227191 326864 227203
rect 409840 227191 409846 227203
rect 409898 227191 409904 227243
rect 414640 227231 414646 227243
rect 409954 227203 414646 227231
rect 315952 227117 315958 227169
rect 316010 227157 316016 227169
rect 409954 227157 409982 227203
rect 414640 227191 414646 227203
rect 414698 227191 414704 227243
rect 414754 227231 414782 227277
rect 414832 227265 414838 227317
rect 414890 227305 414896 227317
rect 422800 227305 422806 227317
rect 414890 227277 422806 227305
rect 414890 227265 414896 227277
rect 422800 227265 422806 227277
rect 422858 227265 422864 227317
rect 423472 227265 423478 227317
rect 423530 227305 423536 227317
rect 431440 227305 431446 227317
rect 423530 227277 431446 227305
rect 423530 227265 423536 227277
rect 431440 227265 431446 227277
rect 431498 227265 431504 227317
rect 432208 227265 432214 227317
rect 432266 227305 432272 227317
rect 442864 227305 442870 227317
rect 432266 227277 442870 227305
rect 432266 227265 432272 227277
rect 442864 227265 442870 227277
rect 442922 227265 442928 227317
rect 434704 227231 434710 227243
rect 414754 227203 434710 227231
rect 434704 227191 434710 227203
rect 434762 227191 434768 227243
rect 434896 227191 434902 227243
rect 434954 227231 434960 227243
rect 442978 227231 443006 227351
rect 527152 227339 527158 227351
rect 527210 227339 527216 227391
rect 434954 227203 443006 227231
rect 434954 227191 434960 227203
rect 443056 227191 443062 227243
rect 443114 227231 443120 227243
rect 450160 227231 450166 227243
rect 443114 227203 450166 227231
rect 443114 227191 443120 227203
rect 450160 227191 450166 227203
rect 450218 227191 450224 227243
rect 316010 227129 409982 227157
rect 316010 227117 316016 227129
rect 410032 227117 410038 227169
rect 410090 227157 410096 227169
rect 422992 227157 422998 227169
rect 410090 227129 422998 227157
rect 410090 227117 410096 227129
rect 422992 227117 422998 227129
rect 423050 227117 423056 227169
rect 423280 227117 423286 227169
rect 423338 227157 423344 227169
rect 446608 227157 446614 227169
rect 423338 227129 446614 227157
rect 423338 227117 423344 227129
rect 446608 227117 446614 227129
rect 446666 227117 446672 227169
rect 316624 227043 316630 227095
rect 316682 227083 316688 227095
rect 422608 227083 422614 227095
rect 316682 227055 422614 227083
rect 316682 227043 316688 227055
rect 422608 227043 422614 227055
rect 422666 227043 422672 227095
rect 423376 227043 423382 227095
rect 423434 227083 423440 227095
rect 429616 227083 429622 227095
rect 423434 227055 429622 227083
rect 423434 227043 423440 227055
rect 429616 227043 429622 227055
rect 429674 227043 429680 227095
rect 439024 227043 439030 227095
rect 439082 227083 439088 227095
rect 458992 227083 458998 227095
rect 439082 227055 458998 227083
rect 439082 227043 439088 227055
rect 458992 227043 458998 227055
rect 459050 227043 459056 227095
rect 315184 226969 315190 227021
rect 315242 227009 315248 227021
rect 423280 227009 423286 227021
rect 315242 226981 423286 227009
rect 315242 226969 315248 226981
rect 423280 226969 423286 226981
rect 423338 226969 423344 227021
rect 432784 226969 432790 227021
rect 432842 227009 432848 227021
rect 437488 227009 437494 227021
rect 432842 226981 437494 227009
rect 432842 226969 432848 226981
rect 437488 226969 437494 226981
rect 437546 226969 437552 227021
rect 437584 226969 437590 227021
rect 437642 227009 437648 227021
rect 464176 227009 464182 227021
rect 437642 226981 464182 227009
rect 437642 226969 437648 226981
rect 464176 226969 464182 226981
rect 464234 226969 464240 227021
rect 333904 226895 333910 226947
rect 333962 226935 333968 226947
rect 429520 226935 429526 226947
rect 333962 226907 429526 226935
rect 333962 226895 333968 226907
rect 429520 226895 429526 226907
rect 429578 226895 429584 226947
rect 432112 226895 432118 226947
rect 432170 226935 432176 226947
rect 443056 226935 443062 226947
rect 432170 226907 443062 226935
rect 432170 226895 432176 226907
rect 443056 226895 443062 226907
rect 443114 226895 443120 226947
rect 326608 226821 326614 226873
rect 326666 226861 326672 226873
rect 418768 226861 418774 226873
rect 326666 226833 418774 226861
rect 326666 226821 326672 226833
rect 418768 226821 418774 226833
rect 418826 226821 418832 226873
rect 418864 226821 418870 226873
rect 418922 226861 418928 226873
rect 429040 226861 429046 226873
rect 418922 226833 429046 226861
rect 418922 226821 418928 226833
rect 429040 226821 429046 226833
rect 429098 226821 429104 226873
rect 438160 226861 438166 226873
rect 429346 226833 438166 226861
rect 348208 226747 348214 226799
rect 348266 226787 348272 226799
rect 348266 226759 418814 226787
rect 348266 226747 348272 226759
rect 317776 226673 317782 226725
rect 317834 226713 317840 226725
rect 418672 226713 418678 226725
rect 317834 226685 418678 226713
rect 317834 226673 317840 226685
rect 418672 226673 418678 226685
rect 418730 226673 418736 226725
rect 418786 226713 418814 226759
rect 419056 226747 419062 226799
rect 419114 226787 419120 226799
rect 429346 226787 429374 226833
rect 438160 226821 438166 226833
rect 438218 226821 438224 226873
rect 419114 226759 429374 226787
rect 419114 226747 419120 226759
rect 429712 226747 429718 226799
rect 429770 226787 429776 226799
rect 446704 226787 446710 226799
rect 429770 226759 446710 226787
rect 429770 226747 429776 226759
rect 446704 226747 446710 226759
rect 446762 226747 446768 226799
rect 418786 226685 429278 226713
rect 318448 226599 318454 226651
rect 318506 226639 318512 226651
rect 418864 226639 418870 226651
rect 318506 226611 418870 226639
rect 318506 226599 318512 226611
rect 418864 226599 418870 226611
rect 418922 226599 418928 226651
rect 426064 226639 426070 226651
rect 419266 226611 426070 226639
rect 307120 226525 307126 226577
rect 307178 226565 307184 226577
rect 419266 226565 419294 226611
rect 426064 226599 426070 226611
rect 426122 226599 426128 226651
rect 428464 226639 428470 226651
rect 426178 226611 428470 226639
rect 307178 226537 419294 226565
rect 307178 226525 307184 226537
rect 419728 226525 419734 226577
rect 419786 226565 419792 226577
rect 426178 226565 426206 226611
rect 428464 226599 428470 226611
rect 428522 226599 428528 226651
rect 429250 226639 429278 226685
rect 429328 226673 429334 226725
rect 429386 226713 429392 226725
rect 452368 226713 452374 226725
rect 429386 226685 452374 226713
rect 429386 226673 429392 226685
rect 452368 226673 452374 226685
rect 452426 226673 452432 226725
rect 433744 226639 433750 226651
rect 429250 226611 433750 226639
rect 433744 226599 433750 226611
rect 433802 226599 433808 226651
rect 435376 226599 435382 226651
rect 435434 226639 435440 226651
rect 439312 226639 439318 226651
rect 435434 226611 439318 226639
rect 435434 226599 435440 226611
rect 439312 226599 439318 226611
rect 439370 226599 439376 226651
rect 419786 226537 426206 226565
rect 419786 226525 419792 226537
rect 426256 226525 426262 226577
rect 426314 226565 426320 226577
rect 527056 226565 527062 226577
rect 426314 226537 439358 226565
rect 426314 226525 426320 226537
rect 319216 226451 319222 226503
rect 319274 226491 319280 226503
rect 418864 226491 418870 226503
rect 319274 226463 418870 226491
rect 319274 226451 319280 226463
rect 418864 226451 418870 226463
rect 418922 226451 418928 226503
rect 419152 226451 419158 226503
rect 419210 226491 419216 226503
rect 420784 226491 420790 226503
rect 419210 226463 420790 226491
rect 419210 226451 419216 226463
rect 420784 226451 420790 226463
rect 420842 226451 420848 226503
rect 422992 226451 422998 226503
rect 423050 226491 423056 226503
rect 423050 226463 428318 226491
rect 423050 226451 423056 226463
rect 305584 226377 305590 226429
rect 305642 226417 305648 226429
rect 409936 226417 409942 226429
rect 305642 226389 409942 226417
rect 305642 226377 305648 226389
rect 409936 226377 409942 226389
rect 409994 226377 410000 226429
rect 427024 226417 427030 226429
rect 410146 226389 427030 226417
rect 307792 226303 307798 226355
rect 307850 226343 307856 226355
rect 410146 226343 410174 226389
rect 427024 226377 427030 226389
rect 427082 226377 427088 226429
rect 427696 226343 427702 226355
rect 307850 226315 410174 226343
rect 410242 226315 427702 226343
rect 307850 226303 307856 226315
rect 304144 226229 304150 226281
rect 304202 226269 304208 226281
rect 410032 226269 410038 226281
rect 304202 226241 410038 226269
rect 304202 226229 304208 226241
rect 410032 226229 410038 226241
rect 410090 226229 410096 226281
rect 306352 226155 306358 226207
rect 306410 226195 306416 226207
rect 410242 226195 410270 226315
rect 427696 226303 427702 226315
rect 427754 226303 427760 226355
rect 428290 226343 428318 226463
rect 428368 226451 428374 226503
rect 428426 226491 428432 226503
rect 428426 226463 439214 226491
rect 428426 226451 428432 226463
rect 428848 226343 428854 226355
rect 428290 226315 428854 226343
rect 428848 226303 428854 226315
rect 428906 226303 428912 226355
rect 435856 226343 435862 226355
rect 429154 226315 435862 226343
rect 410320 226229 410326 226281
rect 410378 226269 410384 226281
rect 426448 226269 426454 226281
rect 410378 226241 426454 226269
rect 410378 226229 410384 226241
rect 426448 226229 426454 226241
rect 426506 226229 426512 226281
rect 306410 226167 410270 226195
rect 306410 226155 306416 226167
rect 410608 226155 410614 226207
rect 410666 226195 410672 226207
rect 412144 226195 412150 226207
rect 410666 226167 412150 226195
rect 410666 226155 410672 226167
rect 412144 226155 412150 226167
rect 412202 226155 412208 226207
rect 413200 226155 413206 226207
rect 413258 226195 413264 226207
rect 429154 226195 429182 226315
rect 435856 226303 435862 226315
rect 435914 226303 435920 226355
rect 429232 226229 429238 226281
rect 429290 226269 429296 226281
rect 429712 226269 429718 226281
rect 429290 226241 429718 226269
rect 429290 226229 429296 226241
rect 429712 226229 429718 226241
rect 429770 226229 429776 226281
rect 431824 226229 431830 226281
rect 431882 226269 431888 226281
rect 438928 226269 438934 226281
rect 431882 226241 438934 226269
rect 431882 226229 431888 226241
rect 438928 226229 438934 226241
rect 438986 226229 438992 226281
rect 439186 226269 439214 226463
rect 439330 226417 439358 226537
rect 439522 226537 527062 226565
rect 439522 226417 439550 226537
rect 527056 226525 527062 226537
rect 527114 226525 527120 226577
rect 439330 226389 439550 226417
rect 460528 226269 460534 226281
rect 439186 226241 460534 226269
rect 460528 226229 460534 226241
rect 460586 226229 460592 226281
rect 413258 226167 429182 226195
rect 413258 226155 413264 226167
rect 429520 226155 429526 226207
rect 429578 226195 429584 226207
rect 448720 226195 448726 226207
rect 429578 226167 448726 226195
rect 429578 226155 429584 226167
rect 448720 226155 448726 226167
rect 448778 226155 448784 226207
rect 304912 226081 304918 226133
rect 304970 226121 304976 226133
rect 418672 226121 418678 226133
rect 304970 226093 418678 226121
rect 304970 226081 304976 226093
rect 418672 226081 418678 226093
rect 418730 226081 418736 226133
rect 418768 226081 418774 226133
rect 418826 226121 418832 226133
rect 425296 226121 425302 226133
rect 418826 226093 425302 226121
rect 418826 226081 418832 226093
rect 425296 226081 425302 226093
rect 425354 226081 425360 226133
rect 425392 226081 425398 226133
rect 425450 226121 425456 226133
rect 439024 226121 439030 226133
rect 425450 226093 439030 226121
rect 425450 226081 425456 226093
rect 439024 226081 439030 226093
rect 439082 226081 439088 226133
rect 439312 226081 439318 226133
rect 439370 226121 439376 226133
rect 484048 226121 484054 226133
rect 439370 226093 484054 226121
rect 439370 226081 439376 226093
rect 484048 226081 484054 226093
rect 484106 226081 484112 226133
rect 359824 226007 359830 226059
rect 359882 226047 359888 226059
rect 413200 226047 413206 226059
rect 359882 226019 413206 226047
rect 359882 226007 359888 226019
rect 413200 226007 413206 226019
rect 413258 226007 413264 226059
rect 418864 226047 418870 226059
rect 418594 226019 418870 226047
rect 355024 225933 355030 225985
rect 355082 225973 355088 225985
rect 418594 225973 418622 226019
rect 418864 226007 418870 226019
rect 418922 226007 418928 226059
rect 418978 226019 434942 226047
rect 418978 225973 419006 226019
rect 434320 225973 434326 225985
rect 355082 225945 418622 225973
rect 418690 225945 419006 225973
rect 419266 225945 434326 225973
rect 355082 225933 355088 225945
rect 358768 225859 358774 225911
rect 358826 225899 358832 225911
rect 418690 225899 418718 225945
rect 358826 225871 418718 225899
rect 358826 225859 358832 225871
rect 418864 225859 418870 225911
rect 418922 225899 418928 225911
rect 419266 225899 419294 225945
rect 434320 225933 434326 225945
rect 434378 225933 434384 225985
rect 434914 225973 434942 226019
rect 434992 226007 434998 226059
rect 435050 226047 435056 226059
rect 454288 226047 454294 226059
rect 435050 226019 454294 226047
rect 435050 226007 435056 226019
rect 454288 226007 454294 226019
rect 454346 226007 454352 226059
rect 436240 225973 436246 225985
rect 434914 225945 436246 225973
rect 436240 225933 436246 225945
rect 436298 225933 436304 225985
rect 436528 225899 436534 225911
rect 418922 225871 419294 225899
rect 419362 225871 436534 225899
rect 418922 225859 418928 225871
rect 362416 225785 362422 225837
rect 362474 225825 362480 225837
rect 419362 225825 419390 225871
rect 436528 225859 436534 225871
rect 436586 225859 436592 225911
rect 362474 225797 419390 225825
rect 362474 225785 362480 225797
rect 419440 225785 419446 225837
rect 419498 225825 419504 225837
rect 419728 225825 419734 225837
rect 419498 225797 419734 225825
rect 419498 225785 419504 225797
rect 419728 225785 419734 225797
rect 419786 225785 419792 225837
rect 420112 225785 420118 225837
rect 420170 225825 420176 225837
rect 425872 225825 425878 225837
rect 420170 225797 425878 225825
rect 420170 225785 420176 225797
rect 425872 225785 425878 225797
rect 425930 225785 425936 225837
rect 426256 225785 426262 225837
rect 426314 225825 426320 225837
rect 427408 225825 427414 225837
rect 426314 225797 427414 225825
rect 426314 225785 426320 225797
rect 427408 225785 427414 225797
rect 427466 225785 427472 225837
rect 427504 225785 427510 225837
rect 427562 225825 427568 225837
rect 432496 225825 432502 225837
rect 427562 225797 432502 225825
rect 427562 225785 427568 225797
rect 432496 225785 432502 225797
rect 432554 225785 432560 225837
rect 437410 225797 457310 225825
rect 352144 225711 352150 225763
rect 352202 225751 352208 225763
rect 410320 225751 410326 225763
rect 352202 225723 410326 225751
rect 352202 225711 352208 225723
rect 410320 225711 410326 225723
rect 410378 225711 410384 225763
rect 410416 225711 410422 225763
rect 410474 225751 410480 225763
rect 420880 225751 420886 225763
rect 410474 225723 420886 225751
rect 410474 225711 410480 225723
rect 420880 225711 420886 225723
rect 420938 225711 420944 225763
rect 437296 225751 437302 225763
rect 429538 225723 437302 225751
rect 362320 225637 362326 225689
rect 362378 225677 362384 225689
rect 411280 225677 411286 225689
rect 362378 225649 411286 225677
rect 362378 225637 362384 225649
rect 411280 225637 411286 225649
rect 411338 225637 411344 225689
rect 411376 225637 411382 225689
rect 411434 225677 411440 225689
rect 415600 225677 415606 225689
rect 411434 225649 415606 225677
rect 411434 225637 411440 225649
rect 415600 225637 415606 225649
rect 415658 225637 415664 225689
rect 417232 225637 417238 225689
rect 417290 225677 417296 225689
rect 418864 225677 418870 225689
rect 417290 225649 418870 225677
rect 417290 225637 417296 225649
rect 418864 225637 418870 225649
rect 418922 225637 418928 225689
rect 419056 225637 419062 225689
rect 419114 225677 419120 225689
rect 419248 225677 419254 225689
rect 419114 225649 419254 225677
rect 419114 225637 419120 225649
rect 419248 225637 419254 225649
rect 419306 225637 419312 225689
rect 429538 225677 429566 225723
rect 437296 225711 437302 225723
rect 437354 225711 437360 225763
rect 419362 225649 429566 225677
rect 351664 225563 351670 225615
rect 351722 225603 351728 225615
rect 418768 225603 418774 225615
rect 351722 225575 418774 225603
rect 351722 225563 351728 225575
rect 418768 225563 418774 225575
rect 418826 225563 418832 225615
rect 419362 225603 419390 225649
rect 429616 225637 429622 225689
rect 429674 225677 429680 225689
rect 437410 225677 437438 225797
rect 437776 225711 437782 225763
rect 437834 225751 437840 225763
rect 457168 225751 457174 225763
rect 437834 225723 457174 225751
rect 437834 225711 437840 225723
rect 457168 225711 457174 225723
rect 457226 225711 457232 225763
rect 457282 225751 457310 225797
rect 512656 225751 512662 225763
rect 457282 225723 512662 225751
rect 512656 225711 512662 225723
rect 512714 225711 512720 225763
rect 429674 225649 437438 225677
rect 429674 225637 429680 225649
rect 418882 225575 419390 225603
rect 420610 225575 420830 225603
rect 360688 225489 360694 225541
rect 360746 225529 360752 225541
rect 418882 225529 418910 225575
rect 360746 225501 418910 225529
rect 360746 225489 360752 225501
rect 418960 225489 418966 225541
rect 419018 225529 419024 225541
rect 420610 225529 420638 225575
rect 419018 225501 420638 225529
rect 419018 225489 419024 225501
rect 420688 225489 420694 225541
rect 420746 225489 420752 225541
rect 420802 225529 420830 225575
rect 420976 225563 420982 225615
rect 421034 225603 421040 225615
rect 424816 225603 424822 225615
rect 421034 225575 424822 225603
rect 421034 225563 421040 225575
rect 424816 225563 424822 225575
rect 424874 225563 424880 225615
rect 426352 225563 426358 225615
rect 426410 225603 426416 225615
rect 521392 225603 521398 225615
rect 426410 225575 521398 225603
rect 426410 225563 426416 225575
rect 521392 225563 521398 225575
rect 521450 225563 521456 225615
rect 433648 225529 433654 225541
rect 420802 225501 433654 225529
rect 433648 225489 433654 225501
rect 433706 225489 433712 225541
rect 433744 225489 433750 225541
rect 433802 225529 433808 225541
rect 443920 225529 443926 225541
rect 433802 225501 443926 225529
rect 433802 225489 433808 225501
rect 443920 225489 443926 225501
rect 443978 225489 443984 225541
rect 354736 225415 354742 225467
rect 354794 225455 354800 225467
rect 420706 225455 420734 225489
rect 354794 225427 420734 225455
rect 354794 225415 354800 225427
rect 420784 225415 420790 225467
rect 420842 225455 420848 225467
rect 425200 225455 425206 225467
rect 420842 225427 425206 225455
rect 420842 225415 420848 225427
rect 425200 225415 425206 225427
rect 425258 225415 425264 225467
rect 427792 225455 427798 225467
rect 426178 225427 427798 225455
rect 354832 225341 354838 225393
rect 354890 225381 354896 225393
rect 420112 225381 420118 225393
rect 354890 225353 420118 225381
rect 354890 225341 354896 225353
rect 420112 225341 420118 225353
rect 420170 225341 420176 225393
rect 421456 225381 421462 225393
rect 420322 225353 421462 225381
rect 355120 225267 355126 225319
rect 355178 225307 355184 225319
rect 420208 225307 420214 225319
rect 355178 225279 420214 225307
rect 355178 225267 355184 225279
rect 420208 225267 420214 225279
rect 420266 225267 420272 225319
rect 365104 225193 365110 225245
rect 365162 225233 365168 225245
rect 420322 225233 420350 225353
rect 421456 225341 421462 225353
rect 421514 225341 421520 225393
rect 422896 225341 422902 225393
rect 422954 225381 422960 225393
rect 426178 225381 426206 225427
rect 427792 225415 427798 225427
rect 427850 225415 427856 225467
rect 427888 225415 427894 225467
rect 427946 225455 427952 225467
rect 445072 225455 445078 225467
rect 427946 225427 445078 225455
rect 427946 225415 427952 225427
rect 445072 225415 445078 225427
rect 445130 225415 445136 225467
rect 422954 225353 426206 225381
rect 422954 225341 422960 225353
rect 426256 225341 426262 225393
rect 426314 225381 426320 225393
rect 489712 225381 489718 225393
rect 426314 225353 489718 225381
rect 426314 225341 426320 225353
rect 489712 225341 489718 225353
rect 489770 225341 489776 225393
rect 421840 225307 421846 225319
rect 365162 225205 420350 225233
rect 420418 225279 421846 225307
rect 365162 225193 365168 225205
rect 363568 225119 363574 225171
rect 363626 225159 363632 225171
rect 420418 225159 420446 225279
rect 421840 225267 421846 225279
rect 421898 225267 421904 225319
rect 423568 225267 423574 225319
rect 423626 225307 423632 225319
rect 431056 225307 431062 225319
rect 423626 225279 431062 225307
rect 423626 225267 423632 225279
rect 431056 225267 431062 225279
rect 431114 225267 431120 225319
rect 431536 225267 431542 225319
rect 431594 225307 431600 225319
rect 433072 225307 433078 225319
rect 431594 225279 433078 225307
rect 431594 225267 431600 225279
rect 433072 225267 433078 225279
rect 433130 225267 433136 225319
rect 438928 225267 438934 225319
rect 438986 225307 438992 225319
rect 442096 225307 442102 225319
rect 438986 225279 442102 225307
rect 438986 225267 438992 225279
rect 442096 225267 442102 225279
rect 442154 225267 442160 225319
rect 420496 225193 420502 225245
rect 420554 225233 420560 225245
rect 435472 225233 435478 225245
rect 420554 225205 435478 225233
rect 420554 225193 420560 225205
rect 435472 225193 435478 225205
rect 435530 225193 435536 225245
rect 422224 225159 422230 225171
rect 363626 225131 420446 225159
rect 420514 225131 422230 225159
rect 363626 225119 363632 225131
rect 366736 225045 366742 225097
rect 366794 225085 366800 225097
rect 420304 225085 420310 225097
rect 366794 225057 420310 225085
rect 366794 225045 366800 225057
rect 420304 225045 420310 225057
rect 420362 225045 420368 225097
rect 363472 224971 363478 225023
rect 363530 225011 363536 225023
rect 420514 225011 420542 225131
rect 422224 225119 422230 225131
rect 422282 225119 422288 225171
rect 423088 225119 423094 225171
rect 423146 225159 423152 225171
rect 448144 225159 448150 225171
rect 423146 225131 448150 225159
rect 423146 225119 423152 225131
rect 448144 225119 448150 225131
rect 448202 225119 448208 225171
rect 420592 225045 420598 225097
rect 420650 225085 420656 225097
rect 434032 225085 434038 225097
rect 420650 225057 434038 225085
rect 420650 225045 420656 225057
rect 434032 225045 434038 225057
rect 434090 225045 434096 225097
rect 363530 224983 420542 225011
rect 363530 224971 363536 224983
rect 421936 224971 421942 225023
rect 421994 225011 422000 225023
rect 435088 225011 435094 225023
rect 421994 224983 435094 225011
rect 421994 224971 422000 224983
rect 435088 224971 435094 224983
rect 435146 224971 435152 225023
rect 444688 225011 444694 225023
rect 436354 224983 444694 225011
rect 368368 224897 368374 224949
rect 368426 224937 368432 224949
rect 381328 224937 381334 224949
rect 368426 224909 381334 224937
rect 368426 224897 368432 224909
rect 381328 224897 381334 224909
rect 381386 224897 381392 224949
rect 395152 224897 395158 224949
rect 395210 224937 395216 224949
rect 436354 224937 436382 224983
rect 444688 224971 444694 224983
rect 444746 224971 444752 225023
rect 395210 224909 436382 224937
rect 395210 224897 395216 224909
rect 436432 224897 436438 224949
rect 436490 224937 436496 224949
rect 449104 224937 449110 224949
rect 436490 224909 449110 224937
rect 436490 224897 436496 224909
rect 449104 224897 449110 224909
rect 449162 224897 449168 224949
rect 359920 224823 359926 224875
rect 359978 224863 359984 224875
rect 374992 224863 374998 224875
rect 359978 224835 374998 224863
rect 359978 224823 359984 224835
rect 374992 224823 374998 224835
rect 375050 224823 375056 224875
rect 395248 224823 395254 224875
rect 395306 224863 395312 224875
rect 443152 224863 443158 224875
rect 395306 224835 443158 224863
rect 395306 224823 395312 224835
rect 443152 224823 443158 224835
rect 443210 224823 443216 224875
rect 394576 224749 394582 224801
rect 394634 224789 394640 224801
rect 441328 224789 441334 224801
rect 394634 224761 441334 224789
rect 394634 224749 394640 224761
rect 441328 224749 441334 224761
rect 441386 224749 441392 224801
rect 144016 224675 144022 224727
rect 144074 224715 144080 224727
rect 174160 224715 174166 224727
rect 144074 224687 174166 224715
rect 144074 224675 144080 224687
rect 174160 224675 174166 224687
rect 174218 224675 174224 224727
rect 348880 224675 348886 224727
rect 348938 224715 348944 224727
rect 424432 224715 424438 224727
rect 348938 224687 424438 224715
rect 348938 224675 348944 224687
rect 424432 224675 424438 224687
rect 424490 224675 424496 224727
rect 424546 224687 425726 224715
rect 395824 224601 395830 224653
rect 395882 224641 395888 224653
rect 405712 224641 405718 224653
rect 395882 224613 405718 224641
rect 395882 224601 395888 224613
rect 405712 224601 405718 224613
rect 405770 224601 405776 224653
rect 417712 224601 417718 224653
rect 417770 224641 417776 224653
rect 418000 224641 418006 224653
rect 417770 224613 418006 224641
rect 417770 224601 417776 224613
rect 418000 224601 418006 224613
rect 418058 224601 418064 224653
rect 418096 224601 418102 224653
rect 418154 224641 418160 224653
rect 424048 224641 424054 224653
rect 418154 224613 424054 224641
rect 418154 224601 418160 224613
rect 424048 224601 424054 224613
rect 424106 224601 424112 224653
rect 424546 224641 424574 224687
rect 424450 224613 424574 224641
rect 374992 224527 374998 224579
rect 375050 224567 375056 224579
rect 420784 224567 420790 224579
rect 375050 224539 420790 224567
rect 375050 224527 375056 224539
rect 420784 224527 420790 224539
rect 420842 224527 420848 224579
rect 420880 224527 420886 224579
rect 420938 224567 420944 224579
rect 424450 224567 424478 224613
rect 420938 224539 424478 224567
rect 425698 224567 425726 224687
rect 425776 224675 425782 224727
rect 425834 224715 425840 224727
rect 426544 224715 426550 224727
rect 425834 224687 426550 224715
rect 425834 224675 425840 224687
rect 426544 224675 426550 224687
rect 426602 224675 426608 224727
rect 432112 224715 432118 224727
rect 426658 224687 432118 224715
rect 426160 224601 426166 224653
rect 426218 224641 426224 224653
rect 426658 224641 426686 224687
rect 432112 224675 432118 224687
rect 432170 224675 432176 224727
rect 432592 224675 432598 224727
rect 432650 224715 432656 224727
rect 452464 224715 452470 224727
rect 432650 224687 452470 224715
rect 432650 224675 432656 224687
rect 452464 224675 452470 224687
rect 452522 224675 452528 224727
rect 426218 224613 426686 224641
rect 426218 224601 426224 224613
rect 430384 224601 430390 224653
rect 430442 224641 430448 224653
rect 433456 224641 433462 224653
rect 430442 224613 433462 224641
rect 430442 224601 430448 224613
rect 433456 224601 433462 224613
rect 433514 224601 433520 224653
rect 426640 224567 426646 224579
rect 425698 224539 426646 224567
rect 420938 224527 420944 224539
rect 426640 224527 426646 224539
rect 426698 224527 426704 224579
rect 427312 224527 427318 224579
rect 427370 224567 427376 224579
rect 428176 224567 428182 224579
rect 427370 224539 428182 224567
rect 427370 224527 427376 224539
rect 428176 224527 428182 224539
rect 428234 224527 428240 224579
rect 429040 224527 429046 224579
rect 429098 224567 429104 224579
rect 438064 224567 438070 224579
rect 429098 224539 438070 224567
rect 429098 224527 429104 224539
rect 438064 224527 438070 224539
rect 438122 224527 438128 224579
rect 354256 224453 354262 224505
rect 354314 224493 354320 224505
rect 438736 224493 438742 224505
rect 354314 224465 438742 224493
rect 354314 224453 354320 224465
rect 438736 224453 438742 224465
rect 438794 224453 438800 224505
rect 354448 224379 354454 224431
rect 354506 224419 354512 224431
rect 421072 224419 421078 224431
rect 354506 224391 421078 224419
rect 354506 224379 354512 224391
rect 421072 224379 421078 224391
rect 421130 224379 421136 224431
rect 422320 224379 422326 224431
rect 422378 224419 422384 224431
rect 436912 224419 436918 224431
rect 422378 224391 436918 224419
rect 422378 224379 422384 224391
rect 436912 224379 436918 224391
rect 436970 224379 436976 224431
rect 351376 224305 351382 224357
rect 351434 224345 351440 224357
rect 439120 224345 439126 224357
rect 351434 224317 439126 224345
rect 351434 224305 351440 224317
rect 439120 224305 439126 224317
rect 439178 224305 439184 224357
rect 364624 224271 364630 224283
rect 351394 224243 364630 224271
rect 325840 224157 325846 224209
rect 325898 224197 325904 224209
rect 338320 224197 338326 224209
rect 325898 224169 338326 224197
rect 325898 224157 325904 224169
rect 338320 224157 338326 224169
rect 338378 224157 338384 224209
rect 351394 224123 351422 224243
rect 364624 224231 364630 224243
rect 364682 224231 364688 224283
rect 391888 224231 391894 224283
rect 391946 224271 391952 224283
rect 444304 224271 444310 224283
rect 391946 224243 444310 224271
rect 391946 224231 391952 224243
rect 444304 224231 444310 224243
rect 444362 224231 444368 224283
rect 351472 224157 351478 224209
rect 351530 224197 351536 224209
rect 351530 224169 378782 224197
rect 351530 224157 351536 224169
rect 336994 224095 351422 224123
rect 328048 224009 328054 224061
rect 328106 224049 328112 224061
rect 336994 224049 337022 224095
rect 363856 224083 363862 224135
rect 363914 224123 363920 224135
rect 364336 224123 364342 224135
rect 363914 224095 364342 224123
rect 363914 224083 363920 224095
rect 364336 224083 364342 224095
rect 364394 224083 364400 224135
rect 378754 224123 378782 224169
rect 396016 224157 396022 224209
rect 396074 224197 396080 224209
rect 405424 224197 405430 224209
rect 396074 224169 405430 224197
rect 396074 224157 396080 224169
rect 405424 224157 405430 224169
rect 405482 224157 405488 224209
rect 405712 224157 405718 224209
rect 405770 224197 405776 224209
rect 439504 224197 439510 224209
rect 405770 224169 439510 224197
rect 405770 224157 405776 224169
rect 439504 224157 439510 224169
rect 439562 224157 439568 224209
rect 395824 224123 395830 224135
rect 364450 224095 378686 224123
rect 378754 224095 395830 224123
rect 328106 224021 337022 224049
rect 328106 224009 328112 224021
rect 348592 224009 348598 224061
rect 348650 224049 348656 224061
rect 364450 224049 364478 224095
rect 348650 224021 364478 224049
rect 348650 224009 348656 224021
rect 364624 224009 364630 224061
rect 364682 224049 364688 224061
rect 378544 224049 378550 224061
rect 364682 224021 378550 224049
rect 364682 224009 364688 224021
rect 378544 224009 378550 224021
rect 378602 224009 378608 224061
rect 378658 224049 378686 224095
rect 395824 224083 395830 224095
rect 395882 224083 395888 224135
rect 395920 224083 395926 224135
rect 395978 224123 395984 224135
rect 417712 224123 417718 224135
rect 395978 224095 417718 224123
rect 395978 224083 395984 224095
rect 417712 224083 417718 224095
rect 417770 224083 417776 224135
rect 427312 224123 427318 224135
rect 417826 224095 427318 224123
rect 417826 224049 417854 224095
rect 427312 224083 427318 224095
rect 427370 224083 427376 224135
rect 442480 224123 442486 224135
rect 427714 224095 442486 224123
rect 378658 224021 417854 224049
rect 418096 224009 418102 224061
rect 418154 224049 418160 224061
rect 427600 224049 427606 224061
rect 418154 224021 427606 224049
rect 418154 224009 418160 224021
rect 427600 224009 427606 224021
rect 427658 224009 427664 224061
rect 207376 223935 207382 223987
rect 207434 223935 207440 223987
rect 379312 223935 379318 223987
rect 379370 223975 379376 223987
rect 403216 223975 403222 223987
rect 379370 223947 403222 223975
rect 379370 223935 379376 223947
rect 403216 223935 403222 223947
rect 403274 223935 403280 223987
rect 405136 223935 405142 223987
rect 405194 223975 405200 223987
rect 406096 223975 406102 223987
rect 405194 223947 406102 223975
rect 405194 223935 405200 223947
rect 406096 223935 406102 223947
rect 406154 223935 406160 223987
rect 418000 223935 418006 223987
rect 418058 223975 418064 223987
rect 418192 223975 418198 223987
rect 418058 223947 418198 223975
rect 418058 223935 418064 223947
rect 418192 223935 418198 223947
rect 418250 223935 418256 223987
rect 418480 223935 418486 223987
rect 418538 223975 418544 223987
rect 427714 223975 427742 224095
rect 442480 224083 442486 224095
rect 442538 224083 442544 224135
rect 428176 224009 428182 224061
rect 428234 224049 428240 224061
rect 440272 224049 440278 224061
rect 428234 224021 440278 224049
rect 428234 224009 428240 224021
rect 440272 224009 440278 224021
rect 440330 224009 440336 224061
rect 418538 223947 427742 223975
rect 418538 223935 418544 223947
rect 204304 223787 204310 223839
rect 204362 223827 204368 223839
rect 207394 223827 207422 223935
rect 330448 223861 330454 223913
rect 330506 223901 330512 223913
rect 363856 223901 363862 223913
rect 330506 223873 363862 223901
rect 330506 223861 330512 223873
rect 363856 223861 363862 223873
rect 363914 223861 363920 223913
rect 364336 223861 364342 223913
rect 364394 223901 364400 223913
rect 396016 223901 396022 223913
rect 364394 223873 396022 223901
rect 364394 223861 364400 223873
rect 396016 223861 396022 223873
rect 396074 223861 396080 223913
rect 405424 223861 405430 223913
rect 405482 223901 405488 223913
rect 418096 223901 418102 223913
rect 405482 223873 418102 223901
rect 405482 223861 405488 223873
rect 418096 223861 418102 223873
rect 418154 223861 418160 223913
rect 427600 223861 427606 223913
rect 427658 223901 427664 223913
rect 427658 223873 443630 223901
rect 427658 223861 427664 223873
rect 443602 223839 443630 223873
rect 207664 223827 207670 223839
rect 204362 223799 207670 223827
rect 204362 223787 204368 223799
rect 207664 223787 207670 223799
rect 207722 223787 207728 223839
rect 330256 223787 330262 223839
rect 330314 223787 330320 223839
rect 338320 223787 338326 223839
rect 338378 223827 338384 223839
rect 364240 223827 364246 223839
rect 338378 223799 364246 223827
rect 338378 223787 338384 223799
rect 364240 223787 364246 223799
rect 364298 223787 364304 223839
rect 364354 223799 374270 223827
rect 330274 223753 330302 223787
rect 364354 223753 364382 223799
rect 330274 223725 364382 223753
rect 374242 223753 374270 223799
rect 378544 223787 378550 223839
rect 378602 223827 378608 223839
rect 379312 223827 379318 223839
rect 378602 223799 379318 223827
rect 378602 223787 378608 223799
rect 379312 223787 379318 223799
rect 379370 223787 379376 223839
rect 379408 223787 379414 223839
rect 379466 223827 379472 223839
rect 417904 223827 417910 223839
rect 379466 223799 417910 223827
rect 379466 223787 379472 223799
rect 417904 223787 417910 223799
rect 417962 223787 417968 223839
rect 418000 223787 418006 223839
rect 418058 223827 418064 223839
rect 441712 223827 441718 223839
rect 418058 223799 441718 223827
rect 418058 223787 418064 223799
rect 441712 223787 441718 223799
rect 441770 223787 441776 223839
rect 443584 223787 443590 223839
rect 443642 223787 443648 223839
rect 445072 223787 445078 223839
rect 445130 223787 445136 223839
rect 451792 223787 451798 223839
rect 451850 223827 451856 223839
rect 452032 223827 452038 223839
rect 451850 223799 452038 223827
rect 451850 223787 451856 223799
rect 452032 223787 452038 223799
rect 452090 223787 452096 223839
rect 483856 223787 483862 223839
rect 483914 223827 483920 223839
rect 503200 223827 503206 223839
rect 483914 223799 503206 223827
rect 483914 223787 483920 223799
rect 503200 223787 503206 223799
rect 503258 223787 503264 223839
rect 445090 223753 445118 223787
rect 374242 223725 445118 223753
rect 204496 223235 204502 223247
rect 204418 223207 204502 223235
rect 204418 223013 204446 223207
rect 204496 223195 204502 223207
rect 204554 223195 204560 223247
rect 204496 223047 204502 223099
rect 204554 223087 204560 223099
rect 204976 223087 204982 223099
rect 204554 223059 204982 223087
rect 204554 223047 204560 223059
rect 204976 223047 204982 223059
rect 205034 223047 205040 223099
rect 204418 222985 204926 223013
rect 204898 222877 204926 222985
rect 204880 222825 204886 222877
rect 204938 222825 204944 222877
rect 641008 222381 641014 222433
rect 641066 222421 641072 222433
rect 649648 222421 649654 222433
rect 641066 222393 649654 222421
rect 641066 222381 641072 222393
rect 649648 222381 649654 222393
rect 649706 222381 649712 222433
rect 144016 221789 144022 221841
rect 144074 221829 144080 221841
rect 171280 221829 171286 221841
rect 144074 221801 171286 221829
rect 144074 221789 144080 221801
rect 171280 221789 171286 221801
rect 171338 221789 171344 221841
rect 199984 221789 199990 221841
rect 200042 221829 200048 221841
rect 200080 221829 200086 221841
rect 200042 221801 200086 221829
rect 200042 221789 200048 221801
rect 200080 221789 200086 221801
rect 200138 221789 200144 221841
rect 141520 221715 141526 221767
rect 141578 221755 141584 221767
rect 198736 221755 198742 221767
rect 141578 221727 198742 221755
rect 141578 221715 141584 221727
rect 198736 221715 198742 221727
rect 198794 221715 198800 221767
rect 641296 221345 641302 221397
rect 641354 221385 641360 221397
rect 650320 221385 650326 221397
rect 641354 221357 650326 221385
rect 641354 221345 641360 221357
rect 650320 221345 650326 221357
rect 650378 221345 650384 221397
rect 42352 221049 42358 221101
rect 42410 221089 42416 221101
rect 45712 221089 45718 221101
rect 42410 221061 45718 221089
rect 42410 221049 42416 221061
rect 45712 221049 45718 221061
rect 45770 221049 45776 221101
rect 641296 220753 641302 220805
rect 641354 220793 641360 220805
rect 650032 220793 650038 220805
rect 641354 220765 650038 220793
rect 641354 220753 641360 220765
rect 650032 220753 650038 220765
rect 650090 220753 650096 220805
rect 42352 220309 42358 220361
rect 42410 220349 42416 220361
rect 45808 220349 45814 220361
rect 42410 220321 45814 220349
rect 42410 220309 42416 220321
rect 45808 220309 45814 220321
rect 45866 220309 45872 220361
rect 42352 219421 42358 219473
rect 42410 219461 42416 219473
rect 45520 219461 45526 219473
rect 42410 219433 45526 219461
rect 42410 219421 42416 219433
rect 45520 219421 45526 219433
rect 45578 219421 45584 219473
rect 144112 218977 144118 219029
rect 144170 219017 144176 219029
rect 149584 219017 149590 219029
rect 144170 218989 149590 219017
rect 144170 218977 144176 218989
rect 149584 218977 149590 218989
rect 149642 218977 149648 219029
rect 144016 218903 144022 218955
rect 144074 218943 144080 218955
rect 165520 218943 165526 218955
rect 144074 218915 165526 218943
rect 144074 218903 144080 218915
rect 165520 218903 165526 218915
rect 165578 218903 165584 218955
rect 141904 218829 141910 218881
rect 141962 218869 141968 218881
rect 199024 218869 199030 218881
rect 141962 218841 199030 218869
rect 141962 218829 141968 218841
rect 199024 218829 199030 218841
rect 199082 218829 199088 218881
rect 142192 218755 142198 218807
rect 142250 218795 142256 218807
rect 198736 218795 198742 218807
rect 142250 218767 198742 218795
rect 142250 218755 142256 218767
rect 198736 218755 198742 218767
rect 198794 218755 198800 218807
rect 140848 218681 140854 218733
rect 140906 218721 140912 218733
rect 198832 218721 198838 218733
rect 140906 218693 198838 218721
rect 140906 218681 140912 218693
rect 198832 218681 198838 218693
rect 198890 218681 198896 218733
rect 149680 218607 149686 218659
rect 149738 218647 149744 218659
rect 198928 218647 198934 218659
rect 149738 218619 198934 218647
rect 149738 218607 149744 218619
rect 198928 218607 198934 218619
rect 198986 218607 198992 218659
rect 155440 218533 155446 218585
rect 155498 218573 155504 218585
rect 198736 218573 198742 218585
rect 155498 218545 198742 218573
rect 155498 218533 155504 218545
rect 198736 218533 198742 218545
rect 198794 218533 198800 218585
rect 144016 218015 144022 218067
rect 144074 218055 144080 218067
rect 159760 218055 159766 218067
rect 144074 218027 159766 218055
rect 144074 218015 144080 218027
rect 159760 218015 159766 218027
rect 159818 218015 159824 218067
rect 141328 215943 141334 215995
rect 141386 215983 141392 215995
rect 199024 215983 199030 215995
rect 141386 215955 199030 215983
rect 141386 215943 141392 215955
rect 199024 215943 199030 215955
rect 199082 215943 199088 215995
rect 141712 215869 141718 215921
rect 141770 215909 141776 215921
rect 198928 215909 198934 215921
rect 141770 215881 198934 215909
rect 141770 215869 141776 215881
rect 198928 215869 198934 215881
rect 198986 215869 198992 215921
rect 164080 215795 164086 215847
rect 164138 215835 164144 215847
rect 198736 215835 198742 215847
rect 164138 215807 198742 215835
rect 164138 215795 164144 215807
rect 198736 215795 198742 215807
rect 198794 215795 198800 215847
rect 175600 215721 175606 215773
rect 175658 215761 175664 215773
rect 198832 215761 198838 215773
rect 175658 215733 198838 215761
rect 175658 215721 175664 215733
rect 198832 215721 198838 215733
rect 198890 215721 198896 215773
rect 181360 215647 181366 215699
rect 181418 215687 181424 215699
rect 198736 215687 198742 215699
rect 181418 215659 198742 215687
rect 181418 215647 181424 215659
rect 198736 215647 198742 215659
rect 198794 215647 198800 215699
rect 187120 215573 187126 215625
rect 187178 215613 187184 215625
rect 198832 215613 198838 215625
rect 187178 215585 198838 215613
rect 187178 215573 187184 215585
rect 198832 215573 198838 215585
rect 198890 215573 198896 215625
rect 144016 213205 144022 213257
rect 144074 213245 144080 213257
rect 154000 213245 154006 213257
rect 144074 213217 154006 213245
rect 144074 213205 144080 213217
rect 154000 213205 154006 213217
rect 154058 213205 154064 213257
rect 146512 213131 146518 213183
rect 146570 213171 146576 213183
rect 148336 213171 148342 213183
rect 146570 213143 148342 213171
rect 146570 213131 146576 213143
rect 148336 213131 148342 213143
rect 148394 213131 148400 213183
rect 139984 213057 139990 213109
rect 140042 213097 140048 213109
rect 198736 213097 198742 213109
rect 140042 213069 198742 213097
rect 140042 213057 140048 213069
rect 198736 213057 198742 213069
rect 198794 213057 198800 213109
rect 144016 210245 144022 210297
rect 144074 210285 144080 210297
rect 185680 210285 185686 210297
rect 144074 210257 185686 210285
rect 144074 210245 144080 210257
rect 185680 210245 185686 210257
rect 185738 210245 185744 210297
rect 639760 210245 639766 210297
rect 639818 210285 639824 210297
rect 679696 210285 679702 210297
rect 639818 210257 679702 210285
rect 639818 210245 639824 210257
rect 679696 210245 679702 210257
rect 679754 210245 679760 210297
rect 144016 207359 144022 207411
rect 144074 207399 144080 207411
rect 148048 207399 148054 207411
rect 144074 207371 148054 207399
rect 144074 207359 144080 207371
rect 148048 207359 148054 207371
rect 148106 207359 148112 207411
rect 204592 207359 204598 207411
rect 204650 207399 204656 207411
rect 204880 207399 204886 207411
rect 204650 207371 204886 207399
rect 204650 207359 204656 207371
rect 204880 207359 204886 207371
rect 204938 207359 204944 207411
rect 674512 205731 674518 205783
rect 674570 205771 674576 205783
rect 675472 205771 675478 205783
rect 674570 205743 675478 205771
rect 674570 205731 674576 205743
rect 675472 205731 675478 205743
rect 675530 205731 675536 205783
rect 146800 205139 146806 205191
rect 146858 205179 146864 205191
rect 156880 205179 156886 205191
rect 146858 205151 156886 205179
rect 146858 205139 146864 205151
rect 156880 205139 156886 205151
rect 156938 205139 156944 205191
rect 675088 205031 675094 205043
rect 675010 205003 675094 205031
rect 675010 204821 675038 205003
rect 675088 204991 675094 205003
rect 675146 204991 675152 205043
rect 675184 204991 675190 205043
rect 675242 205031 675248 205043
rect 675472 205031 675478 205043
rect 675242 205003 675478 205031
rect 675242 204991 675248 205003
rect 675472 204991 675478 205003
rect 675530 204991 675536 205043
rect 674992 204769 674998 204821
rect 675050 204769 675056 204821
rect 146800 204473 146806 204525
rect 146858 204513 146864 204525
rect 182800 204513 182806 204525
rect 146858 204485 182806 204513
rect 146858 204473 146864 204485
rect 182800 204473 182806 204485
rect 182858 204473 182864 204525
rect 42352 204325 42358 204377
rect 42410 204365 42416 204377
rect 44560 204365 44566 204377
rect 42410 204337 44566 204365
rect 42410 204325 42416 204337
rect 44560 204325 44566 204337
rect 44618 204325 44624 204377
rect 144976 201587 144982 201639
rect 145034 201627 145040 201639
rect 179920 201627 179926 201639
rect 145034 201599 179926 201627
rect 145034 201587 145040 201599
rect 179920 201587 179926 201599
rect 179978 201587 179984 201639
rect 200656 201513 200662 201565
rect 200714 201553 200720 201565
rect 200944 201553 200950 201565
rect 200714 201525 200950 201553
rect 200714 201513 200720 201525
rect 200944 201513 200950 201525
rect 201002 201513 201008 201565
rect 42064 201291 42070 201343
rect 42122 201331 42128 201343
rect 42928 201331 42934 201343
rect 42122 201303 42934 201331
rect 42122 201291 42128 201303
rect 42928 201291 42934 201303
rect 42986 201291 42992 201343
rect 674416 201291 674422 201343
rect 674474 201331 674480 201343
rect 675376 201331 675382 201343
rect 674474 201303 675382 201331
rect 674474 201291 674480 201303
rect 675376 201291 675382 201303
rect 675434 201291 675440 201343
rect 37360 200773 37366 200825
rect 37418 200813 37424 200825
rect 41776 200813 41782 200825
rect 37418 200785 41782 200813
rect 37418 200773 37424 200785
rect 41776 200773 41782 200785
rect 41834 200773 41840 200825
rect 42736 198849 42742 198901
rect 42794 198889 42800 198901
rect 43312 198889 43318 198901
rect 42794 198861 43318 198889
rect 42794 198849 42800 198861
rect 43312 198849 43318 198861
rect 43370 198849 43376 198901
rect 42832 198775 42838 198827
rect 42890 198815 42896 198827
rect 43216 198815 43222 198827
rect 42890 198787 43222 198815
rect 42890 198775 42896 198787
rect 43216 198775 43222 198787
rect 43274 198775 43280 198827
rect 144976 198775 144982 198827
rect 145034 198815 145040 198827
rect 162640 198815 162646 198827
rect 145034 198787 162646 198815
rect 145034 198775 145040 198787
rect 162640 198775 162646 198787
rect 162698 198775 162704 198827
rect 144400 198701 144406 198753
rect 144458 198741 144464 198753
rect 197296 198741 197302 198753
rect 144458 198713 197302 198741
rect 144458 198701 144464 198713
rect 197296 198701 197302 198713
rect 197354 198701 197360 198753
rect 41872 198183 41878 198235
rect 41930 198223 41936 198235
rect 42352 198223 42358 198235
rect 41930 198195 42358 198223
rect 41930 198183 41936 198195
rect 42352 198183 42358 198195
rect 42410 198183 42416 198235
rect 674800 197591 674806 197643
rect 674858 197631 674864 197643
rect 675376 197631 675382 197643
rect 674858 197603 675382 197631
rect 674858 197591 674864 197603
rect 675376 197591 675382 197603
rect 675434 197591 675440 197643
rect 41968 197443 41974 197495
rect 42026 197483 42032 197495
rect 42448 197483 42454 197495
rect 42026 197455 42454 197483
rect 42026 197443 42032 197455
rect 42448 197443 42454 197455
rect 42506 197443 42512 197495
rect 41776 197369 41782 197421
rect 41834 197369 41840 197421
rect 41794 197199 41822 197369
rect 41776 197147 41782 197199
rect 41834 197147 41840 197199
rect 674128 196999 674134 197051
rect 674186 197039 674192 197051
rect 675472 197039 675478 197051
rect 674186 197011 675478 197039
rect 674186 196999 674192 197011
rect 675472 196999 675478 197011
rect 675530 196999 675536 197051
rect 674704 196555 674710 196607
rect 674762 196595 674768 196607
rect 675376 196595 675382 196607
rect 674762 196567 675382 196595
rect 674762 196555 674768 196567
rect 675376 196555 675382 196567
rect 675434 196555 675440 196607
rect 639568 195815 639574 195867
rect 639626 195855 639632 195867
rect 639952 195855 639958 195867
rect 639626 195827 639958 195855
rect 639626 195815 639632 195827
rect 639952 195815 639958 195827
rect 640010 195815 640016 195867
rect 42160 195297 42166 195349
rect 42218 195337 42224 195349
rect 42352 195337 42358 195349
rect 42218 195309 42358 195337
rect 42218 195297 42224 195309
rect 42352 195297 42358 195309
rect 42410 195297 42416 195349
rect 42352 195149 42358 195201
rect 42410 195189 42416 195201
rect 43216 195189 43222 195201
rect 42410 195161 43222 195189
rect 42410 195149 42416 195161
rect 43216 195149 43222 195161
rect 43274 195149 43280 195201
rect 42064 194483 42070 194535
rect 42122 194523 42128 194535
rect 47632 194523 47638 194535
rect 42122 194495 47638 194523
rect 42122 194483 42128 194495
rect 47632 194483 47638 194495
rect 47690 194483 47696 194535
rect 42064 193447 42070 193499
rect 42122 193487 42128 193499
rect 43312 193487 43318 193499
rect 42122 193459 43318 193487
rect 42122 193447 42128 193459
rect 43312 193447 43318 193459
rect 43370 193447 43376 193499
rect 144592 193077 144598 193129
rect 144650 193117 144656 193129
rect 148528 193117 148534 193129
rect 144650 193089 148534 193117
rect 144650 193077 144656 193089
rect 148528 193077 148534 193089
rect 148586 193077 148592 193129
rect 146800 193003 146806 193055
rect 146858 193043 146864 193055
rect 191536 193043 191542 193055
rect 146858 193015 191542 193043
rect 146858 193003 146864 193015
rect 191536 193003 191542 193015
rect 191594 193003 191600 193055
rect 42160 192189 42166 192241
rect 42218 192229 42224 192241
rect 43024 192229 43030 192241
rect 42218 192201 43030 192229
rect 42218 192189 42224 192201
rect 43024 192189 43030 192201
rect 43082 192189 43088 192241
rect 42064 191449 42070 191501
rect 42122 191489 42128 191501
rect 42352 191489 42358 191501
rect 42122 191461 42358 191489
rect 42122 191449 42128 191461
rect 42352 191449 42358 191461
rect 42410 191449 42416 191501
rect 42160 191005 42166 191057
rect 42218 191045 42224 191057
rect 43120 191045 43126 191057
rect 42218 191017 43126 191045
rect 42218 191005 42224 191017
rect 43120 191005 43126 191017
rect 43178 191005 43184 191057
rect 144304 190117 144310 190169
rect 144362 190157 144368 190169
rect 188656 190157 188662 190169
rect 144362 190129 188662 190157
rect 144362 190117 144368 190129
rect 188656 190117 188662 190129
rect 188714 190117 188720 190169
rect 42256 189229 42262 189281
rect 42314 189269 42320 189281
rect 42640 189269 42646 189281
rect 42314 189241 42646 189269
rect 42314 189229 42320 189241
rect 42640 189229 42646 189241
rect 42698 189229 42704 189281
rect 42160 187823 42166 187875
rect 42218 187863 42224 187875
rect 42736 187863 42742 187875
rect 42218 187835 42742 187863
rect 42218 187823 42224 187835
rect 42736 187823 42742 187835
rect 42794 187823 42800 187875
rect 146800 187231 146806 187283
rect 146858 187271 146864 187283
rect 185776 187271 185782 187283
rect 146858 187243 185782 187271
rect 146858 187231 146864 187243
rect 185776 187231 185782 187243
rect 185834 187231 185840 187283
rect 200752 187231 200758 187283
rect 200810 187271 200816 187283
rect 201040 187271 201046 187283
rect 200810 187243 201046 187271
rect 200810 187231 200816 187243
rect 201040 187231 201046 187243
rect 201098 187231 201104 187283
rect 42160 187083 42166 187135
rect 42218 187123 42224 187135
rect 42640 187123 42646 187135
rect 42218 187095 42646 187123
rect 42218 187083 42224 187095
rect 42640 187083 42646 187095
rect 42698 187083 42704 187135
rect 42064 186639 42070 186691
rect 42122 186679 42128 186691
rect 42448 186679 42454 186691
rect 42122 186651 42454 186679
rect 42122 186639 42128 186651
rect 42448 186639 42454 186651
rect 42506 186639 42512 186691
rect 146800 184419 146806 184471
rect 146858 184459 146864 184471
rect 180016 184459 180022 184471
rect 146858 184431 180022 184459
rect 146858 184419 146864 184431
rect 180016 184419 180022 184431
rect 180074 184419 180080 184471
rect 146608 184345 146614 184397
rect 146666 184385 146672 184397
rect 182896 184385 182902 184397
rect 146666 184357 182902 184385
rect 146666 184345 146672 184357
rect 182896 184345 182902 184357
rect 182954 184345 182960 184397
rect 655312 184345 655318 184397
rect 655370 184385 655376 184397
rect 674416 184385 674422 184397
rect 655370 184357 674422 184385
rect 655370 184345 655376 184357
rect 674416 184345 674422 184357
rect 674474 184345 674480 184397
rect 661168 183901 661174 183953
rect 661226 183941 661232 183953
rect 674704 183941 674710 183953
rect 661226 183913 674710 183941
rect 661226 183901 661232 183913
rect 674704 183901 674710 183913
rect 674762 183901 674768 183953
rect 144976 182865 144982 182917
rect 145034 182905 145040 182917
rect 146512 182905 146518 182917
rect 145034 182877 146518 182905
rect 145034 182865 145040 182877
rect 146512 182865 146518 182877
rect 146570 182865 146576 182917
rect 666736 182865 666742 182917
rect 666794 182905 666800 182917
rect 674416 182905 674422 182917
rect 666794 182877 674422 182905
rect 666794 182865 666800 182877
rect 674416 182865 674422 182877
rect 674474 182865 674480 182917
rect 144688 181533 144694 181585
rect 144746 181573 144752 181585
rect 148912 181573 148918 181585
rect 144746 181545 148918 181573
rect 144746 181533 144752 181545
rect 148912 181533 148918 181545
rect 148970 181533 148976 181585
rect 146800 181459 146806 181511
rect 146858 181499 146864 181511
rect 168496 181499 168502 181511
rect 146858 181471 168502 181499
rect 146858 181459 146864 181471
rect 168496 181459 168502 181471
rect 168554 181459 168560 181511
rect 200656 181459 200662 181511
rect 200714 181499 200720 181511
rect 200848 181499 200854 181511
rect 200714 181471 200854 181499
rect 200714 181459 200720 181471
rect 200848 181459 200854 181471
rect 200906 181459 200912 181511
rect 144880 181311 144886 181363
rect 144938 181351 144944 181363
rect 146800 181351 146806 181363
rect 144938 181323 146806 181351
rect 144938 181311 144944 181323
rect 146800 181311 146806 181323
rect 146858 181311 146864 181363
rect 144016 178573 144022 178625
rect 144074 178613 144080 178625
rect 177136 178613 177142 178625
rect 144074 178585 177142 178613
rect 144074 178573 144080 178585
rect 177136 178573 177142 178585
rect 177194 178573 177200 178625
rect 144976 175761 144982 175813
rect 145034 175801 145040 175813
rect 149008 175801 149014 175813
rect 145034 175773 149014 175801
rect 145034 175761 145040 175773
rect 149008 175761 149014 175773
rect 149066 175761 149072 175813
rect 144976 172801 144982 172853
rect 145034 172841 145040 172853
rect 149296 172841 149302 172853
rect 145034 172813 149302 172841
rect 145034 172801 145040 172813
rect 149296 172801 149302 172813
rect 149354 172801 149360 172853
rect 144976 169915 144982 169967
rect 145034 169955 145040 169967
rect 151216 169955 151222 169967
rect 145034 169927 151222 169955
rect 145034 169915 145040 169927
rect 151216 169915 151222 169927
rect 151274 169915 151280 169967
rect 144976 167843 144982 167895
rect 145034 167883 145040 167895
rect 156976 167883 156982 167895
rect 145034 167855 156982 167883
rect 145034 167843 145040 167855
rect 156976 167843 156982 167855
rect 157034 167843 157040 167895
rect 641488 167177 641494 167229
rect 641546 167217 641552 167229
rect 674704 167217 674710 167229
rect 641546 167189 674710 167217
rect 641546 167177 641552 167189
rect 674704 167177 674710 167189
rect 674762 167177 674768 167229
rect 144976 167029 144982 167081
rect 145034 167069 145040 167081
rect 149488 167069 149494 167081
rect 145034 167041 149494 167069
rect 145034 167029 145040 167041
rect 149488 167029 149494 167041
rect 149546 167029 149552 167081
rect 144976 164217 144982 164269
rect 145034 164257 145040 164269
rect 149680 164257 149686 164269
rect 145034 164229 149686 164257
rect 145034 164217 145040 164229
rect 149680 164217 149686 164229
rect 149738 164217 149744 164269
rect 642160 164217 642166 164269
rect 642218 164257 642224 164269
rect 674704 164257 674710 164269
rect 642218 164229 674710 164257
rect 642218 164217 642224 164229
rect 674704 164217 674710 164229
rect 674762 164217 674768 164269
rect 144016 164143 144022 164195
rect 144074 164183 144080 164195
rect 194416 164183 194422 164195
rect 144074 164155 194422 164183
rect 144074 164143 144080 164155
rect 194416 164143 194422 164155
rect 194474 164143 194480 164195
rect 642064 164143 642070 164195
rect 642122 164183 642128 164195
rect 674608 164183 674614 164195
rect 642122 164155 674614 164183
rect 642122 164143 642128 164155
rect 674608 164143 674614 164155
rect 674666 164143 674672 164195
rect 675184 163033 675190 163085
rect 675242 163073 675248 163085
rect 676912 163073 676918 163085
rect 675242 163045 676918 163073
rect 675242 163033 675248 163045
rect 676912 163033 676918 163045
rect 676970 163033 676976 163085
rect 675088 162071 675094 162123
rect 675146 162111 675152 162123
rect 676816 162111 676822 162123
rect 675146 162083 676822 162111
rect 675146 162071 675152 162083
rect 676816 162071 676822 162083
rect 676874 162071 676880 162123
rect 144304 161405 144310 161457
rect 144362 161445 144368 161457
rect 148144 161445 148150 161457
rect 144362 161417 148150 161445
rect 144362 161405 144368 161417
rect 148144 161405 148150 161417
rect 148202 161405 148208 161457
rect 144976 161331 144982 161383
rect 145034 161371 145040 161383
rect 171376 161371 171382 161383
rect 145034 161343 171382 161371
rect 145034 161331 145040 161343
rect 171376 161331 171382 161343
rect 171434 161331 171440 161383
rect 144208 161257 144214 161309
rect 144266 161297 144272 161309
rect 174256 161297 174262 161309
rect 144266 161269 174262 161297
rect 144266 161257 144272 161269
rect 174256 161257 174262 161269
rect 174314 161257 174320 161309
rect 144496 161109 144502 161161
rect 144554 161149 144560 161161
rect 144880 161149 144886 161161
rect 144554 161121 144886 161149
rect 144554 161109 144560 161121
rect 144880 161109 144886 161121
rect 144938 161109 144944 161161
rect 675664 160961 675670 161013
rect 675722 160961 675728 161013
rect 674416 160739 674422 160791
rect 674474 160779 674480 160791
rect 675376 160779 675382 160791
rect 674474 160751 675382 160779
rect 674474 160739 674480 160751
rect 675376 160739 675382 160751
rect 675434 160739 675440 160791
rect 675682 160051 675710 160961
rect 675664 159999 675670 160051
rect 675722 159999 675728 160051
rect 144304 158445 144310 158497
rect 144362 158485 144368 158497
rect 147952 158485 147958 158497
rect 144362 158457 147958 158485
rect 144362 158445 144368 158457
rect 147952 158445 147958 158457
rect 148010 158445 148016 158497
rect 674896 157039 674902 157091
rect 674954 157079 674960 157091
rect 675088 157079 675094 157091
rect 674954 157051 675094 157079
rect 674954 157039 674960 157051
rect 675088 157039 675094 157051
rect 675146 157039 675152 157091
rect 674800 156891 674806 156943
rect 674858 156931 674864 156943
rect 675472 156931 675478 156943
rect 674858 156903 675478 156931
rect 674858 156891 674864 156903
rect 675472 156891 675478 156903
rect 675530 156891 675536 156943
rect 144304 156003 144310 156055
rect 144362 156043 144368 156055
rect 149104 156043 149110 156055
rect 144362 156015 149110 156043
rect 144362 156003 144368 156015
rect 149104 156003 149110 156015
rect 149162 156003 149168 156055
rect 144496 155559 144502 155611
rect 144554 155599 144560 155611
rect 165616 155599 165622 155611
rect 144554 155571 165622 155599
rect 144554 155559 144560 155571
rect 165616 155559 165622 155571
rect 165674 155559 165680 155611
rect 144496 152747 144502 152799
rect 144554 152787 144560 152799
rect 159856 152787 159862 152799
rect 144554 152759 159862 152787
rect 144554 152747 144560 152759
rect 159856 152747 159862 152759
rect 159914 152747 159920 152799
rect 144304 152673 144310 152725
rect 144362 152713 144368 152725
rect 202960 152713 202966 152725
rect 144362 152685 202966 152713
rect 144362 152673 144368 152685
rect 202960 152673 202966 152685
rect 203018 152673 203024 152725
rect 674224 152599 674230 152651
rect 674282 152639 674288 152651
rect 675376 152639 675382 152651
rect 674282 152611 675382 152639
rect 674282 152599 674288 152611
rect 675376 152599 675382 152611
rect 675434 152599 675440 152651
rect 674032 152007 674038 152059
rect 674090 152047 674096 152059
rect 675472 152047 675478 152059
rect 674090 152019 675478 152047
rect 674090 152007 674096 152019
rect 675472 152007 675478 152019
rect 675530 152007 675536 152059
rect 674512 151489 674518 151541
rect 674570 151529 674576 151541
rect 675376 151529 675382 151541
rect 674570 151501 675382 151529
rect 674570 151489 674576 151501
rect 675376 151489 675382 151501
rect 675434 151489 675440 151541
rect 144304 149861 144310 149913
rect 144362 149901 144368 149913
rect 154096 149901 154102 149913
rect 144362 149873 154102 149901
rect 144362 149861 144368 149873
rect 154096 149861 154102 149873
rect 154154 149861 154160 149913
rect 144496 149787 144502 149839
rect 144554 149827 144560 149839
rect 203056 149827 203062 149839
rect 144554 149799 203062 149827
rect 144554 149787 144560 149799
rect 203056 149787 203062 149799
rect 203114 149787 203120 149839
rect 640144 149787 640150 149839
rect 640202 149827 640208 149839
rect 643600 149827 643606 149839
rect 640202 149799 643606 149827
rect 640202 149787 640208 149799
rect 643600 149787 643606 149799
rect 643658 149787 643664 149839
rect 144208 149047 144214 149099
rect 144266 149087 144272 149099
rect 144496 149087 144502 149099
rect 144266 149059 144502 149087
rect 144266 149047 144272 149059
rect 144496 149047 144502 149059
rect 144554 149047 144560 149099
rect 144496 147163 144502 147175
rect 144130 147135 144502 147163
rect 144130 146941 144158 147135
rect 144496 147123 144502 147135
rect 144554 147123 144560 147175
rect 144208 147049 144214 147101
rect 144266 147089 144272 147101
rect 147856 147089 147862 147101
rect 144266 147061 147862 147089
rect 144266 147049 144272 147061
rect 147856 147049 147862 147061
rect 147914 147049 147920 147101
rect 144304 146975 144310 147027
rect 144362 147015 144368 147027
rect 162736 147015 162742 147027
rect 144362 146987 162742 147015
rect 144362 146975 144368 146987
rect 162736 146975 162742 146987
rect 162794 146975 162800 147027
rect 144208 146941 144214 146953
rect 144130 146913 144214 146941
rect 144208 146901 144214 146913
rect 144266 146901 144272 146953
rect 144496 146901 144502 146953
rect 144554 146941 144560 146953
rect 163024 146941 163030 146953
rect 144554 146913 163030 146941
rect 144554 146901 144560 146913
rect 163024 146901 163030 146913
rect 163082 146901 163088 146953
rect 144304 144089 144310 144141
rect 144362 144129 144368 144141
rect 147760 144129 147766 144141
rect 144362 144101 147766 144129
rect 144362 144089 144368 144101
rect 147760 144089 147766 144101
rect 147818 144089 147824 144141
rect 144496 144015 144502 144067
rect 144554 144055 144560 144067
rect 162832 144055 162838 144067
rect 144554 144027 162838 144055
rect 144554 144015 144560 144027
rect 162832 144015 162838 144027
rect 162890 144015 162896 144067
rect 674320 142649 674326 142661
rect 659554 142621 674326 142649
rect 642160 142535 642166 142587
rect 642218 142575 642224 142587
rect 659554 142575 659582 142621
rect 674320 142609 674326 142621
rect 674378 142649 674384 142661
rect 679696 142649 679702 142661
rect 674378 142621 679702 142649
rect 674378 142609 674384 142621
rect 679696 142609 679702 142621
rect 679754 142609 679760 142661
rect 642218 142547 659582 142575
rect 642218 142535 642224 142547
rect 144496 142239 144502 142291
rect 144554 142279 144560 142291
rect 157072 142279 157078 142291
rect 144554 142251 157078 142279
rect 144554 142239 144560 142251
rect 157072 142239 157078 142251
rect 157130 142239 157136 142291
rect 144304 141129 144310 141181
rect 144362 141169 144368 141181
rect 203152 141169 203158 141181
rect 144362 141141 203158 141169
rect 144362 141129 144368 141141
rect 203152 141129 203158 141141
rect 203210 141129 203216 141181
rect 143920 139427 143926 139479
rect 143978 139467 143984 139479
rect 144208 139467 144214 139479
rect 143978 139439 144214 139467
rect 143978 139427 143984 139439
rect 144208 139427 144214 139439
rect 144266 139427 144272 139479
rect 655216 138539 655222 138591
rect 655274 138579 655280 138591
rect 674704 138579 674710 138591
rect 655274 138551 674710 138579
rect 655274 138539 655280 138551
rect 674704 138539 674710 138551
rect 674762 138539 674768 138591
rect 144208 138391 144214 138443
rect 144266 138431 144272 138443
rect 151312 138431 151318 138443
rect 144266 138403 151318 138431
rect 144266 138391 144272 138403
rect 151312 138391 151318 138403
rect 151370 138391 151376 138443
rect 655120 138391 655126 138443
rect 655178 138431 655184 138443
rect 674416 138431 674422 138443
rect 655178 138403 674422 138431
rect 655178 138391 655184 138403
rect 674416 138391 674422 138403
rect 674474 138391 674480 138443
rect 144304 138317 144310 138369
rect 144362 138357 144368 138369
rect 162928 138357 162934 138369
rect 144362 138329 162934 138357
rect 144362 138317 144368 138329
rect 162928 138317 162934 138329
rect 162986 138317 162992 138369
rect 144400 138243 144406 138295
rect 144458 138243 144464 138295
rect 144496 138243 144502 138295
rect 144554 138283 144560 138295
rect 203248 138283 203254 138295
rect 144554 138255 203254 138283
rect 144554 138243 144560 138255
rect 203248 138243 203254 138255
rect 203306 138243 203312 138295
rect 144418 138073 144446 138243
rect 143920 138021 143926 138073
rect 143978 138061 143984 138073
rect 144304 138061 144310 138073
rect 143978 138033 144310 138061
rect 143978 138021 143984 138033
rect 144304 138021 144310 138033
rect 144362 138021 144368 138073
rect 144400 138021 144406 138073
rect 144458 138021 144464 138073
rect 655408 135579 655414 135631
rect 655466 135619 655472 135631
rect 674704 135619 674710 135631
rect 655466 135591 674710 135619
rect 655466 135579 655472 135591
rect 674704 135579 674710 135591
rect 674762 135579 674768 135631
rect 144208 135545 144214 135557
rect 144034 135517 144214 135545
rect 144034 135397 144062 135517
rect 144208 135505 144214 135517
rect 144266 135505 144272 135557
rect 144112 135431 144118 135483
rect 144170 135471 144176 135483
rect 197392 135471 197398 135483
rect 144170 135443 197398 135471
rect 144170 135431 144176 135443
rect 197392 135431 197398 135443
rect 197450 135431 197456 135483
rect 203344 135397 203350 135409
rect 144034 135369 203350 135397
rect 203344 135357 203350 135369
rect 203402 135357 203408 135409
rect 640720 135357 640726 135409
rect 640778 135397 640784 135409
rect 674704 135397 674710 135409
rect 640778 135369 674710 135397
rect 640778 135357 640784 135369
rect 674704 135357 674710 135369
rect 674762 135357 674768 135409
rect 144016 132619 144022 132671
rect 144074 132659 144080 132671
rect 147664 132659 147670 132671
rect 144074 132631 147670 132659
rect 144074 132619 144080 132631
rect 147664 132619 147670 132631
rect 147722 132619 147728 132671
rect 144208 132545 144214 132597
rect 144266 132585 144272 132597
rect 194512 132585 194518 132597
rect 144266 132557 194518 132585
rect 144266 132545 144272 132557
rect 194512 132545 194518 132557
rect 194570 132545 194576 132597
rect 144112 132471 144118 132523
rect 144170 132511 144176 132523
rect 204976 132511 204982 132523
rect 144170 132483 204982 132511
rect 144170 132471 144176 132483
rect 204976 132471 204982 132483
rect 205034 132471 205040 132523
rect 643600 132471 643606 132523
rect 643658 132511 643664 132523
rect 674416 132511 674422 132523
rect 643658 132483 674422 132511
rect 643658 132471 643664 132483
rect 674416 132471 674422 132483
rect 674474 132471 674480 132523
rect 144112 129659 144118 129711
rect 144170 129699 144176 129711
rect 191632 129699 191638 129711
rect 144170 129671 191638 129699
rect 144170 129659 144176 129671
rect 191632 129659 191638 129671
rect 191690 129659 191696 129711
rect 144208 129585 144214 129637
rect 144266 129625 144272 129637
rect 203440 129625 203446 129637
rect 144266 129597 203446 129625
rect 144266 129585 144272 129597
rect 203440 129585 203446 129597
rect 203498 129585 203504 129637
rect 144112 126773 144118 126825
rect 144170 126813 144176 126825
rect 188752 126813 188758 126825
rect 144170 126785 188758 126813
rect 144170 126773 144176 126785
rect 188752 126773 188758 126785
rect 188810 126773 188816 126825
rect 144208 126699 144214 126751
rect 144266 126739 144272 126751
rect 203536 126739 203542 126751
rect 144266 126711 203542 126739
rect 144266 126699 144272 126711
rect 203536 126699 203542 126711
rect 203594 126699 203600 126751
rect 200848 126625 200854 126677
rect 200906 126665 200912 126677
rect 201040 126665 201046 126677
rect 200906 126637 201046 126665
rect 200906 126625 200912 126637
rect 201040 126625 201046 126637
rect 201098 126625 201104 126677
rect 144208 124035 144214 124087
rect 144266 124075 144272 124087
rect 185872 124075 185878 124087
rect 144266 124047 185878 124075
rect 144266 124035 144272 124047
rect 185872 124035 185878 124047
rect 185930 124035 185936 124087
rect 144016 123961 144022 124013
rect 144074 124001 144080 124013
rect 203728 124001 203734 124013
rect 144074 123973 203734 124001
rect 144074 123961 144080 123973
rect 203728 123961 203734 123973
rect 203786 123961 203792 124013
rect 144112 123887 144118 123939
rect 144170 123927 144176 123939
rect 203632 123927 203638 123939
rect 144170 123899 203638 123927
rect 144170 123887 144176 123899
rect 203632 123887 203638 123899
rect 203690 123887 203696 123939
rect 642064 121223 642070 121275
rect 642122 121263 642128 121275
rect 674704 121263 674710 121275
rect 642122 121235 674710 121263
rect 642122 121223 642128 121235
rect 674704 121223 674710 121235
rect 674762 121223 674768 121275
rect 642160 121149 642166 121201
rect 642218 121189 642224 121201
rect 674800 121189 674806 121201
rect 642218 121161 674806 121189
rect 642218 121149 642224 121161
rect 674800 121149 674806 121161
rect 674858 121149 674864 121201
rect 641392 121075 641398 121127
rect 641450 121115 641456 121127
rect 674608 121115 674614 121127
rect 641450 121087 674614 121115
rect 641450 121075 641456 121087
rect 674608 121075 674614 121087
rect 674666 121075 674672 121127
rect 144208 121001 144214 121053
rect 144266 121041 144272 121053
rect 203824 121041 203830 121053
rect 144266 121013 203830 121041
rect 144266 121001 144272 121013
rect 203824 121001 203830 121013
rect 203882 121001 203888 121053
rect 200464 120927 200470 120979
rect 200522 120967 200528 120979
rect 200752 120967 200758 120979
rect 200522 120939 200758 120967
rect 200522 120927 200528 120939
rect 200752 120927 200758 120939
rect 200810 120927 200816 120979
rect 200848 120927 200854 120979
rect 200906 120967 200912 120979
rect 201040 120967 201046 120979
rect 200906 120939 201046 120967
rect 200906 120927 200912 120939
rect 201040 120927 201046 120939
rect 201098 120927 201104 120979
rect 674896 119521 674902 119573
rect 674954 119561 674960 119573
rect 675088 119561 675094 119573
rect 674954 119533 675094 119561
rect 674954 119521 674960 119533
rect 675088 119521 675094 119533
rect 675146 119521 675152 119573
rect 674128 118485 674134 118537
rect 674186 118525 674192 118537
rect 675280 118525 675286 118537
rect 674186 118497 675286 118525
rect 674186 118485 674192 118497
rect 675280 118485 675286 118497
rect 675338 118485 675344 118537
rect 144208 118263 144214 118315
rect 144266 118303 144272 118315
rect 180112 118303 180118 118315
rect 144266 118275 180118 118303
rect 144266 118263 144272 118275
rect 180112 118263 180118 118275
rect 180170 118263 180176 118315
rect 144112 118189 144118 118241
rect 144170 118229 144176 118241
rect 182992 118229 182998 118241
rect 144170 118201 182998 118229
rect 144170 118189 144176 118201
rect 182992 118189 182998 118201
rect 183050 118189 183056 118241
rect 144016 118115 144022 118167
rect 144074 118155 144080 118167
rect 203920 118155 203926 118167
rect 144074 118127 203926 118155
rect 144074 118115 144080 118127
rect 203920 118115 203926 118127
rect 203978 118115 203984 118167
rect 144208 115303 144214 115355
rect 144266 115343 144272 115355
rect 168592 115343 168598 115355
rect 144266 115315 168598 115343
rect 144266 115303 144272 115315
rect 168592 115303 168598 115315
rect 168650 115303 168656 115355
rect 144112 115229 144118 115281
rect 144170 115269 144176 115281
rect 204016 115269 204022 115281
rect 144170 115241 204022 115269
rect 144170 115229 144176 115241
rect 204016 115229 204022 115241
rect 204074 115229 204080 115281
rect 674896 114785 674902 114837
rect 674954 114825 674960 114837
rect 675088 114825 675094 114837
rect 674954 114797 675094 114825
rect 674954 114785 674960 114797
rect 675088 114785 675094 114797
rect 675146 114785 675152 114837
rect 674128 114119 674134 114171
rect 674186 114159 674192 114171
rect 675376 114159 675382 114171
rect 674186 114131 675382 114159
rect 674186 114119 674192 114131
rect 675376 114119 675382 114131
rect 675434 114119 675440 114171
rect 674224 113601 674230 113653
rect 674282 113641 674288 113653
rect 675184 113641 675190 113653
rect 674282 113613 675190 113641
rect 674282 113601 674288 113613
rect 675184 113601 675190 113613
rect 675242 113601 675248 113653
rect 674512 113305 674518 113357
rect 674570 113345 674576 113357
rect 675088 113345 675094 113357
rect 674570 113317 675094 113345
rect 674570 113305 674576 113317
rect 675088 113305 675094 113317
rect 675146 113305 675152 113357
rect 144208 112417 144214 112469
rect 144266 112457 144272 112469
rect 204112 112457 204118 112469
rect 144266 112429 204118 112457
rect 144266 112417 144272 112429
rect 204112 112417 204118 112429
rect 204170 112417 204176 112469
rect 144112 112343 144118 112395
rect 144170 112383 144176 112395
rect 204880 112383 204886 112395
rect 144170 112355 204886 112383
rect 144170 112343 144176 112355
rect 204880 112343 204886 112355
rect 204938 112343 204944 112395
rect 674416 111159 674422 111211
rect 674474 111199 674480 111211
rect 675376 111199 675382 111211
rect 674474 111171 675382 111199
rect 674474 111159 674480 111171
rect 675376 111159 675382 111171
rect 675434 111159 675440 111211
rect 144208 109605 144214 109657
rect 144266 109645 144272 109657
rect 174352 109645 174358 109657
rect 144266 109617 174358 109645
rect 144266 109605 144272 109617
rect 174352 109605 174358 109617
rect 174410 109605 174416 109657
rect 144016 109531 144022 109583
rect 144074 109571 144080 109583
rect 177232 109571 177238 109583
rect 144074 109543 177238 109571
rect 144074 109531 144080 109543
rect 177232 109531 177238 109543
rect 177290 109531 177296 109583
rect 144112 109457 144118 109509
rect 144170 109497 144176 109509
rect 204208 109497 204214 109509
rect 144170 109469 204214 109497
rect 144170 109457 144176 109469
rect 204208 109457 204214 109469
rect 204266 109457 204272 109509
rect 674800 107533 674806 107585
rect 674858 107573 674864 107585
rect 675376 107573 675382 107585
rect 674858 107545 675382 107573
rect 674858 107533 674864 107545
rect 675376 107533 675382 107545
rect 675434 107533 675440 107585
rect 674032 106867 674038 106919
rect 674090 106907 674096 106919
rect 675472 106907 675478 106919
rect 674090 106879 675478 106907
rect 674090 106867 674096 106879
rect 675472 106867 675478 106879
rect 675530 106867 675536 106919
rect 144208 106571 144214 106623
rect 144266 106611 144272 106623
rect 171472 106611 171478 106623
rect 144266 106583 171478 106611
rect 144266 106571 144272 106583
rect 171472 106571 171478 106583
rect 171530 106571 171536 106623
rect 200464 106497 200470 106549
rect 200522 106537 200528 106549
rect 200656 106537 200662 106549
rect 200522 106509 200662 106537
rect 200522 106497 200528 106509
rect 200656 106497 200662 106509
rect 200714 106497 200720 106549
rect 674608 106349 674614 106401
rect 674666 106389 674672 106401
rect 675376 106389 675382 106401
rect 674666 106361 675382 106389
rect 674666 106349 674672 106361
rect 675376 106349 675382 106361
rect 675434 106349 675440 106401
rect 674320 105165 674326 105217
rect 674378 105205 674384 105217
rect 675376 105205 675382 105217
rect 674378 105177 675382 105205
rect 674378 105165 674384 105177
rect 675376 105165 675382 105177
rect 675434 105165 675440 105217
rect 144112 103833 144118 103885
rect 144170 103873 144176 103885
rect 165712 103873 165718 103885
rect 144170 103845 165718 103873
rect 144170 103833 144176 103845
rect 165712 103833 165718 103845
rect 165770 103833 165776 103885
rect 144208 103759 144214 103811
rect 144266 103799 144272 103811
rect 202768 103799 202774 103811
rect 144266 103771 202774 103799
rect 144266 103759 144272 103771
rect 202768 103759 202774 103771
rect 202826 103759 202832 103811
rect 144016 103685 144022 103737
rect 144074 103725 144080 103737
rect 202864 103725 202870 103737
rect 144074 103697 202870 103725
rect 144074 103685 144080 103697
rect 202864 103685 202870 103697
rect 202922 103685 202928 103737
rect 144208 100799 144214 100851
rect 144266 100839 144272 100851
rect 202672 100839 202678 100851
rect 144266 100811 202678 100839
rect 144266 100799 144272 100811
rect 202672 100799 202678 100811
rect 202730 100799 202736 100851
rect 652528 100799 652534 100851
rect 652586 100839 652592 100851
rect 668176 100839 668182 100851
rect 652586 100811 668182 100839
rect 652586 100799 652592 100811
rect 668176 100799 668182 100811
rect 668234 100799 668240 100851
rect 144208 97913 144214 97965
rect 144266 97953 144272 97965
rect 202576 97953 202582 97965
rect 144266 97925 202582 97953
rect 144266 97913 144272 97925
rect 202576 97913 202582 97925
rect 202634 97913 202640 97965
rect 204976 96507 204982 96559
rect 205034 96507 205040 96559
rect 204880 96285 204886 96337
rect 204938 96325 204944 96337
rect 204994 96325 205022 96507
rect 663280 96433 663286 96485
rect 663338 96473 663344 96485
rect 665200 96473 665206 96485
rect 663338 96445 665206 96473
rect 663338 96433 663344 96445
rect 665200 96433 665206 96445
rect 665258 96433 665264 96485
rect 204938 96297 205022 96325
rect 204938 96285 204944 96297
rect 144112 95101 144118 95153
rect 144170 95141 144176 95153
rect 202192 95141 202198 95153
rect 144170 95113 202198 95141
rect 144170 95101 144176 95113
rect 202192 95101 202198 95113
rect 202250 95101 202256 95153
rect 144208 95027 144214 95079
rect 144266 95067 144272 95079
rect 201808 95067 201814 95079
rect 144266 95039 201814 95067
rect 144266 95027 144272 95039
rect 201808 95027 201814 95039
rect 201866 95027 201872 95079
rect 197200 94953 197206 95005
rect 197258 94993 197264 95005
rect 198736 94993 198742 95005
rect 197258 94965 198742 94993
rect 197258 94953 197264 94965
rect 198736 94953 198742 94965
rect 198794 94953 198800 95005
rect 191440 94879 191446 94931
rect 191498 94919 191504 94931
rect 198928 94919 198934 94931
rect 191498 94891 198934 94919
rect 191498 94879 191504 94891
rect 198928 94879 198934 94891
rect 198986 94879 198992 94931
rect 144208 93547 144214 93599
rect 144266 93587 144272 93599
rect 149776 93587 149782 93599
rect 144266 93559 149782 93587
rect 144266 93547 144272 93559
rect 149776 93547 149782 93559
rect 149834 93547 149840 93599
rect 635248 92807 635254 92859
rect 635306 92847 635312 92859
rect 662512 92847 662518 92859
rect 635306 92819 662518 92847
rect 635306 92807 635312 92819
rect 662512 92807 662518 92819
rect 662570 92807 662576 92859
rect 635056 92733 635062 92785
rect 635114 92773 635120 92785
rect 663088 92773 663094 92785
rect 635114 92745 663094 92773
rect 635114 92733 635120 92745
rect 663088 92733 663094 92745
rect 663146 92733 663152 92785
rect 641008 92659 641014 92711
rect 641066 92699 641072 92711
rect 659824 92699 659830 92711
rect 641066 92671 659830 92699
rect 641066 92659 641072 92671
rect 659824 92659 659830 92671
rect 659882 92659 659888 92711
rect 635344 92585 635350 92637
rect 635402 92625 635408 92637
rect 658864 92625 658870 92637
rect 635402 92597 658870 92625
rect 635402 92585 635408 92597
rect 658864 92585 658870 92597
rect 658922 92585 658928 92637
rect 634960 92511 634966 92563
rect 635018 92551 635024 92563
rect 658288 92551 658294 92563
rect 635018 92523 658294 92551
rect 635018 92511 635024 92523
rect 658288 92511 658294 92523
rect 658346 92511 658352 92563
rect 635440 92437 635446 92489
rect 635498 92477 635504 92489
rect 659344 92477 659350 92489
rect 635498 92449 659350 92477
rect 635498 92437 635504 92449
rect 659344 92437 659350 92449
rect 659402 92437 659408 92489
rect 635152 92363 635158 92415
rect 635210 92403 635216 92415
rect 661168 92403 661174 92415
rect 635210 92375 661174 92403
rect 635210 92363 635216 92375
rect 661168 92363 661174 92375
rect 661226 92363 661232 92415
rect 634000 92289 634006 92341
rect 634058 92329 634064 92341
rect 660688 92329 660694 92341
rect 634058 92301 660694 92329
rect 634058 92289 634064 92301
rect 660688 92289 660694 92301
rect 660746 92289 660752 92341
rect 640720 92215 640726 92267
rect 640778 92255 640784 92267
rect 661744 92255 661750 92267
rect 640778 92227 661750 92255
rect 640778 92215 640784 92227
rect 661744 92215 661750 92227
rect 661802 92215 661808 92267
rect 152656 92141 152662 92193
rect 152714 92181 152720 92193
rect 198832 92181 198838 92193
rect 152714 92153 198838 92181
rect 152714 92141 152720 92153
rect 198832 92141 198838 92153
rect 198890 92141 198896 92193
rect 640816 92141 640822 92193
rect 640874 92181 640880 92193
rect 657520 92181 657526 92193
rect 640874 92153 657526 92181
rect 640874 92141 640880 92153
rect 657520 92141 657526 92153
rect 657578 92141 657584 92193
rect 151120 92067 151126 92119
rect 151178 92107 151184 92119
rect 198736 92107 198742 92119
rect 151178 92079 198742 92107
rect 151178 92067 151184 92079
rect 198736 92067 198742 92079
rect 198794 92067 198800 92119
rect 156880 91993 156886 92045
rect 156938 92033 156944 92045
rect 199024 92033 199030 92045
rect 156938 92005 199030 92033
rect 156938 91993 156944 92005
rect 199024 91993 199030 92005
rect 199082 91993 199088 92045
rect 188560 91919 188566 91971
rect 188618 91959 188624 91971
rect 199120 91959 199126 91971
rect 188618 91931 199126 91959
rect 188618 91919 188624 91931
rect 199120 91919 199126 91931
rect 199178 91919 199184 91971
rect 185680 91845 185686 91897
rect 185738 91885 185744 91897
rect 198832 91885 198838 91897
rect 185738 91857 198838 91885
rect 185738 91845 185744 91857
rect 198832 91845 198838 91857
rect 198890 91845 198896 91897
rect 182800 91771 182806 91823
rect 182858 91811 182864 91823
rect 198928 91811 198934 91823
rect 182858 91783 198934 91811
rect 182858 91771 182864 91783
rect 198928 91771 198934 91783
rect 198986 91771 198992 91823
rect 144208 90587 144214 90639
rect 144266 90627 144272 90639
rect 160240 90627 160246 90639
rect 144266 90599 160246 90627
rect 144266 90587 144272 90599
rect 160240 90587 160246 90599
rect 160298 90587 160304 90639
rect 144208 89255 144214 89307
rect 144266 89295 144272 89307
rect 163120 89295 163126 89307
rect 144266 89267 163126 89295
rect 144266 89255 144272 89267
rect 163120 89255 163126 89267
rect 163178 89255 163184 89307
rect 168400 89181 168406 89233
rect 168458 89221 168464 89233
rect 198928 89221 198934 89233
rect 168458 89193 198934 89221
rect 168458 89181 168464 89193
rect 198928 89181 198934 89193
rect 198986 89181 198992 89233
rect 174160 89107 174166 89159
rect 174218 89147 174224 89159
rect 199024 89147 199030 89159
rect 174218 89119 199030 89147
rect 174218 89107 174224 89119
rect 199024 89107 199030 89119
rect 199082 89107 199088 89159
rect 177040 89033 177046 89085
rect 177098 89073 177104 89085
rect 198832 89073 198838 89085
rect 177098 89045 198838 89073
rect 177098 89033 177104 89045
rect 198832 89033 198838 89045
rect 198890 89033 198896 89085
rect 179920 88959 179926 89011
rect 179978 88999 179984 89011
rect 198736 88999 198742 89011
rect 179978 88971 198742 88999
rect 179978 88959 179984 88971
rect 198736 88959 198742 88971
rect 198794 88959 198800 89011
rect 194320 88885 194326 88937
rect 194378 88925 194384 88937
rect 199216 88925 199222 88937
rect 194378 88897 199222 88925
rect 194378 88885 194384 88897
rect 199216 88885 199222 88897
rect 199274 88885 199280 88937
rect 635536 87775 635542 87827
rect 635594 87815 635600 87827
rect 652528 87815 652534 87827
rect 635594 87787 652534 87815
rect 635594 87775 635600 87787
rect 652528 87775 652534 87787
rect 652586 87775 652592 87827
rect 144208 87075 144214 87087
rect 144034 87047 144214 87075
rect 144034 86409 144062 87047
rect 144208 87035 144214 87047
rect 144266 87035 144272 87087
rect 144112 86517 144118 86569
rect 144170 86557 144176 86569
rect 163216 86557 163222 86569
rect 144170 86529 163222 86557
rect 144170 86517 144176 86529
rect 163216 86517 163222 86529
rect 163274 86517 163280 86569
rect 202576 86517 202582 86569
rect 202634 86557 202640 86569
rect 204880 86557 204886 86569
rect 202634 86529 204886 86557
rect 202634 86517 202640 86529
rect 204880 86517 204886 86529
rect 204938 86517 204944 86569
rect 144208 86443 144214 86495
rect 144266 86483 144272 86495
rect 202384 86483 202390 86495
rect 144266 86455 202390 86483
rect 144266 86443 144272 86455
rect 202384 86443 202390 86455
rect 202442 86443 202448 86495
rect 640912 86443 640918 86495
rect 640970 86483 640976 86495
rect 652624 86483 652630 86495
rect 640970 86455 652630 86483
rect 640970 86443 640976 86455
rect 652624 86443 652630 86455
rect 652682 86443 652688 86495
rect 144112 86409 144118 86421
rect 144034 86381 144118 86409
rect 144112 86369 144118 86381
rect 144170 86369 144176 86421
rect 151216 86369 151222 86421
rect 151274 86409 151280 86421
rect 199216 86409 199222 86421
rect 151274 86381 199222 86409
rect 151274 86369 151280 86381
rect 199216 86369 199222 86381
rect 199274 86369 199280 86421
rect 200848 86369 200854 86421
rect 200906 86409 200912 86421
rect 201040 86409 201046 86421
rect 200906 86381 201046 86409
rect 200906 86369 200912 86381
rect 201040 86369 201046 86381
rect 201098 86369 201104 86421
rect 154000 86295 154006 86347
rect 154058 86335 154064 86347
rect 199120 86335 199126 86347
rect 154058 86307 199126 86335
rect 154058 86295 154064 86307
rect 199120 86295 199126 86307
rect 199178 86295 199184 86347
rect 202192 86295 202198 86347
rect 202250 86335 202256 86347
rect 202576 86335 202582 86347
rect 202250 86307 202582 86335
rect 202250 86295 202256 86307
rect 202576 86295 202582 86307
rect 202634 86295 202640 86347
rect 159760 86221 159766 86273
rect 159818 86261 159824 86273
rect 198928 86261 198934 86273
rect 159818 86233 198934 86261
rect 159818 86221 159824 86233
rect 198928 86221 198934 86233
rect 198986 86221 198992 86273
rect 162640 86147 162646 86199
rect 162698 86187 162704 86199
rect 199024 86187 199030 86199
rect 162698 86159 199030 86187
rect 162698 86147 162704 86159
rect 199024 86147 199030 86159
rect 199082 86147 199088 86199
rect 165520 86073 165526 86125
rect 165578 86113 165584 86125
rect 198736 86113 198742 86125
rect 165578 86085 198742 86113
rect 165578 86073 165584 86085
rect 198736 86073 198742 86085
rect 198794 86073 198800 86125
rect 171280 85999 171286 86051
rect 171338 86039 171344 86051
rect 198832 86039 198838 86051
rect 171338 86011 198838 86039
rect 171338 85999 171344 86011
rect 198832 85999 198838 86011
rect 198890 85999 198896 86051
rect 146896 83779 146902 83831
rect 146954 83819 146960 83831
rect 163600 83819 163606 83831
rect 146954 83791 163606 83819
rect 146954 83779 146960 83791
rect 163600 83779 163606 83791
rect 163658 83779 163664 83831
rect 641104 83705 641110 83757
rect 641162 83745 641168 83757
rect 653584 83745 653590 83757
rect 641162 83717 653590 83745
rect 641162 83705 641168 83717
rect 653584 83705 653590 83717
rect 653642 83705 653648 83757
rect 144112 83631 144118 83683
rect 144170 83671 144176 83683
rect 163312 83671 163318 83683
rect 144170 83643 163318 83671
rect 144170 83631 144176 83643
rect 163312 83631 163318 83643
rect 163370 83631 163376 83683
rect 635632 83631 635638 83683
rect 635690 83671 635696 83683
rect 653680 83671 653686 83683
rect 635690 83643 653686 83671
rect 635690 83631 635696 83643
rect 653680 83631 653686 83643
rect 653738 83631 653744 83683
rect 635728 83557 635734 83609
rect 635786 83597 635792 83609
rect 653488 83597 653494 83609
rect 635786 83569 653494 83597
rect 635786 83557 635792 83569
rect 653488 83557 653494 83569
rect 653546 83557 653552 83609
rect 146896 83483 146902 83535
rect 146954 83523 146960 83535
rect 148720 83523 148726 83535
rect 146954 83495 148726 83523
rect 146954 83483 146960 83495
rect 148720 83483 148726 83495
rect 148778 83483 148784 83535
rect 197296 83483 197302 83535
rect 197354 83523 197360 83535
rect 200752 83523 200758 83535
rect 197354 83495 200758 83523
rect 197354 83483 197360 83495
rect 200752 83483 200758 83495
rect 200810 83483 200816 83535
rect 194416 83409 194422 83461
rect 194474 83449 194480 83461
rect 199504 83449 199510 83461
rect 194474 83421 199510 83449
rect 194474 83409 194480 83421
rect 199504 83409 199510 83421
rect 199562 83409 199568 83461
rect 191536 83335 191542 83387
rect 191594 83375 191600 83387
rect 198832 83375 198838 83387
rect 191594 83347 198838 83375
rect 191594 83335 191600 83347
rect 198832 83335 198838 83347
rect 198890 83335 198896 83387
rect 188656 83261 188662 83313
rect 188714 83301 188720 83313
rect 198928 83301 198934 83313
rect 188714 83273 198934 83301
rect 188714 83261 188720 83273
rect 198928 83261 198934 83273
rect 198986 83261 198992 83313
rect 156976 83187 156982 83239
rect 157034 83227 157040 83239
rect 198736 83227 198742 83239
rect 157034 83199 198742 83227
rect 157034 83187 157040 83199
rect 198736 83187 198742 83199
rect 198794 83187 198800 83239
rect 146992 82151 146998 82203
rect 147050 82191 147056 82203
rect 160048 82191 160054 82203
rect 147050 82163 160054 82191
rect 147050 82151 147056 82163
rect 160048 82151 160054 82163
rect 160106 82151 160112 82203
rect 640624 81041 640630 81093
rect 640682 81081 640688 81093
rect 663280 81081 663286 81093
rect 640682 81053 663286 81081
rect 640682 81041 640688 81053
rect 663280 81041 663286 81053
rect 663338 81041 663344 81093
rect 641296 80893 641302 80945
rect 641354 80933 641360 80945
rect 663472 80933 663478 80945
rect 641354 80905 663478 80933
rect 641354 80893 641360 80905
rect 663472 80893 663478 80905
rect 663530 80893 663536 80945
rect 662416 80859 662422 80871
rect 641122 80831 662422 80859
rect 635920 80745 635926 80797
rect 635978 80785 635984 80797
rect 641122 80785 641150 80831
rect 662416 80819 662422 80831
rect 662474 80819 662480 80871
rect 635978 80757 641150 80785
rect 635978 80745 635984 80757
rect 641200 80745 641206 80797
rect 641258 80785 641264 80797
rect 653680 80785 653686 80797
rect 641258 80757 653686 80785
rect 641258 80745 641264 80757
rect 653680 80745 653686 80757
rect 653738 80745 653744 80797
rect 144112 80671 144118 80723
rect 144170 80711 144176 80723
rect 162640 80711 162646 80723
rect 144170 80683 162646 80711
rect 144170 80671 144176 80683
rect 162640 80671 162646 80683
rect 162698 80671 162704 80723
rect 201808 80671 201814 80723
rect 201866 80711 201872 80723
rect 202096 80711 202102 80723
rect 201866 80683 202102 80711
rect 201866 80671 201872 80683
rect 202096 80671 202102 80683
rect 202154 80671 202160 80723
rect 635824 80671 635830 80723
rect 635882 80711 635888 80723
rect 640624 80711 640630 80723
rect 635882 80683 640630 80711
rect 635882 80671 635888 80683
rect 640624 80671 640630 80683
rect 640682 80671 640688 80723
rect 641392 80671 641398 80723
rect 641450 80711 641456 80723
rect 653584 80711 653590 80723
rect 641450 80683 653590 80711
rect 641450 80671 641456 80683
rect 653584 80671 653590 80683
rect 653642 80671 653648 80723
rect 168496 80597 168502 80649
rect 168554 80637 168560 80649
rect 198928 80637 198934 80649
rect 168554 80609 198934 80637
rect 168554 80597 168560 80609
rect 198928 80597 198934 80609
rect 198986 80597 198992 80649
rect 177136 80523 177142 80575
rect 177194 80563 177200 80575
rect 199024 80563 199030 80575
rect 177194 80535 199030 80563
rect 177194 80523 177200 80535
rect 199024 80523 199030 80535
rect 199082 80523 199088 80575
rect 180016 80449 180022 80501
rect 180074 80489 180080 80501
rect 198832 80489 198838 80501
rect 180074 80461 198838 80489
rect 180074 80449 180080 80461
rect 198832 80449 198838 80461
rect 198890 80449 198896 80501
rect 185776 80375 185782 80427
rect 185834 80415 185840 80427
rect 198736 80415 198742 80427
rect 185834 80387 198742 80415
rect 185834 80375 185840 80387
rect 198736 80375 198742 80387
rect 198794 80375 198800 80427
rect 182896 80227 182902 80279
rect 182954 80267 182960 80279
rect 198736 80267 198742 80279
rect 182954 80239 198742 80267
rect 182954 80227 182960 80239
rect 198736 80227 198742 80239
rect 198794 80227 198800 80279
rect 144208 78639 144214 78651
rect 144034 78611 144214 78639
rect 144034 77751 144062 78611
rect 144208 78599 144214 78611
rect 144266 78599 144272 78651
rect 144112 77859 144118 77911
rect 144170 77899 144176 77911
rect 163408 77899 163414 77911
rect 144170 77871 163414 77899
rect 144170 77859 144176 77871
rect 163408 77859 163414 77871
rect 163466 77859 163472 77911
rect 144208 77785 144214 77837
rect 144266 77825 144272 77837
rect 163504 77825 163510 77837
rect 144266 77797 163510 77825
rect 144266 77785 144272 77797
rect 163504 77785 163510 77797
rect 163562 77785 163568 77837
rect 144112 77751 144118 77763
rect 144034 77723 144118 77751
rect 144112 77711 144118 77723
rect 144170 77711 144176 77763
rect 149104 77711 149110 77763
rect 149162 77751 149168 77763
rect 199120 77751 199126 77763
rect 149162 77723 199126 77751
rect 149162 77711 149168 77723
rect 199120 77711 199126 77723
rect 199178 77711 199184 77763
rect 641488 77711 641494 77763
rect 641546 77751 641552 77763
rect 657520 77751 657526 77763
rect 641546 77723 657526 77751
rect 641546 77711 641552 77723
rect 657520 77711 657526 77723
rect 657578 77711 657584 77763
rect 149008 77637 149014 77689
rect 149066 77677 149072 77689
rect 198736 77677 198742 77689
rect 149066 77649 198742 77677
rect 149066 77637 149072 77649
rect 198736 77637 198742 77649
rect 198794 77637 198800 77689
rect 642160 77637 642166 77689
rect 642218 77677 642224 77689
rect 663760 77677 663766 77689
rect 642218 77649 663766 77677
rect 642218 77637 642224 77649
rect 663760 77637 663766 77649
rect 663818 77637 663824 77689
rect 149776 77563 149782 77615
rect 149834 77603 149840 77615
rect 198928 77603 198934 77615
rect 149834 77575 198934 77603
rect 149834 77563 149840 77575
rect 198928 77563 198934 77575
rect 198986 77563 198992 77615
rect 165616 77489 165622 77541
rect 165674 77529 165680 77541
rect 199024 77529 199030 77541
rect 165674 77501 199030 77529
rect 165674 77489 165680 77501
rect 199024 77489 199030 77501
rect 199082 77489 199088 77541
rect 171376 77415 171382 77467
rect 171434 77455 171440 77467
rect 198832 77455 198838 77467
rect 171434 77427 198838 77455
rect 171434 77415 171440 77427
rect 198832 77415 198838 77427
rect 198890 77415 198896 77467
rect 174256 77341 174262 77393
rect 174314 77381 174320 77393
rect 198736 77381 198742 77393
rect 174314 77353 198742 77381
rect 174314 77341 174320 77353
rect 198736 77341 198742 77353
rect 198794 77341 198800 77393
rect 144208 77267 144214 77319
rect 144266 77307 144272 77319
rect 155536 77307 155542 77319
rect 144266 77279 155542 77307
rect 144266 77267 144272 77279
rect 155536 77267 155542 77279
rect 155594 77267 155600 77319
rect 641584 76897 641590 76949
rect 641642 76937 641648 76949
rect 659632 76937 659638 76949
rect 641642 76909 659638 76937
rect 641642 76897 641648 76909
rect 659632 76897 659638 76909
rect 659690 76897 659696 76949
rect 658288 76863 658294 76875
rect 640162 76835 658294 76863
rect 636304 76749 636310 76801
rect 636362 76789 636368 76801
rect 640162 76789 640190 76835
rect 658288 76823 658294 76835
rect 658346 76823 658352 76875
rect 636362 76761 640190 76789
rect 636362 76749 636368 76761
rect 641680 76749 641686 76801
rect 641738 76789 641744 76801
rect 658864 76789 658870 76801
rect 641738 76761 658870 76789
rect 641738 76749 641744 76761
rect 658864 76749 658870 76761
rect 658922 76749 658928 76801
rect 636016 76675 636022 76727
rect 636074 76715 636080 76727
rect 656944 76715 656950 76727
rect 636074 76687 656950 76715
rect 636074 76675 636080 76687
rect 656944 76675 656950 76687
rect 657002 76675 657008 76727
rect 636208 76601 636214 76653
rect 636266 76641 636272 76653
rect 660688 76641 660694 76653
rect 636266 76613 660694 76641
rect 636266 76601 636272 76613
rect 660688 76601 660694 76613
rect 660746 76601 660752 76653
rect 636112 76527 636118 76579
rect 636170 76567 636176 76579
rect 661168 76567 661174 76579
rect 636170 76539 661174 76567
rect 636170 76527 636176 76539
rect 661168 76527 661174 76539
rect 661226 76527 661232 76579
rect 634768 76453 634774 76505
rect 634826 76493 634832 76505
rect 661744 76493 661750 76505
rect 634826 76465 661750 76493
rect 634826 76453 634832 76465
rect 661744 76453 661750 76465
rect 661802 76453 661808 76505
rect 634864 76379 634870 76431
rect 634922 76419 634928 76431
rect 660112 76419 660118 76431
rect 634922 76391 660118 76419
rect 634922 76379 634928 76391
rect 660112 76379 660118 76391
rect 660170 76379 660176 76431
rect 636400 76305 636406 76357
rect 636458 76345 636464 76357
rect 662512 76345 662518 76357
rect 636458 76317 662518 76345
rect 636458 76305 636464 76317
rect 662512 76305 662518 76317
rect 662570 76305 662576 76357
rect 144208 75343 144214 75395
rect 144266 75383 144272 75395
rect 159760 75383 159766 75395
rect 144266 75355 159766 75383
rect 144266 75343 144272 75355
rect 159760 75343 159766 75355
rect 159818 75343 159824 75395
rect 144016 75195 144022 75247
rect 144074 75235 144080 75247
rect 144208 75235 144214 75247
rect 144074 75207 144214 75235
rect 144074 75195 144080 75207
rect 144208 75195 144214 75207
rect 144266 75195 144272 75247
rect 143920 74973 143926 75025
rect 143978 75013 143984 75025
rect 144112 75013 144118 75025
rect 143978 74985 144118 75013
rect 143978 74973 143984 74985
rect 144112 74973 144118 74985
rect 144170 74973 144176 75025
rect 146896 74899 146902 74951
rect 146954 74939 146960 74951
rect 151120 74939 151126 74951
rect 146954 74911 151126 74939
rect 146954 74899 146960 74911
rect 151120 74899 151126 74911
rect 151178 74899 151184 74951
rect 154096 74825 154102 74877
rect 154154 74865 154160 74877
rect 198928 74865 198934 74877
rect 154154 74837 198934 74865
rect 154154 74825 154160 74837
rect 198928 74825 198934 74837
rect 198986 74825 198992 74877
rect 157072 74751 157078 74803
rect 157130 74791 157136 74803
rect 199120 74791 199126 74803
rect 157130 74763 199126 74791
rect 157130 74751 157136 74763
rect 199120 74751 199126 74763
rect 199178 74751 199184 74803
rect 160240 74677 160246 74729
rect 160298 74717 160304 74729
rect 199024 74717 199030 74729
rect 160298 74689 199030 74717
rect 160298 74677 160304 74689
rect 199024 74677 199030 74689
rect 199082 74677 199088 74729
rect 159856 74603 159862 74655
rect 159914 74643 159920 74655
rect 198736 74643 198742 74655
rect 159914 74615 198742 74643
rect 159914 74603 159920 74615
rect 198736 74603 198742 74615
rect 198794 74603 198800 74655
rect 163024 74529 163030 74581
rect 163082 74569 163088 74581
rect 198832 74569 198838 74581
rect 163082 74541 198838 74569
rect 163082 74529 163088 74541
rect 198832 74529 198838 74541
rect 198890 74529 198896 74581
rect 143920 73715 143926 73767
rect 143978 73755 143984 73767
rect 159952 73755 159958 73767
rect 143978 73727 159958 73755
rect 143978 73715 143984 73727
rect 159952 73715 159958 73727
rect 160010 73715 160016 73767
rect 143920 72013 143926 72065
rect 143978 72053 143984 72065
rect 160144 72053 160150 72065
rect 143978 72025 160150 72053
rect 143978 72013 143984 72025
rect 160144 72013 160150 72025
rect 160202 72013 160208 72065
rect 197392 71939 197398 71991
rect 197450 71979 197456 71991
rect 200752 71979 200758 71991
rect 197450 71951 200758 71979
rect 197450 71939 197456 71951
rect 200752 71939 200758 71951
rect 200810 71939 200816 71991
rect 194512 71865 194518 71917
rect 194570 71905 194576 71917
rect 199600 71905 199606 71917
rect 194570 71877 199606 71905
rect 194570 71865 194576 71877
rect 199600 71865 199606 71877
rect 199658 71865 199664 71917
rect 191632 71791 191638 71843
rect 191690 71831 191696 71843
rect 198832 71831 198838 71843
rect 191690 71803 198838 71831
rect 191690 71791 191696 71803
rect 198832 71791 198838 71803
rect 198890 71791 198896 71843
rect 188752 71717 188758 71769
rect 188810 71757 188816 71769
rect 198928 71757 198934 71769
rect 188810 71729 198934 71757
rect 188810 71717 188816 71729
rect 198928 71717 198934 71729
rect 198986 71717 198992 71769
rect 151312 71643 151318 71695
rect 151370 71683 151376 71695
rect 198736 71683 198742 71695
rect 151370 71655 198742 71683
rect 151370 71643 151376 71655
rect 198736 71643 198742 71655
rect 198794 71643 198800 71695
rect 146896 70015 146902 70067
rect 146954 70055 146960 70067
rect 159856 70055 159862 70067
rect 146954 70027 159862 70055
rect 146954 70015 146960 70027
rect 159856 70015 159862 70027
rect 159914 70015 159920 70067
rect 147472 69053 147478 69105
rect 147530 69093 147536 69105
rect 199024 69093 199030 69105
rect 147530 69065 199030 69093
rect 147530 69053 147536 69065
rect 199024 69053 199030 69065
rect 199082 69053 199088 69105
rect 168592 68979 168598 69031
rect 168650 69019 168656 69031
rect 199120 69019 199126 69031
rect 168650 68991 199126 69019
rect 168650 68979 168656 68991
rect 199120 68979 199126 68991
rect 199178 68979 199184 69031
rect 180112 68905 180118 68957
rect 180170 68945 180176 68957
rect 198928 68945 198934 68957
rect 180170 68917 198934 68945
rect 180170 68905 180176 68917
rect 198928 68905 198934 68917
rect 198986 68905 198992 68957
rect 185872 68831 185878 68883
rect 185930 68871 185936 68883
rect 198832 68871 198838 68883
rect 185930 68843 198838 68871
rect 185930 68831 185936 68843
rect 198832 68831 198838 68843
rect 198890 68831 198896 68883
rect 182992 68757 182998 68809
rect 183050 68797 183056 68809
rect 198736 68797 198742 68809
rect 183050 68769 198742 68797
rect 183050 68757 183056 68769
rect 198736 68757 198742 68769
rect 198794 68757 198800 68809
rect 143920 66907 143926 66959
rect 143978 66947 143984 66959
rect 160240 66947 160246 66959
rect 143978 66919 160246 66947
rect 143978 66907 143984 66919
rect 160240 66907 160246 66919
rect 160298 66907 160304 66959
rect 143920 66759 143926 66811
rect 143978 66799 143984 66811
rect 160336 66799 160342 66811
rect 143978 66771 160342 66799
rect 143978 66759 143984 66771
rect 160336 66759 160342 66771
rect 160394 66759 160400 66811
rect 200848 66315 200854 66367
rect 200906 66355 200912 66367
rect 200906 66327 201086 66355
rect 200906 66315 200912 66327
rect 201058 66293 201086 66327
rect 143824 66241 143830 66293
rect 143882 66281 143888 66293
rect 167056 66281 167062 66293
rect 143882 66253 167062 66281
rect 143882 66241 143888 66253
rect 167056 66241 167062 66253
rect 167114 66241 167120 66293
rect 201040 66241 201046 66293
rect 201098 66241 201104 66293
rect 147376 66167 147382 66219
rect 147434 66207 147440 66219
rect 199120 66207 199126 66219
rect 147434 66179 199126 66207
rect 147434 66167 147440 66179
rect 199120 66167 199126 66179
rect 199178 66167 199184 66219
rect 147280 66093 147286 66145
rect 147338 66133 147344 66145
rect 199216 66133 199222 66145
rect 147338 66105 199222 66133
rect 147338 66093 147344 66105
rect 199216 66093 199222 66105
rect 199274 66093 199280 66145
rect 165712 66019 165718 66071
rect 165770 66059 165776 66071
rect 199024 66059 199030 66071
rect 165770 66031 199030 66059
rect 165770 66019 165776 66031
rect 199024 66019 199030 66031
rect 199082 66019 199088 66071
rect 171472 65945 171478 65997
rect 171530 65985 171536 65997
rect 198832 65985 198838 65997
rect 171530 65957 198838 65985
rect 171530 65945 171536 65957
rect 198832 65945 198838 65957
rect 198890 65945 198896 65997
rect 174352 65871 174358 65923
rect 174410 65911 174416 65923
rect 198736 65911 198742 65923
rect 174410 65883 198742 65911
rect 174410 65871 174416 65883
rect 198736 65871 198742 65883
rect 198794 65871 198800 65923
rect 177232 65797 177238 65849
rect 177290 65837 177296 65849
rect 198928 65837 198934 65849
rect 177290 65809 198934 65837
rect 177290 65797 177296 65809
rect 198928 65797 198934 65809
rect 198986 65797 198992 65849
rect 152656 65353 152662 65405
rect 152714 65393 152720 65405
rect 155152 65393 155158 65405
rect 152714 65365 155158 65393
rect 152714 65353 152720 65365
rect 155152 65353 155158 65365
rect 155210 65353 155216 65405
rect 146896 64095 146902 64147
rect 146954 64135 146960 64147
rect 160432 64135 160438 64147
rect 146954 64107 160438 64135
rect 146954 64095 146960 64107
rect 160432 64095 160438 64107
rect 160490 64095 160496 64147
rect 143920 63355 143926 63407
rect 143978 63395 143984 63407
rect 164272 63395 164278 63407
rect 143978 63367 164278 63395
rect 143978 63355 143984 63367
rect 164272 63355 164278 63367
rect 164330 63355 164336 63407
rect 146992 63281 146998 63333
rect 147050 63321 147056 63333
rect 199120 63321 199126 63333
rect 147050 63293 199126 63321
rect 147050 63281 147056 63293
rect 199120 63281 199126 63293
rect 199178 63281 199184 63333
rect 151120 63207 151126 63259
rect 151178 63247 151184 63259
rect 199024 63247 199030 63259
rect 151178 63219 199030 63247
rect 151178 63207 151184 63219
rect 199024 63207 199030 63219
rect 199082 63207 199088 63259
rect 155536 63133 155542 63185
rect 155594 63173 155600 63185
rect 198928 63173 198934 63185
rect 155594 63145 198934 63173
rect 155594 63133 155600 63145
rect 198928 63133 198934 63145
rect 198986 63133 198992 63185
rect 160048 63059 160054 63111
rect 160106 63099 160112 63111
rect 198832 63099 198838 63111
rect 160106 63071 198838 63099
rect 160106 63059 160112 63071
rect 198832 63059 198838 63071
rect 198890 63059 198896 63111
rect 163600 62985 163606 63037
rect 163658 63025 163664 63037
rect 198736 63025 198742 63037
rect 163658 62997 198742 63025
rect 163658 62985 163664 62997
rect 198736 62985 198742 62997
rect 198794 62985 198800 63037
rect 202000 61505 202006 61557
rect 202058 61545 202064 61557
rect 203056 61545 203062 61557
rect 202058 61517 203062 61545
rect 202058 61505 202064 61517
rect 203056 61505 203062 61517
rect 203114 61505 203120 61557
rect 202288 61431 202294 61483
rect 202346 61471 202352 61483
rect 202960 61471 202966 61483
rect 202346 61443 202966 61471
rect 202346 61431 202352 61443
rect 202960 61431 202966 61443
rect 203018 61431 203024 61483
rect 202192 61357 202198 61409
rect 202250 61397 202256 61409
rect 203344 61397 203350 61409
rect 202250 61369 203350 61397
rect 202250 61357 202256 61369
rect 203344 61357 203350 61369
rect 203402 61357 203408 61409
rect 202480 61283 202486 61335
rect 202538 61323 202544 61335
rect 203248 61323 203254 61335
rect 202538 61295 203254 61323
rect 202538 61283 202544 61295
rect 203248 61283 203254 61295
rect 203306 61283 203312 61335
rect 203248 60839 203254 60891
rect 203306 60879 203312 60891
rect 203728 60879 203734 60891
rect 203306 60851 203734 60879
rect 203306 60839 203312 60851
rect 203728 60839 203734 60851
rect 203786 60839 203792 60891
rect 146896 60617 146902 60669
rect 146954 60657 146960 60669
rect 160528 60657 160534 60669
rect 146954 60629 160534 60657
rect 146954 60617 146960 60629
rect 160528 60617 160534 60629
rect 160586 60617 160592 60669
rect 146992 60543 146998 60595
rect 147050 60583 147056 60595
rect 147050 60555 164126 60583
rect 147050 60543 147056 60555
rect 138160 60469 138166 60521
rect 138218 60509 138224 60521
rect 159088 60509 159094 60521
rect 138218 60481 159094 60509
rect 138218 60469 138224 60481
rect 159088 60469 159094 60481
rect 159146 60469 159152 60521
rect 164098 60435 164126 60555
rect 198928 60435 198934 60447
rect 164098 60407 198934 60435
rect 198928 60395 198934 60407
rect 198986 60395 198992 60447
rect 640144 60395 640150 60447
rect 640202 60435 640208 60447
rect 663568 60435 663574 60447
rect 640202 60407 663574 60435
rect 640202 60395 640208 60407
rect 663568 60395 663574 60407
rect 663626 60395 663632 60447
rect 164272 60321 164278 60373
rect 164330 60361 164336 60373
rect 198832 60361 198838 60373
rect 164330 60333 198838 60361
rect 164330 60321 164336 60333
rect 198832 60321 198838 60333
rect 198890 60321 198896 60373
rect 167056 60247 167062 60299
rect 167114 60287 167120 60299
rect 198736 60287 198742 60299
rect 167114 60259 198742 60287
rect 167114 60247 167120 60259
rect 198736 60247 198742 60259
rect 198794 60247 198800 60299
rect 204016 59063 204022 59115
rect 204074 59103 204080 59115
rect 204976 59103 204982 59115
rect 204074 59075 204982 59103
rect 204074 59063 204080 59075
rect 204976 59063 204982 59075
rect 205034 59063 205040 59115
rect 204784 58915 204790 58967
rect 204842 58955 204848 58967
rect 204976 58955 204982 58967
rect 204842 58927 204982 58955
rect 204842 58915 204848 58927
rect 204976 58915 204982 58927
rect 205034 58915 205040 58967
rect 204112 57287 204118 57339
rect 204170 57327 204176 57339
rect 204496 57327 204502 57339
rect 204170 57299 204502 57327
rect 204170 57287 204176 57299
rect 204496 57287 204502 57299
rect 204554 57287 204560 57339
rect 204208 56251 204214 56303
rect 204266 56291 204272 56303
rect 204688 56291 204694 56303
rect 204266 56263 204694 56291
rect 204266 56251 204272 56263
rect 204688 56251 204694 56263
rect 204746 56251 204752 56303
rect 204976 54771 204982 54823
rect 205034 54771 205040 54823
rect 204994 54219 205022 54771
rect 639568 54623 639574 54675
rect 639626 54663 639632 54675
rect 639952 54663 639958 54675
rect 639626 54635 639958 54663
rect 639626 54623 639632 54635
rect 639952 54623 639958 54635
rect 640010 54623 640016 54675
rect 205936 54219 205942 54231
rect 204994 54191 205942 54219
rect 205936 54179 205942 54191
rect 205994 54179 206000 54231
rect 215152 54219 215158 54231
rect 206050 54191 215158 54219
rect 201040 54105 201046 54157
rect 201098 54145 201104 54157
rect 206050 54145 206078 54191
rect 215152 54179 215158 54191
rect 215210 54179 215216 54231
rect 632272 54179 632278 54231
rect 632330 54219 632336 54231
rect 634960 54219 634966 54231
rect 632330 54191 634966 54219
rect 632330 54179 632336 54191
rect 634960 54179 634966 54191
rect 635018 54179 635024 54231
rect 201098 54117 206078 54145
rect 201098 54105 201104 54117
rect 206320 54105 206326 54157
rect 206378 54145 206384 54157
rect 214960 54145 214966 54157
rect 206378 54117 214966 54145
rect 206378 54105 206384 54117
rect 214960 54105 214966 54117
rect 215018 54105 215024 54157
rect 633712 54105 633718 54157
rect 633770 54145 633776 54157
rect 636208 54145 636214 54157
rect 633770 54117 636214 54145
rect 633770 54105 633776 54117
rect 636208 54105 636214 54117
rect 636266 54105 636272 54157
rect 200656 54031 200662 54083
rect 200714 54071 200720 54083
rect 214768 54071 214774 54083
rect 200714 54043 214774 54071
rect 200714 54031 200720 54043
rect 214768 54031 214774 54043
rect 214826 54031 214832 54083
rect 633328 54031 633334 54083
rect 633386 54071 633392 54083
rect 636016 54071 636022 54083
rect 633386 54043 636022 54071
rect 633386 54031 633392 54043
rect 636016 54031 636022 54043
rect 636074 54031 636080 54083
rect 201136 53957 201142 54009
rect 201194 53997 201200 54009
rect 201194 53969 206462 53997
rect 201194 53957 201200 53969
rect 204976 53883 204982 53935
rect 205034 53923 205040 53935
rect 206128 53923 206134 53935
rect 205034 53895 206134 53923
rect 205034 53883 205040 53895
rect 206128 53883 206134 53895
rect 206186 53883 206192 53935
rect 199696 53809 199702 53861
rect 199754 53849 199760 53861
rect 206320 53849 206326 53861
rect 199754 53821 206326 53849
rect 199754 53809 199760 53821
rect 206320 53809 206326 53821
rect 206378 53809 206384 53861
rect 206434 53849 206462 53969
rect 632560 53957 632566 54009
rect 632618 53997 632624 54009
rect 635824 53997 635830 54009
rect 632618 53969 635830 53997
rect 632618 53957 632624 53969
rect 635824 53957 635830 53969
rect 635882 53957 635888 54009
rect 631888 53883 631894 53935
rect 631946 53923 631952 53935
rect 635440 53923 635446 53935
rect 631946 53895 635446 53923
rect 631946 53883 631952 53895
rect 635440 53883 635446 53895
rect 635498 53883 635504 53935
rect 206434 53821 214190 53849
rect 201424 53735 201430 53787
rect 201482 53775 201488 53787
rect 201482 53747 213470 53775
rect 201482 53735 201488 53747
rect 201232 53661 201238 53713
rect 201290 53701 201296 53713
rect 201290 53673 211982 53701
rect 201290 53661 201296 53673
rect 211954 53639 211982 53673
rect 213442 53639 213470 53747
rect 214162 53639 214190 53821
rect 629296 53809 629302 53861
rect 629354 53849 629360 53861
rect 634768 53849 634774 53861
rect 629354 53821 634774 53849
rect 629354 53809 629360 53821
rect 634768 53809 634774 53821
rect 634826 53809 634832 53861
rect 630352 53735 630358 53787
rect 630410 53775 630416 53787
rect 635248 53775 635254 53787
rect 630410 53747 635254 53775
rect 630410 53735 630416 53747
rect 635248 53735 635254 53747
rect 635306 53735 635312 53787
rect 630064 53661 630070 53713
rect 630122 53701 630128 53713
rect 635152 53701 635158 53713
rect 630122 53673 635158 53701
rect 630122 53661 630128 53673
rect 635152 53661 635158 53673
rect 635210 53661 635216 53713
rect 204304 53587 204310 53639
rect 204362 53627 204368 53639
rect 207472 53627 207478 53639
rect 204362 53599 207478 53627
rect 204362 53587 204368 53599
rect 207472 53587 207478 53599
rect 207530 53587 207536 53639
rect 207568 53587 207574 53639
rect 207626 53627 207632 53639
rect 209728 53627 209734 53639
rect 207626 53599 209734 53627
rect 207626 53587 207632 53599
rect 209728 53587 209734 53599
rect 209786 53587 209792 53639
rect 210736 53587 210742 53639
rect 210794 53627 210800 53639
rect 211552 53627 211558 53639
rect 210794 53599 211558 53627
rect 210794 53587 210800 53599
rect 211552 53587 211558 53599
rect 211610 53587 211616 53639
rect 211936 53587 211942 53639
rect 211994 53587 212000 53639
rect 213424 53587 213430 53639
rect 213482 53587 213488 53639
rect 214144 53587 214150 53639
rect 214202 53587 214208 53639
rect 214768 53587 214774 53639
rect 214826 53627 214832 53639
rect 215632 53627 215638 53639
rect 214826 53599 215638 53627
rect 214826 53587 214832 53599
rect 215632 53587 215638 53599
rect 215690 53587 215696 53639
rect 631504 53587 631510 53639
rect 631562 53627 631568 53639
rect 635632 53627 635638 53639
rect 631562 53599 635638 53627
rect 631562 53587 631568 53599
rect 635632 53587 635638 53599
rect 635690 53587 635696 53639
rect 199792 53513 199798 53565
rect 199850 53553 199856 53565
rect 210064 53553 210070 53565
rect 199850 53525 210070 53553
rect 199850 53513 199856 53525
rect 210064 53513 210070 53525
rect 210122 53513 210128 53565
rect 631120 53513 631126 53565
rect 631178 53553 631184 53565
rect 635920 53553 635926 53565
rect 631178 53525 635926 53553
rect 631178 53513 631184 53525
rect 635920 53513 635926 53525
rect 635978 53513 635984 53565
rect 163504 53439 163510 53491
rect 163562 53479 163568 53491
rect 212848 53479 212854 53491
rect 163562 53451 212854 53479
rect 163562 53439 163568 53451
rect 212848 53439 212854 53451
rect 212906 53439 212912 53491
rect 627760 53439 627766 53491
rect 627818 53479 627824 53491
rect 635728 53479 635734 53491
rect 627818 53451 635734 53479
rect 627818 53439 627824 53451
rect 635728 53439 635734 53451
rect 635786 53439 635792 53491
rect 202096 53365 202102 53417
rect 202154 53405 202160 53417
rect 204304 53405 204310 53417
rect 202154 53377 204310 53405
rect 202154 53365 202160 53377
rect 204304 53365 204310 53377
rect 204362 53365 204368 53417
rect 204496 53365 204502 53417
rect 204554 53405 204560 53417
rect 206320 53405 206326 53417
rect 204554 53377 206326 53405
rect 204554 53365 204560 53377
rect 206320 53365 206326 53377
rect 206378 53365 206384 53417
rect 206512 53365 206518 53417
rect 206570 53405 206576 53417
rect 211216 53405 211222 53417
rect 206570 53377 211222 53405
rect 206570 53365 206576 53377
rect 211216 53365 211222 53377
rect 211274 53365 211280 53417
rect 160432 53291 160438 53343
rect 160490 53331 160496 53343
rect 210256 53331 210262 53343
rect 160490 53303 210262 53331
rect 160490 53291 160496 53303
rect 210256 53291 210262 53303
rect 210314 53291 210320 53343
rect 204112 53217 204118 53269
rect 204170 53257 204176 53269
rect 204496 53257 204502 53269
rect 204170 53229 204502 53257
rect 204170 53217 204176 53229
rect 204496 53217 204502 53229
rect 204554 53217 204560 53269
rect 204592 53217 204598 53269
rect 204650 53257 204656 53269
rect 205552 53257 205558 53269
rect 204650 53229 205558 53257
rect 204650 53217 204656 53229
rect 205552 53217 205558 53229
rect 205610 53217 205616 53269
rect 206896 53217 206902 53269
rect 206954 53257 206960 53269
rect 215824 53257 215830 53269
rect 206954 53229 215830 53257
rect 206954 53217 206960 53229
rect 215824 53217 215830 53229
rect 215882 53217 215888 53269
rect 160336 53143 160342 53195
rect 160394 53183 160400 53195
rect 210640 53183 210646 53195
rect 160394 53155 210646 53183
rect 160394 53143 160400 53155
rect 210640 53143 210646 53155
rect 210698 53143 210704 53195
rect 204400 53069 204406 53121
rect 204458 53109 204464 53121
rect 205264 53109 205270 53121
rect 204458 53081 205270 53109
rect 204458 53069 204464 53081
rect 205264 53069 205270 53081
rect 205322 53069 205328 53121
rect 205840 53069 205846 53121
rect 205898 53109 205904 53121
rect 227920 53109 227926 53121
rect 205898 53081 227926 53109
rect 205898 53069 205904 53081
rect 227920 53069 227926 53081
rect 227978 53069 227984 53121
rect 160240 52995 160246 53047
rect 160298 53035 160304 53047
rect 211024 53035 211030 53047
rect 160298 53007 211030 53035
rect 160298 52995 160304 53007
rect 211024 52995 211030 53007
rect 211082 52995 211088 53047
rect 163408 52921 163414 52973
rect 163466 52961 163472 52973
rect 213232 52961 213238 52973
rect 163466 52933 213238 52961
rect 163466 52921 163472 52933
rect 213232 52921 213238 52933
rect 213290 52921 213296 52973
rect 160144 52847 160150 52899
rect 160202 52887 160208 52899
rect 211696 52887 211702 52899
rect 160202 52859 211702 52887
rect 160202 52847 160208 52859
rect 211696 52847 211702 52859
rect 211754 52847 211760 52899
rect 163312 52773 163318 52825
rect 163370 52813 163376 52825
rect 213904 52813 213910 52825
rect 163370 52785 213910 52813
rect 163370 52773 163376 52785
rect 213904 52773 213910 52785
rect 213962 52773 213968 52825
rect 159952 52699 159958 52751
rect 160010 52739 160016 52751
rect 212080 52739 212086 52751
rect 160010 52711 212086 52739
rect 160010 52699 160016 52711
rect 212080 52699 212086 52711
rect 212138 52699 212144 52751
rect 160528 52625 160534 52677
rect 160586 52665 160592 52677
rect 209872 52665 209878 52677
rect 160586 52637 209878 52665
rect 160586 52625 160592 52637
rect 209872 52625 209878 52637
rect 209930 52625 209936 52677
rect 159952 52551 159958 52603
rect 160010 52591 160016 52603
rect 211408 52591 211414 52603
rect 160010 52563 211414 52591
rect 160010 52551 160016 52563
rect 211408 52551 211414 52563
rect 211466 52551 211472 52603
rect 162640 52477 162646 52529
rect 162698 52517 162704 52529
rect 213616 52517 213622 52529
rect 162698 52489 213622 52517
rect 162698 52477 162704 52489
rect 213616 52477 213622 52489
rect 213674 52477 213680 52529
rect 162928 52403 162934 52455
rect 162986 52443 162992 52455
rect 222544 52443 222550 52455
rect 162986 52415 222550 52443
rect 162986 52403 162992 52415
rect 222544 52403 222550 52415
rect 222602 52403 222608 52455
rect 163216 52329 163222 52381
rect 163274 52369 163280 52381
rect 218704 52369 218710 52381
rect 163274 52341 218710 52369
rect 163274 52329 163280 52341
rect 218704 52329 218710 52341
rect 218762 52329 218768 52381
rect 162832 52255 162838 52307
rect 162890 52295 162896 52307
rect 223504 52295 223510 52307
rect 162890 52267 223510 52295
rect 162890 52255 162896 52267
rect 223504 52255 223510 52267
rect 223562 52255 223568 52307
rect 163120 52181 163126 52233
rect 163178 52221 163184 52233
rect 221296 52221 221302 52233
rect 163178 52193 221302 52221
rect 163178 52181 163184 52193
rect 221296 52181 221302 52193
rect 221354 52181 221360 52233
rect 162736 52107 162742 52159
rect 162794 52147 162800 52159
rect 224272 52147 224278 52159
rect 162794 52119 224278 52147
rect 162794 52107 162800 52119
rect 224272 52107 224278 52119
rect 224330 52107 224336 52159
rect 204688 52033 204694 52085
rect 204746 52073 204752 52085
rect 205168 52073 205174 52085
rect 204746 52045 205174 52073
rect 204746 52033 204752 52045
rect 205168 52033 205174 52045
rect 205226 52033 205232 52085
rect 205360 52033 205366 52085
rect 205418 52073 205424 52085
rect 634096 52073 634102 52085
rect 205418 52045 634102 52073
rect 205418 52033 205424 52045
rect 634096 52033 634102 52045
rect 634154 52033 634160 52085
rect 159952 51959 159958 52011
rect 160010 51999 160016 52011
rect 212464 51999 212470 52011
rect 160010 51971 212470 51999
rect 160010 51959 160016 51971
rect 212464 51959 212470 51971
rect 212522 51959 212528 52011
rect 212656 51959 212662 52011
rect 212714 51999 212720 52011
rect 639760 51999 639766 52011
rect 212714 51971 639766 51999
rect 212714 51959 212720 51971
rect 639760 51959 639766 51971
rect 639818 51959 639824 52011
rect 204784 51885 204790 51937
rect 204842 51925 204848 51937
rect 205072 51925 205078 51937
rect 204842 51897 205078 51925
rect 204842 51885 204848 51897
rect 205072 51885 205078 51897
rect 205130 51885 205136 51937
rect 206032 51885 206038 51937
rect 206090 51925 206096 51937
rect 639664 51925 639670 51937
rect 206090 51897 639670 51925
rect 206090 51885 206096 51897
rect 639664 51885 639670 51897
rect 639722 51885 639728 51937
rect 205936 51811 205942 51863
rect 205994 51851 206000 51863
rect 210832 51851 210838 51863
rect 205994 51823 210838 51851
rect 205994 51811 206000 51823
rect 210832 51811 210838 51823
rect 210890 51811 210896 51863
rect 204496 51663 204502 51715
rect 204554 51703 204560 51715
rect 212272 51703 212278 51715
rect 204554 51675 212278 51703
rect 204554 51663 204560 51675
rect 212272 51663 212278 51675
rect 212330 51663 212336 51715
rect 204592 51589 204598 51641
rect 204650 51629 204656 51641
rect 213040 51629 213046 51641
rect 204650 51601 213046 51629
rect 204650 51589 204656 51601
rect 213040 51589 213046 51601
rect 213098 51589 213104 51641
rect 202960 51515 202966 51567
rect 203018 51555 203024 51567
rect 215248 51555 215254 51567
rect 203018 51527 215254 51555
rect 203018 51515 203024 51527
rect 215248 51515 215254 51527
rect 215306 51515 215312 51567
rect 145552 51367 145558 51419
rect 145610 51407 145616 51419
rect 238000 51407 238006 51419
rect 145610 51379 238006 51407
rect 145610 51367 145616 51379
rect 238000 51367 238006 51379
rect 238058 51367 238064 51419
rect 145744 51293 145750 51345
rect 145802 51333 145808 51345
rect 237136 51333 237142 51345
rect 145802 51305 237142 51333
rect 145802 51293 145808 51305
rect 237136 51293 237142 51305
rect 237194 51293 237200 51345
rect 143920 51219 143926 51271
rect 143978 51259 143984 51271
rect 145552 51259 145558 51271
rect 143978 51231 145558 51259
rect 143978 51219 143984 51231
rect 145552 51219 145558 51231
rect 145610 51219 145616 51271
rect 145840 51219 145846 51271
rect 145898 51259 145904 51271
rect 236368 51259 236374 51271
rect 145898 51231 236374 51259
rect 145898 51219 145904 51231
rect 236368 51219 236374 51231
rect 236426 51219 236432 51271
rect 146416 51145 146422 51197
rect 146474 51185 146480 51197
rect 237520 51185 237526 51197
rect 146474 51157 237526 51185
rect 146474 51145 146480 51157
rect 237520 51145 237526 51157
rect 237578 51145 237584 51197
rect 144400 51071 144406 51123
rect 144458 51111 144464 51123
rect 234544 51111 234550 51123
rect 144458 51083 234550 51111
rect 144458 51071 144464 51083
rect 234544 51071 234550 51083
rect 234602 51071 234608 51123
rect 144592 50997 144598 51049
rect 144650 51037 144656 51049
rect 234160 51037 234166 51049
rect 144650 51009 234166 51037
rect 144650 50997 144656 51009
rect 234160 50997 234166 51009
rect 234218 50997 234224 51049
rect 144784 50923 144790 50975
rect 144842 50963 144848 50975
rect 234928 50963 234934 50975
rect 144842 50935 234934 50963
rect 144842 50923 144848 50935
rect 234928 50923 234934 50935
rect 234986 50923 234992 50975
rect 145936 50849 145942 50901
rect 145994 50889 146000 50901
rect 235792 50889 235798 50901
rect 145994 50861 235798 50889
rect 145994 50849 146000 50861
rect 235792 50849 235798 50861
rect 235850 50849 235856 50901
rect 146032 50775 146038 50827
rect 146090 50815 146096 50827
rect 235312 50815 235318 50827
rect 146090 50787 235318 50815
rect 146090 50775 146096 50787
rect 235312 50775 235318 50787
rect 235370 50775 235376 50827
rect 145168 50701 145174 50753
rect 145226 50741 145232 50753
rect 230896 50741 230902 50753
rect 145226 50713 230902 50741
rect 145226 50701 145232 50713
rect 230896 50701 230902 50713
rect 230954 50701 230960 50753
rect 145264 50627 145270 50679
rect 145322 50667 145328 50679
rect 232720 50667 232726 50679
rect 145322 50639 232726 50667
rect 145322 50627 145328 50639
rect 232720 50627 232726 50639
rect 232778 50627 232784 50679
rect 146512 50553 146518 50605
rect 146570 50593 146576 50605
rect 232336 50593 232342 50605
rect 146570 50565 232342 50593
rect 146570 50553 146576 50565
rect 232336 50553 232342 50565
rect 232394 50553 232400 50605
rect 146608 50479 146614 50531
rect 146666 50519 146672 50531
rect 230992 50519 230998 50531
rect 146666 50491 230998 50519
rect 146666 50479 146672 50491
rect 230992 50479 230998 50491
rect 231050 50479 231056 50531
rect 146704 50405 146710 50457
rect 146762 50445 146768 50457
rect 233104 50445 233110 50457
rect 146762 50417 233110 50445
rect 146762 50405 146768 50417
rect 233104 50405 233110 50417
rect 233162 50405 233168 50457
rect 146800 50331 146806 50383
rect 146858 50371 146864 50383
rect 231376 50371 231382 50383
rect 146858 50343 231382 50371
rect 146858 50331 146864 50343
rect 231376 50331 231382 50343
rect 231434 50331 231440 50383
rect 145552 50257 145558 50309
rect 145610 50297 145616 50309
rect 227536 50297 227542 50309
rect 145610 50269 227542 50297
rect 145610 50257 145616 50269
rect 227536 50257 227542 50269
rect 227594 50257 227600 50309
rect 144688 50183 144694 50235
rect 144746 50223 144752 50235
rect 228784 50223 228790 50235
rect 144746 50195 228790 50223
rect 144746 50183 144752 50195
rect 228784 50183 228790 50195
rect 228842 50183 228848 50235
rect 144880 50109 144886 50161
rect 144938 50149 144944 50161
rect 228688 50149 228694 50161
rect 144938 50121 228694 50149
rect 144938 50109 144944 50121
rect 228688 50109 228694 50121
rect 228746 50109 228752 50161
rect 144976 50035 144982 50087
rect 145034 50075 145040 50087
rect 229168 50075 229174 50087
rect 145034 50047 229174 50075
rect 145034 50035 145040 50047
rect 229168 50035 229174 50047
rect 229226 50035 229232 50087
rect 145072 49961 145078 50013
rect 145130 50001 145136 50013
rect 230128 50001 230134 50013
rect 145130 49973 230134 50001
rect 145130 49961 145136 49973
rect 230128 49961 230134 49973
rect 230186 49961 230192 50013
rect 144112 49887 144118 49939
rect 144170 49927 144176 49939
rect 226960 49927 226966 49939
rect 144170 49899 226966 49927
rect 144170 49887 144176 49899
rect 226960 49887 226966 49899
rect 227018 49887 227024 49939
rect 144016 49813 144022 49865
rect 144074 49853 144080 49865
rect 226096 49853 226102 49865
rect 144074 49825 226102 49853
rect 144074 49813 144080 49825
rect 226096 49813 226102 49825
rect 226154 49813 226160 49865
rect 144304 49739 144310 49791
rect 144362 49779 144368 49791
rect 225712 49779 225718 49791
rect 144362 49751 225718 49779
rect 144362 49739 144368 49751
rect 225712 49739 225718 49751
rect 225770 49739 225776 49791
rect 146128 49665 146134 49717
rect 146186 49705 146192 49717
rect 241936 49705 241942 49717
rect 146186 49677 241942 49705
rect 146186 49665 146192 49677
rect 241936 49665 241942 49677
rect 241994 49665 242000 49717
rect 145360 49591 145366 49643
rect 145418 49631 145424 49643
rect 239728 49631 239734 49643
rect 145418 49603 239734 49631
rect 145418 49591 145424 49603
rect 239728 49591 239734 49603
rect 239786 49591 239792 49643
rect 144496 49517 144502 49569
rect 144554 49557 144560 49569
rect 226480 49557 226486 49569
rect 144554 49529 226486 49557
rect 144554 49517 144560 49529
rect 226480 49517 226486 49529
rect 226538 49517 226544 49569
rect 146224 49443 146230 49495
rect 146282 49483 146288 49495
rect 241168 49483 241174 49495
rect 146282 49455 241174 49483
rect 146282 49443 146288 49455
rect 241168 49443 241174 49455
rect 241226 49443 241232 49495
rect 145456 49295 145462 49347
rect 145514 49335 145520 49347
rect 238960 49335 238966 49347
rect 145514 49307 238966 49335
rect 145514 49295 145520 49307
rect 238960 49295 238966 49307
rect 239018 49295 239024 49347
rect 146320 49221 146326 49273
rect 146378 49261 146384 49273
rect 240784 49261 240790 49273
rect 146378 49233 240790 49261
rect 146378 49221 146384 49233
rect 240784 49221 240790 49233
rect 240842 49221 240848 49273
rect 145648 49147 145654 49199
rect 145706 49187 145712 49199
rect 237616 49187 237622 49199
rect 145706 49159 237622 49187
rect 145706 49147 145712 49159
rect 237616 49147 237622 49159
rect 237674 49147 237680 49199
rect 202576 48925 202582 48977
rect 202634 48965 202640 48977
rect 214288 48965 214294 48977
rect 202634 48937 214294 48965
rect 202634 48925 202640 48937
rect 214288 48925 214294 48937
rect 214346 48925 214352 48977
rect 216304 48925 216310 48977
rect 216362 48965 216368 48977
rect 264880 48965 264886 48977
rect 216362 48937 264886 48965
rect 216362 48925 216368 48937
rect 264880 48925 264886 48937
rect 264938 48925 264944 48977
rect 627184 48925 627190 48977
rect 627242 48965 627248 48977
rect 636112 48965 636118 48977
rect 627242 48937 636118 48965
rect 627242 48925 627248 48937
rect 636112 48925 636118 48937
rect 636170 48925 636176 48977
rect 202672 48851 202678 48903
rect 202730 48891 202736 48903
rect 215056 48891 215062 48903
rect 202730 48863 215062 48891
rect 202730 48851 202736 48863
rect 215056 48851 215062 48863
rect 215114 48851 215120 48903
rect 215152 48851 215158 48903
rect 215210 48891 215216 48903
rect 226576 48891 226582 48903
rect 215210 48863 226582 48891
rect 215210 48851 215216 48863
rect 226576 48851 226582 48863
rect 226634 48851 226640 48903
rect 202768 48777 202774 48829
rect 202826 48817 202832 48829
rect 215440 48817 215446 48829
rect 202826 48789 215446 48817
rect 202826 48777 202832 48789
rect 215440 48777 215446 48789
rect 215498 48777 215504 48829
rect 204688 48629 204694 48681
rect 204746 48669 204752 48681
rect 208912 48669 208918 48681
rect 204746 48641 208918 48669
rect 204746 48629 204752 48641
rect 208912 48629 208918 48641
rect 208970 48629 208976 48681
rect 204496 48555 204502 48607
rect 204554 48595 204560 48607
rect 217648 48595 217654 48607
rect 204554 48567 217654 48595
rect 204554 48555 204560 48567
rect 217648 48555 217654 48567
rect 217706 48555 217712 48607
rect 203824 48481 203830 48533
rect 203882 48521 203888 48533
rect 216880 48521 216886 48533
rect 203882 48493 216886 48521
rect 203882 48481 203888 48493
rect 216880 48481 216886 48493
rect 216938 48481 216944 48533
rect 203728 48407 203734 48459
rect 203786 48447 203792 48459
rect 203786 48419 209246 48447
rect 203786 48407 203792 48419
rect 209218 48373 209246 48419
rect 209296 48407 209302 48459
rect 209354 48447 209360 48459
rect 235408 48447 235414 48459
rect 209354 48419 235414 48447
rect 209354 48407 209360 48419
rect 235408 48407 235414 48419
rect 235466 48407 235472 48459
rect 217264 48373 217270 48385
rect 209218 48345 217270 48373
rect 217264 48333 217270 48345
rect 217322 48333 217328 48385
rect 628912 48259 628918 48311
rect 628970 48299 628976 48311
rect 663376 48299 663382 48311
rect 628970 48271 663382 48299
rect 628970 48259 628976 48271
rect 663376 48259 663382 48271
rect 663434 48259 663440 48311
rect 147664 48185 147670 48237
rect 147722 48225 147728 48237
rect 201616 48225 201622 48237
rect 147722 48197 201622 48225
rect 147722 48185 147728 48197
rect 201616 48185 201622 48197
rect 201674 48185 201680 48237
rect 203440 48185 203446 48237
rect 203498 48225 203504 48237
rect 211600 48225 211606 48237
rect 203498 48197 211606 48225
rect 203498 48185 203504 48197
rect 211600 48185 211606 48197
rect 211658 48185 211664 48237
rect 216112 48225 216118 48237
rect 211714 48197 216118 48225
rect 147568 48111 147574 48163
rect 147626 48151 147632 48163
rect 211714 48151 211742 48197
rect 216112 48185 216118 48197
rect 216170 48185 216176 48237
rect 147626 48123 211742 48151
rect 147626 48111 147632 48123
rect 216016 48111 216022 48163
rect 216074 48151 216080 48163
rect 639376 48151 639382 48163
rect 216074 48123 639382 48151
rect 216074 48111 216080 48123
rect 639376 48111 639382 48123
rect 639434 48111 639440 48163
rect 202384 48037 202390 48089
rect 202442 48077 202448 48089
rect 216496 48077 216502 48089
rect 202442 48049 216502 48077
rect 202442 48037 202448 48049
rect 216496 48037 216502 48049
rect 216554 48037 216560 48089
rect 216592 48037 216598 48089
rect 216650 48077 216656 48089
rect 224752 48077 224758 48089
rect 216650 48049 224758 48077
rect 216650 48037 216656 48049
rect 224752 48037 224758 48049
rect 224810 48037 224816 48089
rect 148144 47963 148150 48015
rect 148202 48003 148208 48015
rect 230512 48003 230518 48015
rect 148202 47975 230518 48003
rect 148202 47963 148208 47975
rect 230512 47963 230518 47975
rect 230570 47963 230576 48015
rect 203344 47889 203350 47941
rect 203402 47929 203408 47941
rect 203402 47901 208862 47929
rect 203402 47889 203408 47901
rect 203248 47815 203254 47867
rect 203306 47855 203312 47867
rect 208720 47855 208726 47867
rect 203306 47827 208726 47855
rect 203306 47815 203312 47827
rect 208720 47815 208726 47827
rect 208778 47815 208784 47867
rect 208834 47781 208862 47901
rect 208912 47889 208918 47941
rect 208970 47929 208976 47941
rect 221680 47929 221686 47941
rect 208970 47901 221686 47929
rect 208970 47889 208976 47901
rect 221680 47889 221686 47901
rect 221738 47889 221744 47941
rect 211600 47815 211606 47867
rect 211658 47855 211664 47867
rect 219088 47855 219094 47867
rect 211658 47827 219094 47855
rect 211658 47815 211664 47827
rect 219088 47815 219094 47827
rect 219146 47815 219152 47867
rect 219472 47781 219478 47793
rect 208834 47753 219478 47781
rect 219472 47741 219478 47753
rect 219530 47741 219536 47793
rect 148528 47667 148534 47719
rect 148586 47707 148592 47719
rect 231952 47707 231958 47719
rect 148586 47679 231958 47707
rect 148586 47667 148592 47679
rect 231952 47667 231958 47679
rect 232010 47667 232016 47719
rect 627952 47667 627958 47719
rect 628010 47707 628016 47719
rect 663184 47707 663190 47719
rect 628010 47679 663190 47707
rect 628010 47667 628016 47679
rect 663184 47667 663190 47679
rect 663242 47667 663248 47719
rect 148912 47593 148918 47645
rect 148970 47633 148976 47645
rect 229744 47633 229750 47645
rect 148970 47605 229750 47633
rect 148970 47593 148976 47605
rect 229744 47593 229750 47605
rect 229802 47593 229808 47645
rect 208720 47519 208726 47571
rect 208778 47559 208784 47571
rect 219856 47559 219862 47571
rect 208778 47531 219862 47559
rect 208778 47519 208784 47531
rect 219856 47519 219862 47531
rect 219914 47519 219920 47571
rect 201616 47445 201622 47497
rect 201674 47485 201680 47497
rect 208336 47485 208342 47497
rect 201674 47457 208342 47485
rect 201674 47445 201680 47457
rect 208336 47445 208342 47457
rect 208394 47445 208400 47497
rect 148336 47371 148342 47423
rect 148394 47411 148400 47423
rect 209296 47411 209302 47423
rect 148394 47383 209302 47411
rect 148394 47371 148400 47383
rect 209296 47371 209302 47383
rect 209354 47371 209360 47423
rect 209392 47371 209398 47423
rect 209450 47411 209456 47423
rect 233584 47411 233590 47423
rect 209450 47383 233590 47411
rect 209450 47371 209456 47383
rect 233584 47371 233590 47383
rect 233642 47371 233648 47423
rect 209602 46865 215486 46893
rect 149488 46779 149494 46831
rect 149546 46819 149552 46831
rect 209392 46819 209398 46831
rect 149546 46791 209398 46819
rect 149546 46779 149552 46791
rect 209392 46779 209398 46791
rect 209450 46779 209456 46831
rect 149680 46705 149686 46757
rect 149738 46745 149744 46757
rect 209602 46745 209630 46865
rect 215458 46819 215486 46865
rect 217840 46853 217846 46905
rect 217898 46893 217904 46905
rect 639952 46893 639958 46905
rect 217898 46865 639958 46893
rect 217898 46853 217904 46865
rect 639952 46853 639958 46865
rect 640010 46853 640016 46905
rect 233296 46819 233302 46831
rect 215458 46791 233302 46819
rect 233296 46779 233302 46791
rect 233354 46779 233360 46831
rect 149738 46717 209630 46745
rect 149738 46705 149744 46717
rect 209680 46705 209686 46757
rect 209738 46745 209744 46757
rect 215152 46745 215158 46757
rect 209738 46717 215158 46745
rect 209738 46705 209744 46717
rect 215152 46705 215158 46717
rect 215210 46705 215216 46757
rect 215248 46705 215254 46757
rect 215306 46745 215312 46757
rect 223120 46745 223126 46757
rect 215306 46717 223126 46745
rect 215306 46705 215312 46717
rect 223120 46705 223126 46717
rect 223178 46705 223184 46757
rect 149296 46631 149302 46683
rect 149354 46671 149360 46683
rect 161296 46671 161302 46683
rect 149354 46643 161302 46671
rect 149354 46631 149360 46643
rect 161296 46631 161302 46643
rect 161354 46631 161360 46683
rect 181360 46631 181366 46683
rect 181418 46671 181424 46683
rect 221776 46671 221782 46683
rect 181418 46643 221782 46671
rect 181418 46631 181424 46643
rect 221776 46631 221782 46643
rect 221834 46631 221840 46683
rect 202480 46557 202486 46609
rect 202538 46597 202544 46609
rect 202538 46569 208286 46597
rect 202538 46557 202544 46569
rect 147856 46483 147862 46535
rect 147914 46523 147920 46535
rect 147914 46495 208190 46523
rect 147914 46483 147920 46495
rect 202288 46409 202294 46461
rect 202346 46449 202352 46461
rect 202346 46421 208094 46449
rect 202346 46409 202352 46421
rect 147952 46335 147958 46387
rect 148010 46375 148016 46387
rect 207856 46375 207862 46387
rect 148010 46347 207862 46375
rect 148010 46335 148016 46347
rect 207856 46335 207862 46347
rect 207914 46335 207920 46387
rect 202000 46261 202006 46313
rect 202058 46301 202064 46313
rect 207952 46301 207958 46313
rect 202058 46273 207958 46301
rect 202058 46261 202064 46273
rect 207952 46261 207958 46273
rect 208010 46261 208016 46313
rect 208066 46301 208094 46421
rect 208162 46375 208190 46495
rect 208258 46449 208286 46569
rect 208528 46557 208534 46609
rect 208586 46597 208592 46609
rect 216592 46597 216598 46609
rect 208586 46569 216598 46597
rect 208586 46557 208592 46569
rect 216592 46557 216598 46569
rect 216650 46557 216656 46609
rect 216688 46557 216694 46609
rect 216746 46597 216752 46609
rect 639856 46597 639862 46609
rect 216746 46569 639862 46597
rect 216746 46557 216752 46569
rect 639856 46557 639862 46569
rect 639914 46557 639920 46609
rect 208336 46483 208342 46535
rect 208394 46523 208400 46535
rect 220912 46523 220918 46535
rect 208394 46495 220918 46523
rect 208394 46483 208400 46495
rect 220912 46483 220918 46495
rect 220970 46483 220976 46535
rect 221776 46483 221782 46535
rect 221834 46523 221840 46535
rect 228304 46523 228310 46535
rect 221834 46495 228310 46523
rect 221834 46483 221840 46495
rect 228304 46483 228310 46495
rect 228362 46483 228368 46535
rect 222160 46449 222166 46461
rect 208258 46421 222166 46449
rect 222160 46409 222166 46421
rect 222218 46409 222224 46461
rect 224656 46375 224662 46387
rect 208162 46347 224662 46375
rect 224656 46335 224662 46347
rect 224714 46335 224720 46387
rect 225328 46301 225334 46313
rect 208066 46273 225334 46301
rect 225328 46261 225334 46273
rect 225386 46261 225392 46313
rect 147760 46187 147766 46239
rect 147818 46227 147824 46239
rect 223888 46227 223894 46239
rect 147818 46199 223894 46227
rect 147818 46187 147824 46199
rect 223888 46187 223894 46199
rect 223946 46187 223952 46239
rect 202192 46113 202198 46165
rect 202250 46153 202256 46165
rect 222064 46153 222070 46165
rect 202250 46125 222070 46153
rect 202250 46113 202256 46125
rect 222064 46113 222070 46125
rect 222122 46113 222128 46165
rect 205168 45151 205174 45203
rect 205226 45191 205232 45203
rect 403120 45191 403126 45203
rect 205226 45163 403126 45191
rect 205226 45151 205232 45163
rect 403120 45151 403126 45163
rect 403178 45151 403184 45203
rect 206992 45077 206998 45129
rect 207050 45117 207056 45129
rect 408880 45117 408886 45129
rect 207050 45089 408886 45117
rect 207050 45077 207056 45089
rect 408880 45077 408886 45089
rect 408938 45077 408944 45129
rect 207376 45003 207382 45055
rect 207434 45043 207440 45055
rect 406288 45043 406294 45055
rect 207434 45015 406294 45043
rect 207434 45003 207440 45015
rect 406288 45003 406294 45015
rect 406346 45003 406352 45055
rect 208048 44929 208054 44981
rect 208106 44969 208112 44981
rect 446512 44969 446518 44981
rect 208106 44941 446518 44969
rect 208106 44929 208112 44941
rect 446512 44929 446518 44941
rect 446570 44929 446576 44981
rect 209200 44855 209206 44907
rect 209258 44895 209264 44907
rect 499984 44895 499990 44907
rect 209258 44867 499990 44895
rect 209258 44855 209264 44867
rect 499984 44855 499990 44867
rect 500042 44855 500048 44907
rect 205264 44781 205270 44833
rect 205322 44821 205328 44833
rect 508240 44821 508246 44833
rect 205322 44793 508246 44821
rect 205322 44781 205328 44793
rect 508240 44781 508246 44793
rect 508298 44781 508304 44833
rect 209584 44707 209590 44759
rect 209642 44747 209648 44759
rect 523888 44747 523894 44759
rect 209642 44719 523894 44747
rect 209642 44707 209648 44719
rect 523888 44707 523894 44719
rect 523946 44707 523952 44759
rect 205552 44633 205558 44685
rect 205610 44673 205616 44685
rect 521200 44673 521206 44685
rect 205610 44645 521206 44673
rect 205610 44633 205616 44645
rect 521200 44633 521206 44645
rect 521258 44633 521264 44685
rect 613456 44633 613462 44685
rect 613514 44673 613520 44685
rect 635536 44673 635542 44685
rect 613514 44645 635542 44673
rect 613514 44633 613520 44645
rect 635536 44633 635542 44645
rect 635594 44633 635600 44685
rect 508240 43227 508246 43279
rect 508298 43267 508304 43279
rect 508298 43239 520382 43267
rect 508298 43227 508304 43239
rect 520354 43205 520382 43239
rect 520336 43153 520342 43205
rect 520394 43153 520400 43205
rect 206608 42339 206614 42391
rect 206666 42379 206672 42391
rect 310096 42379 310102 42391
rect 206666 42351 310102 42379
rect 206666 42339 206672 42351
rect 310096 42339 310102 42351
rect 310154 42339 310160 42391
rect 201328 42117 201334 42169
rect 201386 42157 201392 42169
rect 405232 42157 405238 42169
rect 201386 42129 405238 42157
rect 201386 42117 201392 42129
rect 405232 42117 405238 42129
rect 405290 42117 405296 42169
rect 207664 42043 207670 42095
rect 207722 42083 207728 42095
rect 460048 42083 460054 42095
rect 207722 42055 460054 42083
rect 207722 42043 207728 42055
rect 460048 42043 460054 42055
rect 460106 42043 460112 42095
rect 459184 41969 459190 42021
rect 459242 42009 459248 42021
rect 463696 42009 463702 42021
rect 459242 41981 463702 42009
rect 459242 41969 459248 41981
rect 463696 41969 463702 41981
rect 463754 41969 463760 42021
rect 403120 41895 403126 41947
rect 403178 41935 403184 41947
rect 403178 41907 405182 41935
rect 403178 41895 403184 41907
rect 405154 41861 405182 41907
rect 409090 41861 409392 41868
rect 405154 41840 409392 41861
rect 405154 41833 409118 41840
rect 514864 41747 514870 41799
rect 514922 41747 514928 41799
rect 208432 41673 208438 41725
rect 208490 41713 208496 41725
rect 514882 41713 514910 41747
rect 208490 41685 514910 41713
rect 208490 41673 208496 41685
rect 499984 40341 499990 40393
rect 500042 40381 500048 40393
rect 500042 40353 501182 40381
rect 500042 40341 500048 40353
rect 501154 40307 501182 40353
rect 512560 40307 512566 40319
rect 501154 40279 512566 40307
rect 512560 40267 512566 40279
rect 512618 40267 512624 40319
rect 446512 37381 446518 37433
rect 446570 37421 446576 37433
rect 459184 37421 459190 37433
rect 446570 37393 459190 37421
rect 446570 37381 446576 37393
rect 459184 37381 459190 37393
rect 459242 37381 459248 37433
<< via1 >>
rect 447766 1005671 447818 1005723
rect 95062 1005523 95114 1005575
rect 437206 1005523 437258 1005575
rect 93622 1005449 93674 1005501
rect 100726 1005449 100778 1005501
rect 108694 1005449 108746 1005501
rect 433270 1005449 433322 1005501
rect 469174 1005597 469226 1005649
rect 440566 1005449 440618 1005501
rect 441622 1005449 441674 1005501
rect 93718 1005375 93770 1005427
rect 115222 1005375 115274 1005427
rect 358678 1005375 358730 1005427
rect 379126 1005375 379178 1005427
rect 431638 1005375 431690 1005427
rect 466486 1005523 466538 1005575
rect 443446 1005449 443498 1005501
rect 470998 1005449 471050 1005501
rect 504598 1005449 504650 1005501
rect 441814 1005375 441866 1005427
rect 471862 1005375 471914 1005427
rect 498742 1005375 498794 1005427
rect 512662 1005375 512714 1005427
rect 92566 1005301 92618 1005353
rect 109462 1005301 109514 1005353
rect 298294 1005301 298346 1005353
rect 308758 1005301 308810 1005353
rect 365014 1005301 365066 1005353
rect 383638 1005301 383690 1005353
rect 425302 1005301 425354 1005353
rect 434710 1005301 434762 1005353
rect 434806 1005301 434858 1005353
rect 437782 1005301 437834 1005353
rect 440566 1005301 440618 1005353
rect 92374 1005227 92426 1005279
rect 106582 1005227 106634 1005279
rect 217270 1005227 217322 1005279
rect 218902 1005227 218954 1005279
rect 299542 1005227 299594 1005279
rect 309622 1005227 309674 1005279
rect 424534 1005227 424586 1005279
rect 440854 1005227 440906 1005279
rect 198742 1005153 198794 1005205
rect 207286 1005153 207338 1005205
rect 305302 1005153 305354 1005205
rect 314230 1005153 314282 1005205
rect 325462 1005153 325514 1005205
rect 331222 1005153 331274 1005205
rect 358006 1005153 358058 1005205
rect 383542 1005153 383594 1005205
rect 426070 1005153 426122 1005205
rect 452950 1005301 453002 1005353
rect 441046 1005227 441098 1005279
rect 472054 1005227 472106 1005279
rect 502294 1005227 502346 1005279
rect 516790 1005227 516842 1005279
rect 521398 1005227 521450 1005279
rect 554518 1005227 554570 1005279
rect 572854 1005375 572906 1005427
rect 435574 1005079 435626 1005131
rect 440758 1005079 440810 1005131
rect 443446 1005153 443498 1005205
rect 447766 1005153 447818 1005205
rect 469366 1005153 469418 1005205
rect 508630 1005153 508682 1005205
rect 523990 1005153 524042 1005205
rect 553750 1005153 553802 1005205
rect 571894 1005227 571946 1005279
rect 562486 1005153 562538 1005205
rect 572950 1005153 573002 1005205
rect 434710 1005005 434762 1005057
rect 437206 1005005 437258 1005057
rect 100726 1004931 100778 1004983
rect 114166 1004931 114218 1004983
rect 512662 1004857 512714 1004909
rect 521206 1004857 521258 1004909
rect 356758 1003895 356810 1003947
rect 377206 1003895 377258 1003947
rect 359062 1003821 359114 1003873
rect 379990 1003821 380042 1003873
rect 428086 1003821 428138 1003873
rect 466486 1003821 466538 1003873
rect 501142 1003821 501194 1003873
rect 519478 1003821 519530 1003873
rect 551734 1003821 551786 1003873
rect 570646 1003821 570698 1003873
rect 355990 1003747 356042 1003799
rect 377110 1003747 377162 1003799
rect 423382 1003747 423434 1003799
rect 469270 1003747 469322 1003799
rect 556534 1003747 556586 1003799
rect 574486 1003747 574538 1003799
rect 195286 1003673 195338 1003725
rect 211702 1003673 211754 1003725
rect 359926 1003673 359978 1003725
rect 380086 1003673 380138 1003725
rect 426454 1003673 426506 1003725
rect 470134 1003673 470186 1003725
rect 500374 1003673 500426 1003725
rect 521014 1003673 521066 1003725
rect 552598 1003673 552650 1003725
rect 573046 1003673 573098 1003725
rect 144214 1002563 144266 1002615
rect 151510 1002563 151562 1002615
rect 143734 1002489 143786 1002541
rect 152854 1002489 152906 1002541
rect 502774 1002489 502826 1002541
rect 515446 1002489 515498 1002541
rect 559126 1002489 559178 1002541
rect 566134 1002489 566186 1002541
rect 143926 1002415 143978 1002467
rect 153622 1002415 153674 1002467
rect 489526 1002415 489578 1002467
rect 144022 1002341 144074 1002393
rect 150358 1002341 150410 1002393
rect 503446 1002415 503498 1002467
rect 513526 1002415 513578 1002467
rect 559894 1002415 559946 1002467
rect 564502 1002415 564554 1002467
rect 518614 1002341 518666 1002393
rect 560566 1002341 560618 1002393
rect 564694 1002341 564746 1002393
rect 564790 1002341 564842 1002393
rect 568726 1002341 568778 1002393
rect 144310 1002267 144362 1002319
rect 178486 1002267 178538 1002319
rect 505078 1002267 505130 1002319
rect 521494 1002267 521546 1002319
rect 561526 1002267 561578 1002319
rect 565366 1002267 565418 1002319
rect 573046 1002193 573098 1002245
rect 573334 1002193 573386 1002245
rect 452950 1002045 453002 1002097
rect 461590 1002045 461642 1002097
rect 469366 1002045 469418 1002097
rect 472150 1002045 472202 1002097
rect 566134 1001601 566186 1001653
rect 570166 1001601 570218 1001653
rect 513526 1001453 513578 1001505
rect 515734 1001453 515786 1001505
rect 572854 1001453 572906 1001505
rect 574102 1001453 574154 1001505
rect 434038 1001083 434090 1001135
rect 472630 1001083 472682 1001135
rect 432502 1001009 432554 1001061
rect 472534 1001009 472586 1001061
rect 564502 1001009 564554 1001061
rect 567766 1001009 567818 1001061
rect 571894 1001009 571946 1001061
rect 573238 1001009 573290 1001061
rect 430870 1000935 430922 1000987
rect 472342 1000935 472394 1000987
rect 510934 1000935 510986 1000987
rect 516694 1000935 516746 1000987
rect 195094 1000861 195146 1000913
rect 208150 1000861 208202 1000913
rect 428950 1000861 429002 1000913
rect 472630 1000861 472682 1000913
rect 143830 1000787 143882 1000839
rect 160246 1000787 160298 1000839
rect 361558 1000787 361610 1000839
rect 383638 1000787 383690 1000839
rect 427318 1000787 427370 1000839
rect 472438 1000787 472490 1000839
rect 509302 1000787 509354 1000839
rect 516694 1000787 516746 1000839
rect 469174 1000713 469226 1000765
rect 469558 1000713 469610 1000765
rect 298198 1000343 298250 1000395
rect 305302 1000343 305354 1000395
rect 613462 999825 613514 999877
rect 625558 999825 625610 999877
rect 610582 999751 610634 999803
rect 625462 999751 625514 999803
rect 601846 999677 601898 999729
rect 625846 999677 625898 999729
rect 379126 999603 379178 999655
rect 381430 999603 381482 999655
rect 596182 999603 596234 999655
rect 625750 999603 625802 999655
rect 246646 999529 246698 999581
rect 260758 999529 260810 999581
rect 590710 999529 590762 999581
rect 625366 999529 625418 999581
rect 144118 999455 144170 999507
rect 155158 999455 155210 999507
rect 247702 999455 247754 999507
rect 258838 999455 258890 999507
rect 497590 999455 497642 999507
rect 516694 999455 516746 999507
rect 565366 999455 565418 999507
rect 61846 999381 61898 999433
rect 74710 999381 74762 999433
rect 92950 999381 93002 999433
rect 123862 999381 123914 999433
rect 143734 999381 143786 999433
rect 156886 999381 156938 999433
rect 195190 999381 195242 999433
rect 226006 999381 226058 999433
rect 246550 999381 246602 999433
rect 259606 999381 259658 999433
rect 298102 999381 298154 999433
rect 311254 999381 311306 999433
rect 377110 999381 377162 999433
rect 379030 999381 379082 999433
rect 466582 999381 466634 999433
rect 472246 999381 472298 999433
rect 540310 999381 540362 999433
rect 570262 999381 570314 999433
rect 506326 999307 506378 999359
rect 516694 999307 516746 999359
rect 590614 999455 590666 999507
rect 625846 999455 625898 999507
rect 590518 999381 590570 999433
rect 625654 999381 625706 999433
rect 571030 999307 571082 999359
rect 461590 998715 461642 998767
rect 466582 998715 466634 998767
rect 567766 998567 567818 998619
rect 570838 998567 570890 998619
rect 195382 997901 195434 997953
rect 209398 997901 209450 997953
rect 328342 997901 328394 997953
rect 367894 997901 367946 997953
rect 371446 997901 371498 997953
rect 555190 997901 555242 997953
rect 559894 997901 559946 997953
rect 570262 997901 570314 997953
rect 610678 997901 610730 997953
rect 325462 997827 325514 997879
rect 350134 997827 350186 997879
rect 557302 997827 557354 997879
rect 596182 997827 596234 997879
rect 318454 997753 318506 997805
rect 369046 997753 369098 997805
rect 556150 997753 556202 997805
rect 590518 997753 590570 997805
rect 564694 997679 564746 997731
rect 590614 997679 590666 997731
rect 573334 997605 573386 997657
rect 590710 997605 590762 997657
rect 573238 997531 573290 997583
rect 610582 997531 610634 997583
rect 559894 997457 559946 997509
rect 570550 997457 570602 997509
rect 572950 997457 573002 997509
rect 601846 997457 601898 997509
rect 574486 997383 574538 997435
rect 613462 997383 613514 997435
rect 377206 997087 377258 997139
rect 382006 997087 382058 997139
rect 510262 996569 510314 996621
rect 521110 996569 521162 996621
rect 259126 996495 259178 996547
rect 263926 996495 263978 996547
rect 379990 996495 380042 996547
rect 380278 996495 380330 996547
rect 507862 996495 507914 996547
rect 521206 996495 521258 996547
rect 316342 996421 316394 996473
rect 162646 996125 162698 996177
rect 213334 996125 213386 996177
rect 265078 996125 265130 996177
rect 276502 996125 276554 996177
rect 302326 996125 302378 996177
rect 316342 996125 316394 996177
rect 423286 996347 423338 996399
rect 440758 996347 440810 996399
rect 511894 996199 511946 996251
rect 399862 996125 399914 996177
rect 408886 996125 408938 996177
rect 408982 996125 409034 996177
rect 423286 996125 423338 996177
rect 436438 996125 436490 996177
rect 513430 996125 513482 996177
rect 563734 996125 563786 996177
rect 164086 996051 164138 996103
rect 215638 996051 215690 996103
rect 218902 996051 218954 996103
rect 266902 996051 266954 996103
rect 266998 996051 267050 996103
rect 318646 996051 318698 996103
rect 367126 996051 367178 996103
rect 437782 996051 437834 996103
rect 471862 996051 471914 996103
rect 511126 996051 511178 996103
rect 562774 996051 562826 996103
rect 103894 995977 103946 996029
rect 115222 995977 115274 996029
rect 164182 995977 164234 996029
rect 276502 995977 276554 996029
rect 92374 995903 92426 995955
rect 92470 995903 92522 995955
rect 101494 995903 101546 995955
rect 106486 995903 106538 995955
rect 113398 995903 113450 995955
rect 144118 995903 144170 995955
rect 144406 995903 144458 995955
rect 151990 995903 152042 995955
rect 195670 995903 195722 995955
rect 200278 995903 200330 995955
rect 200950 995903 201002 995955
rect 213046 995903 213098 995955
rect 216790 995903 216842 995955
rect 246454 995903 246506 995955
rect 254902 995829 254954 995881
rect 257302 995829 257354 995881
rect 81046 995755 81098 995807
rect 84790 995755 84842 995807
rect 91510 995755 91562 995807
rect 105430 995755 105482 995807
rect 113398 995755 113450 995807
rect 118102 995755 118154 995807
rect 132406 995755 132458 995807
rect 142966 995755 143018 995807
rect 143734 995755 143786 995807
rect 164086 995755 164138 995807
rect 165622 995755 165674 995807
rect 188086 995755 188138 995807
rect 202870 995755 202922 995807
rect 236470 995755 236522 995807
rect 245686 995755 245738 995807
rect 246550 995755 246602 995807
rect 250486 995755 250538 995807
rect 254038 995755 254090 995807
rect 268534 995755 268586 995807
rect 273718 995755 273770 995807
rect 74902 995681 74954 995733
rect 82486 995681 82538 995733
rect 85366 995681 85418 995733
rect 99766 995681 99818 995733
rect 141046 995681 141098 995733
rect 143830 995681 143882 995733
rect 163990 995681 164042 995733
rect 166198 995681 166250 995733
rect 188854 995681 188906 995733
rect 204214 995681 204266 995733
rect 250390 995681 250442 995733
rect 255670 995681 255722 995733
rect 133078 995607 133130 995659
rect 146806 995607 146858 995659
rect 194422 995607 194474 995659
rect 195094 995607 195146 995659
rect 139318 995533 139370 995585
rect 143926 995533 143978 995585
rect 191926 995533 191978 995585
rect 195190 995533 195242 995585
rect 82294 995459 82346 995511
rect 99670 995459 99722 995511
rect 184342 995459 184394 995511
rect 201526 995459 201578 995511
rect 370198 995903 370250 995955
rect 374518 995903 374570 995955
rect 287446 995607 287498 995659
rect 298294 995829 298346 995881
rect 299446 995829 299498 995881
rect 304726 995829 304778 995881
rect 368854 995829 368906 995881
rect 436438 995977 436490 996029
rect 470998 995977 471050 996029
rect 511894 995977 511946 996029
rect 513430 995977 513482 996029
rect 564790 995977 564842 996029
rect 625366 995977 625418 996029
rect 291190 995755 291242 995807
rect 305686 995755 305738 995807
rect 297334 995681 297386 995733
rect 298102 995681 298154 995733
rect 302422 995681 302474 995733
rect 310294 995755 310346 995807
rect 360982 995755 361034 995807
rect 365782 995755 365834 995807
rect 371446 995755 371498 995807
rect 399862 995903 399914 995955
rect 472342 995903 472394 995955
rect 383542 995829 383594 995881
rect 472438 995829 472490 995881
rect 523510 995903 523562 995955
rect 523894 995829 523946 995881
rect 625462 995903 625514 995955
rect 610678 995829 610730 995881
rect 616342 995829 616394 995881
rect 625654 995829 625706 995881
rect 383638 995755 383690 995807
rect 384982 995755 385034 995807
rect 389398 995755 389450 995807
rect 472630 995755 472682 995807
rect 474070 995755 474122 995807
rect 477718 995755 477770 995807
rect 480982 995755 481034 995807
rect 523990 995755 524042 995807
rect 527830 995755 527882 995807
rect 528982 995755 529034 995807
rect 529846 995755 529898 995807
rect 537142 995755 537194 995807
rect 540310 995755 540362 995807
rect 563734 995755 563786 995807
rect 567478 995755 567530 995807
rect 625846 995755 625898 995807
rect 626518 995755 626570 995807
rect 630934 995755 630986 995807
rect 631510 995755 631562 995807
rect 634582 995755 634634 995807
rect 365878 995681 365930 995733
rect 377302 995681 377354 995733
rect 383734 995681 383786 995733
rect 384406 995681 384458 995733
rect 472534 995681 472586 995733
rect 473302 995681 473354 995733
rect 524086 995681 524138 995733
rect 528406 995681 528458 995733
rect 625750 995681 625802 995733
rect 627094 995681 627146 995733
rect 291766 995607 291818 995659
rect 307318 995607 307370 995659
rect 472726 995607 472778 995659
rect 474646 995607 474698 995659
rect 523798 995607 523850 995659
rect 525334 995607 525386 995659
rect 562774 995607 562826 995659
rect 567382 995607 567434 995659
rect 625942 995607 625994 995659
rect 627862 995607 627914 995659
rect 287926 995533 287978 995585
rect 302326 995533 302378 995585
rect 472246 995533 472298 995585
rect 476374 995533 476426 995585
rect 302230 995459 302282 995511
rect 466582 995459 466634 995511
rect 482038 995533 482090 995585
rect 523702 995533 523754 995585
rect 524758 995533 524810 995585
rect 625558 995533 625610 995585
rect 630166 995533 630218 995585
rect 81622 995385 81674 995437
rect 103126 995385 103178 995437
rect 129334 995385 129386 995437
rect 146806 995385 146858 995437
rect 183766 995385 183818 995437
rect 206614 995385 206666 995437
rect 472150 995385 472202 995437
rect 478294 995459 478346 995511
rect 523606 995459 523658 995511
rect 526102 995459 526154 995511
rect 85702 995311 85754 995363
rect 92470 995311 92522 995363
rect 133990 995311 134042 995363
rect 144310 995311 144362 995363
rect 133414 995237 133466 995289
rect 144406 995237 144458 995289
rect 469462 995237 469514 995289
rect 482710 995385 482762 995437
rect 521110 995385 521162 995437
rect 537142 995385 537194 995437
rect 518614 995311 518666 995363
rect 530566 995311 530618 995363
rect 521302 995163 521354 995215
rect 633718 995163 633770 995215
rect 485590 995089 485642 995141
rect 643990 995089 644042 995141
rect 226006 995015 226058 995067
rect 642454 995015 642506 995067
rect 320758 994719 320810 994771
rect 325462 994719 325514 994771
rect 227542 994423 227594 994475
rect 236758 994423 236810 994475
rect 238966 994423 239018 994475
rect 630838 994349 630890 994401
rect 632374 994349 632426 994401
rect 247798 994127 247850 994179
rect 250486 994127 250538 994179
rect 82582 994053 82634 994105
rect 133942 994053 133994 994105
rect 243094 993979 243146 994031
rect 247702 993979 247754 994031
rect 235798 993905 235850 993957
rect 246454 993905 246506 993957
rect 180502 993831 180554 993883
rect 198742 993831 198794 993883
rect 234934 993831 234986 993883
rect 247702 993831 247754 993883
rect 77686 993757 77738 993809
rect 100726 993757 100778 993809
rect 131830 993757 131882 993809
rect 158614 993757 158666 993809
rect 182998 993757 183050 993809
rect 210166 993757 210218 993809
rect 232150 993757 232202 993809
rect 243094 993757 243146 993809
rect 259126 994053 259178 994105
rect 574102 993979 574154 994031
rect 635254 993979 635306 994031
rect 570646 993831 570698 993883
rect 636118 993831 636170 993883
rect 77302 993683 77354 993735
rect 108214 993683 108266 993735
rect 128470 993683 128522 993735
rect 159478 993683 159530 993735
rect 181366 993683 181418 993735
rect 212662 993683 212714 993735
rect 232534 993683 232586 993735
rect 470134 993757 470186 993809
rect 484150 993757 484202 993809
rect 515734 993757 515786 993809
rect 535318 993757 535370 993809
rect 570550 993757 570602 993809
rect 637366 993757 637418 993809
rect 243286 993683 243338 993735
rect 247606 993683 247658 993735
rect 283510 993683 283562 993735
rect 302422 993683 302474 993735
rect 506614 993683 506666 993735
rect 538966 993683 539018 993735
rect 557974 993683 558026 993735
rect 641014 993683 641066 993735
rect 179830 993609 179882 993661
rect 211030 993609 211082 993661
rect 238966 993609 239018 993661
rect 279286 993609 279338 993661
rect 282838 993609 282890 993661
rect 313846 993609 313898 993661
rect 362326 993609 362378 993661
rect 398806 993609 398858 993661
rect 429718 993609 429770 993661
rect 487798 993609 487850 993661
rect 530614 993609 530666 993661
rect 630838 993609 630890 993661
rect 638902 993609 638954 993661
rect 643606 993609 643658 993661
rect 115318 993461 115370 993513
rect 126742 993461 126794 993513
rect 115222 993387 115274 993439
rect 162646 993387 162698 993439
rect 126742 993313 126794 993365
rect 162934 993461 162986 993513
rect 214390 993535 214442 993587
rect 265750 993535 265802 993587
rect 317494 993535 317546 993587
rect 328342 993535 328394 993587
rect 469462 993535 469514 993587
rect 479158 993535 479210 993587
rect 489526 993535 489578 993587
rect 331222 992129 331274 992181
rect 332566 992129 332618 992181
rect 547126 992129 547178 992181
rect 650902 992129 650954 992181
rect 633718 990649 633770 990701
rect 640438 990649 640490 990701
rect 643990 990649 644042 990701
rect 649846 990649 649898 990701
rect 640726 989761 640778 989813
rect 649558 989761 649610 989813
rect 638518 989317 638570 989369
rect 649942 989317 649994 989369
rect 616342 989243 616394 989295
rect 643222 989243 643274 989295
rect 223126 987763 223178 987815
rect 235606 987763 235658 987815
rect 518422 987763 518474 987815
rect 527542 987763 527594 987815
rect 642454 987763 642506 987815
rect 647350 987763 647402 987815
rect 219382 987097 219434 987149
rect 221878 987097 221930 987149
rect 154486 986727 154538 986779
rect 163990 986727 164042 986779
rect 374422 986505 374474 986557
rect 397750 986505 397802 986557
rect 570262 986505 570314 986557
rect 592438 986505 592490 986557
rect 273622 986431 273674 986483
rect 284278 986431 284330 986483
rect 316918 986431 316970 986483
rect 320758 986431 320810 986483
rect 326806 986431 326858 986483
rect 349078 986431 349130 986483
rect 377494 986431 377546 986483
rect 414070 986431 414122 986483
rect 445078 986431 445130 986483
rect 478966 986431 479018 986483
rect 521398 986431 521450 986483
rect 543766 986431 543818 986483
rect 573142 986431 573194 986483
rect 608758 986431 608810 986483
rect 73366 986357 73418 986409
rect 93622 986357 93674 986409
rect 138262 986357 138314 986409
rect 164086 986357 164138 986409
rect 273718 986357 273770 986409
rect 300406 986357 300458 986409
rect 323926 986357 323978 986409
rect 365398 986357 365450 986409
rect 374518 986357 374570 986409
rect 430294 986357 430346 986409
rect 440662 986357 440714 986409
rect 495094 986357 495146 986409
rect 518518 986357 518570 986409
rect 560086 986357 560138 986409
rect 570454 986357 570506 986409
rect 624886 986357 624938 986409
rect 203158 986283 203210 986335
rect 213046 986283 213098 986335
rect 640438 986283 640490 986335
rect 646102 986283 646154 986335
rect 89590 985839 89642 985891
rect 93718 985839 93770 985891
rect 90646 985765 90698 985817
rect 45142 985469 45194 985521
rect 63286 985469 63338 985521
rect 50518 985395 50570 985447
rect 122038 985395 122090 985447
rect 181462 985469 181514 985521
rect 47734 985321 47786 985373
rect 186934 985321 186986 985373
rect 187318 985321 187370 985373
rect 63286 985247 63338 985299
rect 90646 985247 90698 985299
rect 251734 985247 251786 985299
rect 45046 985173 45098 985225
rect 316726 985173 316778 985225
rect 44950 985099 45002 985151
rect 381622 985099 381674 985151
rect 444886 985099 444938 985151
rect 462742 985099 462794 985151
rect 44854 985025 44906 985077
rect 446422 985025 446474 985077
rect 42550 984951 42602 985003
rect 511414 984951 511466 985003
rect 633622 984951 633674 985003
rect 641110 984951 641162 985003
rect 643222 984877 643274 984929
rect 650134 984877 650186 984929
rect 65206 983841 65258 983893
rect 94966 983841 95018 983893
rect 44758 983767 44810 983819
rect 115318 983767 115370 983819
rect 44566 983693 44618 983745
rect 115222 983693 115274 983745
rect 44662 983619 44714 983671
rect 118102 983619 118154 983671
rect 567382 983619 567434 983671
rect 652246 983619 652298 983671
rect 65110 983545 65162 983597
rect 145270 983545 145322 983597
rect 567478 983545 567530 983597
rect 652342 983545 652394 983597
rect 65014 983471 65066 983523
rect 195670 983471 195722 983523
rect 568726 983471 568778 983523
rect 652438 983471 652490 983523
rect 64918 980807 64970 980859
rect 243286 980807 243338 980859
rect 643606 980807 643658 980859
rect 649750 980807 649802 980859
rect 64822 980733 64874 980785
rect 298486 980733 298538 980785
rect 647350 980733 647402 980785
rect 649462 980733 649514 980785
rect 64630 980659 64682 980711
rect 316918 980659 316970 980711
rect 630838 980659 630890 980711
rect 673942 980659 673994 980711
rect 64726 980585 64778 980637
rect 410326 980585 410378 980637
rect 630742 980585 630794 980637
rect 674518 980585 674570 980637
rect 646102 980511 646154 980563
rect 649366 980511 649418 980563
rect 53302 970595 53354 970647
rect 59542 970595 59594 970647
rect 42166 967265 42218 967317
rect 42550 967265 42602 967317
rect 42166 960975 42218 961027
rect 42358 960975 42410 961027
rect 673942 958977 673994 959029
rect 675478 958977 675530 959029
rect 675094 958385 675146 958437
rect 675382 958385 675434 958437
rect 675190 956979 675242 957031
rect 675478 956979 675530 957031
rect 42358 956165 42410 956217
rect 59350 956165 59402 956217
rect 42070 955203 42122 955255
rect 42934 955203 42986 955255
rect 669526 954685 669578 954737
rect 675382 954685 675434 954737
rect 42166 954611 42218 954663
rect 43030 954611 43082 954663
rect 674038 953871 674090 953923
rect 675478 953871 675530 953923
rect 649462 953279 649514 953331
rect 653686 953279 653738 953331
rect 674134 952021 674186 952073
rect 675478 952021 675530 952073
rect 655222 944843 655274 944895
rect 674710 944843 674762 944895
rect 655126 944621 655178 944673
rect 674710 944621 674762 944673
rect 652342 943141 652394 943193
rect 672886 943141 672938 943193
rect 672310 942549 672362 942601
rect 674422 942549 674474 942601
rect 654358 942031 654410 942083
rect 674710 942031 674762 942083
rect 652438 941883 652490 941935
rect 674614 941883 674666 941935
rect 672886 941809 672938 941861
rect 673846 941809 673898 941861
rect 53206 941735 53258 941787
rect 59542 941735 59594 941787
rect 652246 939071 652298 939123
rect 674902 939071 674954 939123
rect 654454 927453 654506 927505
rect 666742 927453 666794 927505
rect 50326 927379 50378 927431
rect 59542 927379 59594 927431
rect 649462 927379 649514 927431
rect 679798 927379 679850 927431
rect 47446 912949 47498 913001
rect 59542 912949 59594 913001
rect 654454 912949 654506 913001
rect 660982 912949 661034 913001
rect 42646 908065 42698 908117
rect 53206 908065 53258 908117
rect 42262 907473 42314 907525
rect 50326 907473 50378 907525
rect 42646 904809 42698 904861
rect 44662 904809 44714 904861
rect 654454 901479 654506 901531
rect 663958 901479 664010 901531
rect 53206 898593 53258 898645
rect 59542 898593 59594 898645
rect 42358 889639 42410 889691
rect 44566 889639 44618 889691
rect 50422 884163 50474 884215
rect 59542 884163 59594 884215
rect 654454 878391 654506 878443
rect 660886 878391 660938 878443
rect 40054 872619 40106 872671
rect 40438 872619 40490 872671
rect 674230 872101 674282 872153
rect 675478 872101 675530 872153
rect 674902 871879 674954 871931
rect 675574 871879 675626 871931
rect 39958 869807 40010 869859
rect 40438 869807 40490 869859
rect 674998 868993 675050 869045
rect 675478 868993 675530 869045
rect 674326 868327 674378 868379
rect 675382 868327 675434 868379
rect 673654 867809 673706 867861
rect 675382 867809 675434 867861
rect 654454 867291 654506 867343
rect 663766 867291 663818 867343
rect 674902 866847 674954 866899
rect 675094 866847 675146 866899
rect 666646 865293 666698 865345
rect 675382 865293 675434 865345
rect 675382 862925 675434 862977
rect 675382 862555 675434 862607
rect 50326 855377 50378 855429
rect 59542 855377 59594 855429
rect 654454 855377 654506 855429
rect 661174 855377 661226 855429
rect 39958 852491 40010 852543
rect 40054 852343 40106 852395
rect 674806 846719 674858 846771
rect 675094 846719 675146 846771
rect 675382 846719 675434 846771
rect 675574 846719 675626 846771
rect 40054 846645 40106 846697
rect 40150 846645 40202 846697
rect 53398 840947 53450 840999
rect 59542 840947 59594 840999
rect 654454 832363 654506 832415
rect 669718 832363 669770 832415
rect 50614 829477 50666 829529
rect 58198 829477 58250 829529
rect 39958 826591 40010 826643
rect 40150 826591 40202 826643
rect 674422 826517 674474 826569
rect 674710 826517 674762 826569
rect 675478 826517 675530 826569
rect 675670 826517 675722 826569
rect 42358 823853 42410 823905
rect 50422 823853 50474 823905
rect 42358 822225 42410 822277
rect 53206 822225 53258 822277
rect 42454 821855 42506 821907
rect 58966 821855 59018 821907
rect 654454 820819 654506 820871
rect 667030 820819 667082 820871
rect 40150 817859 40202 817911
rect 43318 817859 43370 817911
rect 47542 812161 47594 812213
rect 59542 812161 59594 812213
rect 654454 809275 654506 809327
rect 664054 809275 664106 809327
rect 674422 806389 674474 806441
rect 674614 806389 674666 806441
rect 675286 806389 675338 806441
rect 675670 806389 675722 806441
rect 42262 805131 42314 805183
rect 44758 805131 44810 805183
rect 42454 803577 42506 803629
rect 42934 803577 42986 803629
rect 40246 803429 40298 803481
rect 42454 803429 42506 803481
rect 41974 802393 42026 802445
rect 43030 802393 43082 802445
rect 43510 800839 43562 800891
rect 44854 800839 44906 800891
rect 42262 800247 42314 800299
rect 43414 800247 43466 800299
rect 41878 800173 41930 800225
rect 41878 799729 41930 799781
rect 42166 798027 42218 798079
rect 42454 798027 42506 798079
rect 53206 797805 53258 797857
rect 59542 797805 59594 797857
rect 42070 797287 42122 797339
rect 43510 797287 43562 797339
rect 42166 796251 42218 796303
rect 43126 796251 43178 796303
rect 43126 796103 43178 796155
rect 43414 796103 43466 796155
rect 42166 794993 42218 795045
rect 42742 794993 42794 795045
rect 42166 793809 42218 793861
rect 42454 793809 42506 793861
rect 42166 793143 42218 793195
rect 43030 793143 43082 793195
rect 43126 792107 43178 792159
rect 43606 792107 43658 792159
rect 43030 791959 43082 792011
rect 43606 791959 43658 792011
rect 42262 790035 42314 790087
rect 42838 790035 42890 790087
rect 42166 789887 42218 789939
rect 43126 789887 43178 789939
rect 42262 788851 42314 788903
rect 42934 788851 42986 788903
rect 42166 787001 42218 787053
rect 43030 787001 43082 787053
rect 42166 786409 42218 786461
rect 42454 786409 42506 786461
rect 654454 786261 654506 786313
rect 666838 786261 666890 786313
rect 42070 785595 42122 785647
rect 42742 785595 42794 785647
rect 674518 784929 674570 784981
rect 675382 784929 675434 784981
rect 672214 783449 672266 783501
rect 675382 783449 675434 783501
rect 674998 783005 675050 783057
rect 675382 783005 675434 783057
rect 672502 782265 672554 782317
rect 674614 782265 674666 782317
rect 675382 782265 675434 782317
rect 663862 780489 663914 780541
rect 675094 780489 675146 780541
rect 42742 780415 42794 780467
rect 50614 780415 50666 780467
rect 674422 780415 674474 780467
rect 675478 780415 675530 780467
rect 42454 779897 42506 779949
rect 47542 779897 47594 779949
rect 672694 779749 672746 779801
rect 675382 779749 675434 779801
rect 672022 779305 672074 779357
rect 675478 779305 675530 779357
rect 42742 778861 42794 778913
rect 53398 778861 53450 778913
rect 672118 778565 672170 778617
rect 675382 778565 675434 778617
rect 672406 777603 672458 777655
rect 675478 777603 675530 777655
rect 675094 777011 675146 777063
rect 675382 777011 675434 777063
rect 674806 775457 674858 775509
rect 675382 775457 675434 775509
rect 654454 774717 654506 774769
rect 669814 774717 669866 774769
rect 674230 773607 674282 773659
rect 675382 773607 675434 773659
rect 53398 771831 53450 771883
rect 59542 771831 59594 771883
rect 660982 767761 661034 767813
rect 674710 767761 674762 767813
rect 666742 766873 666794 766925
rect 674710 766873 674762 766925
rect 663958 765837 664010 765889
rect 674326 765837 674378 765889
rect 672310 765245 672362 765297
rect 674710 765245 674762 765297
rect 672598 763987 672650 764039
rect 674710 763987 674762 764039
rect 654454 763247 654506 763299
rect 661078 763247 661130 763299
rect 670966 763173 671018 763225
rect 672886 763173 672938 763225
rect 674710 763173 674762 763225
rect 672886 762507 672938 762559
rect 674710 762507 674762 762559
rect 42934 758067 42986 758119
rect 43222 758067 43274 758119
rect 42934 757919 42986 757971
rect 44950 757919 45002 757971
rect 50422 757475 50474 757527
rect 58198 757475 58250 757527
rect 42454 757253 42506 757305
rect 43510 757253 43562 757305
rect 41974 757105 42026 757157
rect 43702 757105 43754 757157
rect 41878 757031 41930 757083
rect 43606 757031 43658 757083
rect 41782 756957 41834 757009
rect 42070 756957 42122 757009
rect 43318 756957 43370 757009
rect 41782 756735 41834 756787
rect 42166 754071 42218 754123
rect 42934 754071 42986 754123
rect 42934 753923 42986 753975
rect 43222 753923 43274 753975
rect 42070 753035 42122 753087
rect 43126 753035 43178 753087
rect 42934 751851 42986 751903
rect 42070 751777 42122 751829
rect 42742 751777 42794 751829
rect 42838 751777 42890 751829
rect 42934 751703 42986 751755
rect 43702 751703 43754 751755
rect 42070 751111 42122 751163
rect 42838 751111 42890 751163
rect 42838 750963 42890 751015
rect 43606 750963 43658 751015
rect 42166 750371 42218 750423
rect 43126 750371 43178 750423
rect 43126 750223 43178 750275
rect 43510 750223 43562 750275
rect 674038 750223 674090 750275
rect 674422 750223 674474 750275
rect 42070 749927 42122 749979
rect 42934 749927 42986 749979
rect 42262 748891 42314 748943
rect 42838 748891 42890 748943
rect 649558 748817 649610 748869
rect 679798 748817 679850 748869
rect 42166 747411 42218 747463
rect 42454 747411 42506 747463
rect 42070 746079 42122 746131
rect 43126 746079 43178 746131
rect 42166 745635 42218 745687
rect 43030 745635 43082 745687
rect 42166 743785 42218 743837
rect 42742 743785 42794 743837
rect 42070 743045 42122 743097
rect 42838 743045 42890 743097
rect 47542 743045 47594 743097
rect 58582 743045 58634 743097
rect 42166 742379 42218 742431
rect 42934 742379 42986 742431
rect 674902 737865 674954 737917
rect 675382 737865 675434 737917
rect 672502 737643 672554 737695
rect 675478 737643 675530 737695
rect 660982 737347 661034 737399
rect 675094 737347 675146 737399
rect 654454 737273 654506 737325
rect 663958 737273 664010 737325
rect 42646 737199 42698 737251
rect 53398 737199 53450 737251
rect 42358 736681 42410 736733
rect 50422 736681 50474 736733
rect 674134 735645 674186 735697
rect 675478 735645 675530 735697
rect 42358 735423 42410 735475
rect 58966 735423 59018 735475
rect 675190 734905 675242 734957
rect 675382 734905 675434 734957
rect 672310 733573 672362 733625
rect 675478 733573 675530 733625
rect 675190 732315 675242 732367
rect 675478 732315 675530 732367
rect 675094 732019 675146 732071
rect 675382 732019 675434 732071
rect 674710 730465 674762 730517
rect 675478 730465 675530 730517
rect 50422 728615 50474 728667
rect 59542 728615 59594 728667
rect 674614 728615 674666 728667
rect 675478 728615 675530 728667
rect 674806 726321 674858 726373
rect 675094 726321 675146 726373
rect 663766 722473 663818 722525
rect 674326 722473 674378 722525
rect 660886 721881 660938 721933
rect 674806 721881 674858 721933
rect 661174 720845 661226 720897
rect 674326 720845 674378 720897
rect 672598 720253 672650 720305
rect 674806 720253 674858 720305
rect 674038 720031 674090 720083
rect 674326 720031 674378 720083
rect 671926 718995 671978 719047
rect 674806 718995 674858 719047
rect 42262 718699 42314 718751
rect 44950 718699 45002 718751
rect 672886 717811 672938 717863
rect 674518 717811 674570 717863
rect 672598 717145 672650 717197
rect 672886 717145 672938 717197
rect 43126 717071 43178 717123
rect 45046 717071 45098 717123
rect 670966 717071 671018 717123
rect 679702 717071 679754 717123
rect 40246 714999 40298 715051
rect 41878 714999 41930 715051
rect 53398 714259 53450 714311
rect 59542 714259 59594 714311
rect 654454 714259 654506 714311
rect 664150 714259 664202 714311
rect 41590 714111 41642 714163
rect 43510 714111 43562 714163
rect 41494 714037 41546 714089
rect 41686 714037 41738 714089
rect 43606 714037 43658 714089
rect 41974 713815 42026 713867
rect 43318 713815 43370 713867
rect 41782 713519 41834 713571
rect 43318 711521 43370 711573
rect 42934 711447 42986 711499
rect 43126 711447 43178 711499
rect 43414 711373 43466 711425
rect 42934 711299 42986 711351
rect 43702 711225 43754 711277
rect 42166 710855 42218 710907
rect 43414 710855 43466 710907
rect 672214 710485 672266 710537
rect 674422 710485 674474 710537
rect 42166 709893 42218 709945
rect 42358 709893 42410 709945
rect 672406 709893 672458 709945
rect 674806 709893 674858 709945
rect 672022 709005 672074 709057
rect 674422 709005 674474 709057
rect 42166 707895 42218 707947
rect 43702 707895 43754 707947
rect 672694 707377 672746 707429
rect 674422 707377 674474 707429
rect 42934 707229 42986 707281
rect 43606 707229 43658 707281
rect 672118 706785 672170 706837
rect 674806 706785 674858 706837
rect 42550 706415 42602 706467
rect 43510 706415 43562 706467
rect 42262 705601 42314 705653
rect 43126 705601 43178 705653
rect 42070 703677 42122 703729
rect 42838 703677 42890 703729
rect 42166 702863 42218 702915
rect 42934 702863 42986 702915
rect 649654 702715 649706 702767
rect 679798 702715 679850 702767
rect 672502 702641 672554 702693
rect 674806 702641 674858 702693
rect 42166 702271 42218 702323
rect 42550 702271 42602 702323
rect 42070 700569 42122 700621
rect 43030 700569 43082 700621
rect 42166 700051 42218 700103
rect 42838 700051 42890 700103
rect 670966 699903 671018 699955
rect 679702 699903 679754 699955
rect 42358 699829 42410 699881
rect 59542 699829 59594 699881
rect 42646 693983 42698 694035
rect 53398 693983 53450 694035
rect 672214 692873 672266 692925
rect 675382 692873 675434 692925
rect 42646 692429 42698 692481
rect 50422 692429 50474 692481
rect 672406 692429 672458 692481
rect 674806 692429 674858 692481
rect 675478 692429 675530 692481
rect 654838 691245 654890 691297
rect 666934 691245 666986 691297
rect 674326 690653 674378 690705
rect 675478 690653 675530 690705
rect 675094 689765 675146 689817
rect 675382 689765 675434 689817
rect 672118 688581 672170 688633
rect 675478 688581 675530 688633
rect 674230 687323 674282 687375
rect 675478 687323 675530 687375
rect 669622 686213 669674 686265
rect 675382 686213 675434 686265
rect 50422 685473 50474 685525
rect 58678 685473 58730 685525
rect 674518 685473 674570 685525
rect 675478 685473 675530 685525
rect 674902 683623 674954 683675
rect 675478 683623 675530 683675
rect 667030 677481 667082 677533
rect 674806 677481 674858 677533
rect 649750 676815 649802 676867
rect 653686 676815 653738 676867
rect 669718 676445 669770 676497
rect 674422 676445 674474 676497
rect 664054 675853 664106 675905
rect 674806 675853 674858 675905
rect 42358 675631 42410 675683
rect 45046 675631 45098 675683
rect 671926 674817 671978 674869
rect 674422 674817 674474 674869
rect 41590 674521 41642 674573
rect 43126 674521 43178 674573
rect 672694 674003 672746 674055
rect 674422 674003 674474 674055
rect 670966 673115 671018 673167
rect 672502 673115 672554 673167
rect 674806 673115 674858 673167
rect 40246 672153 40298 672205
rect 41014 672153 41066 672205
rect 41686 672005 41738 672057
rect 42646 672005 42698 672057
rect 42262 671931 42314 671983
rect 42454 671931 42506 671983
rect 43318 671339 43370 671391
rect 45142 671339 45194 671391
rect 53398 671043 53450 671095
rect 58390 671043 58442 671095
rect 672598 670969 672650 671021
rect 675094 670969 675146 671021
rect 43126 670821 43178 670873
rect 43510 670821 43562 670873
rect 41878 670747 41930 670799
rect 43222 670747 43274 670799
rect 41782 670599 41834 670651
rect 41974 670599 42026 670651
rect 42934 670599 42986 670651
rect 41782 670303 41834 670355
rect 674422 669563 674474 669615
rect 674902 669563 674954 669615
rect 42454 669193 42506 669245
rect 42838 668897 42890 668949
rect 654454 668157 654506 668209
rect 661270 668157 661322 668209
rect 42166 667861 42218 667913
rect 43318 667861 43370 667913
rect 42166 666677 42218 666729
rect 42934 666677 42986 666729
rect 42166 664827 42218 664879
rect 42838 664827 42890 664879
rect 42838 664679 42890 664731
rect 43606 664679 43658 664731
rect 42166 664161 42218 664213
rect 43126 664161 43178 664213
rect 43126 664013 43178 664065
rect 43510 664013 43562 664065
rect 42550 663495 42602 663547
rect 42166 663347 42218 663399
rect 42262 662385 42314 662437
rect 43030 662385 43082 662437
rect 672310 661645 672362 661697
rect 674710 661645 674762 661697
rect 42166 661053 42218 661105
rect 42838 661053 42890 661105
rect 42166 659647 42218 659699
rect 42934 659647 42986 659699
rect 42070 659055 42122 659107
rect 42550 659055 42602 659107
rect 42166 656835 42218 656887
rect 42838 656835 42890 656887
rect 42070 656761 42122 656813
rect 43126 656761 43178 656813
rect 42838 656687 42890 656739
rect 59542 656687 59594 656739
rect 649750 656687 649802 656739
rect 679798 656687 679850 656739
rect 672406 650915 672458 650967
rect 674806 650915 674858 650967
rect 674614 650841 674666 650893
rect 674998 650841 675050 650893
rect 42454 649731 42506 649783
rect 51862 649731 51914 649783
rect 42454 649509 42506 649561
rect 53398 649509 53450 649561
rect 671926 648251 671978 648303
rect 675286 648251 675338 648303
rect 672886 648029 672938 648081
rect 675190 648029 675242 648081
rect 674806 647585 674858 647637
rect 675094 647585 675146 647637
rect 674614 646401 674666 646453
rect 675382 646401 675434 646453
rect 666742 645217 666794 645269
rect 675190 645217 675242 645269
rect 654454 645143 654506 645195
rect 669718 645143 669770 645195
rect 674806 645069 674858 645121
rect 675094 645069 675146 645121
rect 671638 644551 671690 644603
rect 675478 644551 675530 644603
rect 51862 644477 51914 644529
rect 59542 644477 59594 644529
rect 672310 644033 672362 644085
rect 675478 644033 675530 644085
rect 672598 643367 672650 643419
rect 675382 643367 675434 643419
rect 671446 642257 671498 642309
rect 675478 642257 675530 642309
rect 675190 641813 675242 641865
rect 675382 641813 675434 641865
rect 670870 633599 670922 633651
rect 674998 633599 675050 633651
rect 669814 632489 669866 632541
rect 674710 632489 674762 632541
rect 42262 632415 42314 632467
rect 45142 632415 45194 632467
rect 666838 631749 666890 631801
rect 674710 631749 674762 631801
rect 670966 630713 671018 630765
rect 672502 630713 672554 630765
rect 661078 630565 661130 630617
rect 674134 630565 674186 630617
rect 672694 630491 672746 630543
rect 673846 630491 673898 630543
rect 42934 628419 42986 628471
rect 43606 628419 43658 628471
rect 42454 627901 42506 627953
rect 47734 627901 47786 627953
rect 40054 627827 40106 627879
rect 41206 627827 41258 627879
rect 43126 627827 43178 627879
rect 43414 627827 43466 627879
rect 47638 627827 47690 627879
rect 58390 627827 58442 627879
rect 671734 627827 671786 627879
rect 673846 627827 673898 627879
rect 41686 627753 41738 627805
rect 43510 627753 43562 627805
rect 41494 627679 41546 627731
rect 43126 627679 43178 627731
rect 41782 627383 41834 627435
rect 42070 627383 42122 627435
rect 43030 627383 43082 627435
rect 41782 627161 41834 627213
rect 42934 625163 42986 625215
rect 43414 625163 43466 625215
rect 42166 624645 42218 624697
rect 42454 624645 42506 624697
rect 42166 623461 42218 623513
rect 42934 623461 42986 623513
rect 42454 623313 42506 623365
rect 42934 623313 42986 623365
rect 654454 622055 654506 622107
rect 669910 622055 669962 622107
rect 42166 621611 42218 621663
rect 43030 621611 43082 621663
rect 43030 621463 43082 621515
rect 43510 621463 43562 621515
rect 42166 620353 42218 620405
rect 43126 620353 43178 620405
rect 43126 620205 43178 620257
rect 43606 620205 43658 620257
rect 672214 619169 672266 619221
rect 673846 619169 673898 619221
rect 42070 617837 42122 617889
rect 42454 617837 42506 617889
rect 672118 617837 672170 617889
rect 673846 617837 673898 617889
rect 42166 617171 42218 617223
rect 43126 617171 43178 617223
rect 42166 616653 42218 616705
rect 42934 616653 42986 616705
rect 42166 615839 42218 615891
rect 43030 615839 43082 615891
rect 42166 613989 42218 614041
rect 42838 613989 42890 614041
rect 42166 613619 42218 613671
rect 42454 613619 42506 613671
rect 42454 613471 42506 613523
rect 58390 613471 58442 613523
rect 649846 613471 649898 613523
rect 679702 613471 679754 613523
rect 654454 613397 654506 613449
rect 669526 613397 669578 613449
rect 42070 612805 42122 612857
rect 42742 612805 42794 612857
rect 42742 607699 42794 607751
rect 51862 607699 51914 607751
rect 42742 606811 42794 606863
rect 53398 606811 53450 606863
rect 672214 603629 672266 603681
rect 674614 603629 674666 603681
rect 675286 603629 675338 603681
rect 673750 602815 673802 602867
rect 674806 602815 674858 602867
rect 675478 602815 675530 602867
rect 672022 602667 672074 602719
rect 675382 602667 675434 602719
rect 663766 602075 663818 602127
rect 671830 602001 671882 602053
rect 675190 602001 675242 602053
rect 672118 601927 672170 601979
rect 675094 601927 675146 601979
rect 51862 601853 51914 601905
rect 59542 601853 59594 601905
rect 675190 601853 675242 601905
rect 671350 599781 671402 599833
rect 675382 599781 675434 599833
rect 671542 599263 671594 599315
rect 675382 599263 675434 599315
rect 654454 599041 654506 599093
rect 666838 599041 666890 599093
rect 672694 598375 672746 598427
rect 675478 598375 675530 598427
rect 672502 597117 672554 597169
rect 675478 597117 675530 597169
rect 675190 596821 675242 596873
rect 675382 596821 675434 596873
rect 670870 590309 670922 590361
rect 679702 590309 679754 590361
rect 42550 589199 42602 589251
rect 45238 589199 45290 589251
rect 53398 587423 53450 587475
rect 59542 587423 59594 587475
rect 42550 586535 42602 586587
rect 43030 586535 43082 586587
rect 663958 586313 664010 586365
rect 674422 586313 674474 586365
rect 42454 586091 42506 586143
rect 43030 586091 43082 586143
rect 40054 585943 40106 585995
rect 42454 585943 42506 585995
rect 664150 585425 664202 585477
rect 674422 585425 674474 585477
rect 42838 585055 42890 585107
rect 43126 585055 43178 585107
rect 654454 585055 654506 585107
rect 661174 585055 661226 585107
rect 671734 584833 671786 584885
rect 674614 584833 674666 584885
rect 42550 584759 42602 584811
rect 43126 584759 43178 584811
rect 655126 584759 655178 584811
rect 674710 584759 674762 584811
rect 42838 584685 42890 584737
rect 50518 584685 50570 584737
rect 41782 584167 41834 584219
rect 42166 584167 42218 584219
rect 42934 584167 42986 584219
rect 41782 583945 41834 583997
rect 672406 583575 672458 583627
rect 674710 583575 674762 583627
rect 670966 583353 671018 583405
rect 674710 583353 674762 583405
rect 679990 583353 680042 583405
rect 42166 582095 42218 582147
rect 42454 582095 42506 582147
rect 42070 581429 42122 581481
rect 42838 581429 42890 581481
rect 42070 580245 42122 580297
rect 43222 580245 43274 580297
rect 43318 580023 43370 580075
rect 43606 580023 43658 580075
rect 42166 578987 42218 579039
rect 43126 578987 43178 579039
rect 672406 578839 672458 578891
rect 672790 578839 672842 578891
rect 42070 578395 42122 578447
rect 42934 578395 42986 578447
rect 42166 577655 42218 577707
rect 43030 577655 43082 577707
rect 42262 576027 42314 576079
rect 42934 576027 42986 576079
rect 671926 575361 671978 575413
rect 674710 575361 674762 575413
rect 671446 574473 671498 574525
rect 674710 574473 674762 574525
rect 672310 573585 672362 573637
rect 674422 573585 674474 573637
rect 42070 573437 42122 573489
rect 42838 573437 42890 573489
rect 654454 573141 654506 573193
rect 663958 573141 664010 573193
rect 672886 572993 672938 573045
rect 674710 572993 674762 573045
rect 42166 572623 42218 572675
rect 42454 572623 42506 572675
rect 42262 572475 42314 572527
rect 42454 572475 42506 572527
rect 671638 571957 671690 572009
rect 674422 571957 674474 572009
rect 672598 571365 672650 571417
rect 674710 571365 674762 571417
rect 42166 570995 42218 571047
rect 43030 570995 43082 571047
rect 42358 570255 42410 570307
rect 59542 570255 59594 570307
rect 42070 570181 42122 570233
rect 42454 570181 42506 570233
rect 42070 569663 42122 569715
rect 42838 569663 42890 569715
rect 649942 567369 649994 567421
rect 679798 567369 679850 567421
rect 34486 564483 34538 564535
rect 53398 564483 53450 564535
rect 654454 564409 654506 564461
rect 666646 564409 666698 564461
rect 672214 564409 672266 564461
rect 674998 564409 675050 564461
rect 42454 563447 42506 563499
rect 50518 563447 50570 563499
rect 673750 561597 673802 561649
rect 675094 561597 675146 561649
rect 674230 559525 674282 559577
rect 675382 559525 675434 559577
rect 672214 558711 672266 558763
rect 672790 558711 672842 558763
rect 53398 558637 53450 558689
rect 59542 558637 59594 558689
rect 674134 558045 674186 558097
rect 675382 558045 675434 558097
rect 660886 555825 660938 555877
rect 675190 555825 675242 555877
rect 674326 555011 674378 555063
rect 675478 555011 675530 555063
rect 674038 554493 674090 554545
rect 675382 554493 675434 554545
rect 674998 553901 675050 553953
rect 675478 553901 675530 553953
rect 674902 553161 674954 553213
rect 675382 553161 675434 553213
rect 674518 551903 674570 551955
rect 675478 551903 675530 551955
rect 675190 551533 675242 551585
rect 675382 551533 675434 551585
rect 654454 550127 654506 550179
rect 661078 550127 661130 550179
rect 674614 550053 674666 550105
rect 675478 550053 675530 550105
rect 674806 548203 674858 548255
rect 675382 548203 675434 548255
rect 42646 546205 42698 546257
rect 45334 546205 45386 546257
rect 42358 545539 42410 545591
rect 42646 545539 42698 545591
rect 41974 544577 42026 544629
rect 42934 544577 42986 544629
rect 50518 543689 50570 543741
rect 59542 543689 59594 543741
rect 40150 542875 40202 542927
rect 41974 542875 42026 542927
rect 43702 541469 43754 541521
rect 53302 541469 53354 541521
rect 655318 541469 655370 541521
rect 674710 541469 674762 541521
rect 666934 541321 666986 541373
rect 674422 541321 674474 541373
rect 41686 541247 41738 541299
rect 43414 541247 43466 541299
rect 674326 541025 674378 541077
rect 674998 541025 675050 541077
rect 41782 540951 41834 541003
rect 42166 540951 42218 541003
rect 43318 540951 43370 541003
rect 41782 540729 41834 540781
rect 661270 540729 661322 540781
rect 674710 540729 674762 540781
rect 672214 539841 672266 539893
rect 674710 539841 674762 539893
rect 42934 538731 42986 538783
rect 43510 538731 43562 538783
rect 42166 538139 42218 538191
rect 43702 538139 43754 538191
rect 42070 537029 42122 537081
rect 42838 537029 42890 537081
rect 42070 535771 42122 535823
rect 43126 535771 43178 535823
rect 43222 535771 43274 535823
rect 676630 535697 676682 535749
rect 679798 535697 679850 535749
rect 43222 535549 43274 535601
rect 42166 535253 42218 535305
rect 42742 535253 42794 535305
rect 42166 534439 42218 534491
rect 43030 534439 43082 534491
rect 43030 534291 43082 534343
rect 43414 534291 43466 534343
rect 42070 533699 42122 533751
rect 42934 533699 42986 533751
rect 42934 533551 42986 533603
rect 43510 533551 43562 533603
rect 42262 532811 42314 532863
rect 42646 532811 42698 532863
rect 672118 532737 672170 532789
rect 673846 532737 673898 532789
rect 42166 531331 42218 531383
rect 43126 531331 43178 531383
rect 671830 530813 671882 530865
rect 673846 530813 673898 530865
rect 42262 530295 42314 530347
rect 42838 530295 42890 530347
rect 672502 529851 672554 529903
rect 673846 529851 673898 529903
rect 671542 529777 671594 529829
rect 673750 529777 673802 529829
rect 42262 529629 42314 529681
rect 43030 529629 43082 529681
rect 672022 529185 672074 529237
rect 673846 529185 673898 529237
rect 42166 527631 42218 527683
rect 42934 527631 42986 527683
rect 42070 527187 42122 527239
rect 42646 527187 42698 527239
rect 42358 527039 42410 527091
rect 59446 527039 59498 527091
rect 654454 527039 654506 527091
rect 669814 527039 669866 527091
rect 672694 526891 672746 526943
rect 673846 526891 673898 526943
rect 671350 526817 671402 526869
rect 673750 526817 673802 526869
rect 42166 526447 42218 526499
rect 42742 526447 42794 526499
rect 650038 521267 650090 521319
rect 679798 521267 679850 521319
rect 654454 517937 654506 517989
rect 663862 517937 663914 517989
rect 50614 512683 50666 512735
rect 59542 512683 59594 512735
rect 654454 504025 654506 504077
rect 666646 504025 666698 504077
rect 53398 498253 53450 498305
rect 58102 498253 58154 498305
rect 674038 498031 674090 498083
rect 674998 498031 675050 498083
rect 674230 497883 674282 497935
rect 674710 497883 674762 497935
rect 674902 497883 674954 497935
rect 674230 497661 674282 497713
rect 674326 497587 674378 497639
rect 674518 497587 674570 497639
rect 669718 497291 669770 497343
rect 674422 497291 674474 497343
rect 669910 496477 669962 496529
rect 674422 496477 674474 496529
rect 655222 495515 655274 495567
rect 674710 495515 674762 495567
rect 674806 494257 674858 494309
rect 679702 494257 679754 494309
rect 654454 492481 654506 492533
rect 663862 492481 663914 492533
rect 53302 483823 53354 483875
rect 59542 483823 59594 483875
rect 654454 480937 654506 480989
rect 666934 480937 666986 480989
rect 650134 478125 650186 478177
rect 679798 478125 679850 478177
rect 654454 469985 654506 470037
rect 660982 469985 661034 470037
rect 50518 469467 50570 469519
rect 59542 469467 59594 469519
rect 654358 457923 654410 457975
rect 660982 457923 661034 457975
rect 45430 455037 45482 455089
rect 59542 455037 59594 455089
rect 654454 446379 654506 446431
rect 669718 446379 669770 446431
rect 45526 440681 45578 440733
rect 59542 440681 59594 440733
rect 42646 436907 42698 436959
rect 50614 436907 50666 436959
rect 42646 436093 42698 436145
rect 53398 436093 53450 436145
rect 654358 432023 654410 432075
rect 664054 432023 664106 432075
rect 53398 426251 53450 426303
rect 59350 426251 59402 426303
rect 654454 423291 654506 423343
rect 669622 423291 669674 423343
rect 41878 419961 41930 420013
rect 42358 419961 42410 420013
rect 42646 418555 42698 418607
rect 44662 418555 44714 418607
rect 42166 413523 42218 413575
rect 43222 413523 43274 413575
rect 41782 413375 41834 413427
rect 41782 413153 41834 413205
rect 53494 411821 53546 411873
rect 57814 411821 57866 411873
rect 42166 411303 42218 411355
rect 42358 411303 42410 411355
rect 42358 411155 42410 411207
rect 43126 411155 43178 411207
rect 42070 410489 42122 410541
rect 47446 410489 47498 410541
rect 661174 409897 661226 409949
rect 674422 409897 674474 409949
rect 42166 409453 42218 409505
rect 42742 409453 42794 409505
rect 666838 409305 666890 409357
rect 674710 409305 674762 409357
rect 655030 408935 655082 408987
rect 669526 408935 669578 408987
rect 663958 408417 664010 408469
rect 674710 408417 674762 408469
rect 42166 408195 42218 408247
rect 42838 408195 42890 408247
rect 42070 407455 42122 407507
rect 43126 407455 43178 407507
rect 42166 406863 42218 406915
rect 43030 406863 43082 406915
rect 42166 403829 42218 403881
rect 42934 403829 42986 403881
rect 42070 402941 42122 402993
rect 42358 402941 42410 402993
rect 654454 397465 654506 397517
rect 663958 397465 664010 397517
rect 42358 393913 42410 393965
rect 50518 393913 50570 393965
rect 42358 393173 42410 393225
rect 45430 393173 45482 393225
rect 42358 392285 42410 392337
rect 53302 392285 53354 392337
rect 650230 391693 650282 391745
rect 679798 391693 679850 391745
rect 653878 385921 653930 385973
rect 669622 385921 669674 385973
rect 674326 384293 674378 384345
rect 675094 384293 675146 384345
rect 674134 383109 674186 383161
rect 675382 383109 675434 383161
rect 45718 383035 45770 383087
rect 59542 383035 59594 383087
rect 674614 382443 674666 382495
rect 675478 382443 675530 382495
rect 674710 378151 674762 378203
rect 675382 378151 675434 378203
rect 674422 377559 674474 377611
rect 675382 377559 675434 377611
rect 654166 377189 654218 377241
rect 666742 377189 666794 377241
rect 674518 376819 674570 376871
rect 675478 376819 675530 376871
rect 674038 375709 674090 375761
rect 675478 375709 675530 375761
rect 42166 375191 42218 375243
rect 45430 375191 45482 375243
rect 37366 372527 37418 372579
rect 42934 372527 42986 372579
rect 42070 370159 42122 370211
rect 42262 370159 42314 370211
rect 43318 370159 43370 370211
rect 42166 369937 42218 369989
rect 42358 369937 42410 369989
rect 42358 369789 42410 369841
rect 50518 368679 50570 368731
rect 59542 368679 59594 368731
rect 42070 368087 42122 368139
rect 42358 368087 42410 368139
rect 42070 367347 42122 367399
rect 50326 367347 50378 367399
rect 42070 366237 42122 366289
rect 43030 366237 43082 366289
rect 43030 366089 43082 366141
rect 43318 366089 43370 366141
rect 42166 364979 42218 365031
rect 42742 364979 42794 365031
rect 42070 364239 42122 364291
rect 42934 364239 42986 364291
rect 42358 364091 42410 364143
rect 42838 364091 42890 364143
rect 661078 363869 661130 363921
rect 674422 363869 674474 363921
rect 42166 363647 42218 363699
rect 43126 363647 43178 363699
rect 654454 363351 654506 363403
rect 661174 363351 661226 363403
rect 669814 363277 669866 363329
rect 674614 363277 674666 363329
rect 655126 363055 655178 363107
rect 674710 363055 674762 363107
rect 42262 362093 42314 362145
rect 43030 362093 43082 362145
rect 42358 350697 42410 350749
rect 53398 350697 53450 350749
rect 42646 349661 42698 349713
rect 53494 349661 53546 349713
rect 42358 349069 42410 349121
rect 45526 349069 45578 349121
rect 650326 345591 650378 345643
rect 679798 345591 679850 345643
rect 674518 340929 674570 340981
rect 675478 340929 675530 340981
rect 53302 339819 53354 339871
rect 59542 339819 59594 339871
rect 654166 339819 654218 339871
rect 666742 339819 666794 339871
rect 674038 339523 674090 339575
rect 675382 339523 675434 339575
rect 674326 336563 674378 336615
rect 675382 336563 675434 336615
rect 674902 336267 674954 336319
rect 675094 336267 675146 336319
rect 674710 332715 674762 332767
rect 675382 332715 675434 332767
rect 674230 332197 674282 332249
rect 675478 332197 675530 332249
rect 42358 331975 42410 332027
rect 45622 331975 45674 332027
rect 674998 331753 675050 331805
rect 675382 331753 675434 331805
rect 653974 329755 654026 329807
rect 663766 329755 663818 329807
rect 37270 329311 37322 329363
rect 41782 329311 41834 329363
rect 37366 329163 37418 329215
rect 41686 329163 41738 329215
rect 37174 328349 37226 328401
rect 43126 328275 43178 328327
rect 43318 328275 43370 328327
rect 43030 328053 43082 328105
rect 41686 327239 41738 327291
rect 42358 327239 42410 327291
rect 41782 327017 41834 327069
rect 41782 326721 41834 326773
rect 53398 325463 53450 325515
rect 59542 325463 59594 325515
rect 42070 324871 42122 324923
rect 42742 324871 42794 324923
rect 42166 324131 42218 324183
rect 53206 324131 53258 324183
rect 42166 323095 42218 323147
rect 43030 323095 43082 323147
rect 43030 322947 43082 322999
rect 43318 322947 43370 322999
rect 42070 321763 42122 321815
rect 43126 321763 43178 321815
rect 42166 321245 42218 321297
rect 42358 321245 42410 321297
rect 42166 320579 42218 320631
rect 43030 320579 43082 320631
rect 663862 319913 663914 319965
rect 674710 319913 674762 319965
rect 666646 318877 666698 318929
rect 674422 318877 674474 318929
rect 666934 318285 666986 318337
rect 674710 318285 674762 318337
rect 42070 316879 42122 316931
rect 43414 316879 43466 316931
rect 45526 311033 45578 311085
rect 59542 311033 59594 311085
rect 42262 307481 42314 307533
rect 45718 307481 45770 307533
rect 42262 306741 42314 306793
rect 50518 306741 50570 306793
rect 42838 305483 42890 305535
rect 59062 305483 59114 305535
rect 650422 299563 650474 299615
rect 679798 299563 679850 299615
rect 674902 299489 674954 299541
rect 676822 299489 676874 299541
rect 675190 299415 675242 299467
rect 676918 299415 676970 299467
rect 675286 299341 675338 299393
rect 677014 299341 677066 299393
rect 45718 296677 45770 296729
rect 59542 296677 59594 296729
rect 674326 295937 674378 295989
rect 675382 295937 675434 295989
rect 674614 295345 674666 295397
rect 675478 295345 675530 295397
rect 674422 292681 674474 292733
rect 675190 292681 675242 292733
rect 42646 289055 42698 289107
rect 43222 289055 43274 289107
rect 45910 289055 45962 289107
rect 674902 288537 674954 288589
rect 675478 288537 675530 288589
rect 39958 287945 40010 287997
rect 42646 287945 42698 287997
rect 674038 287723 674090 287775
rect 675382 287723 675434 287775
rect 673942 287205 673994 287257
rect 675478 287205 675530 287257
rect 37366 286835 37418 286887
rect 42742 286835 42794 286887
rect 674230 286761 674282 286813
rect 675382 286761 675434 286813
rect 41782 283801 41834 283853
rect 42166 283801 42218 283853
rect 43318 283801 43370 283853
rect 41782 283357 41834 283409
rect 653782 282395 653834 282447
rect 660886 282395 660938 282447
rect 45814 282247 45866 282299
rect 57622 282247 57674 282299
rect 42166 281729 42218 281781
rect 42646 281729 42698 281781
rect 42166 281063 42218 281115
rect 47542 281063 47594 281115
rect 42166 279879 42218 279931
rect 42742 279879 42794 279931
rect 42166 278547 42218 278599
rect 42550 278547 42602 278599
rect 42166 277807 42218 277859
rect 43126 277807 43178 277859
rect 43222 277807 43274 277859
rect 43222 277585 43274 277637
rect 42070 277363 42122 277415
rect 42838 277363 42890 277415
rect 64630 275143 64682 275195
rect 67222 275143 67274 275195
rect 64726 275069 64778 275121
rect 66838 275069 66890 275121
rect 512758 274995 512810 275047
rect 649366 274995 649418 275047
rect 669718 274921 669770 274973
rect 674710 274921 674762 274973
rect 522262 274551 522314 274603
rect 522550 274551 522602 274603
rect 42262 274477 42314 274529
rect 42742 274477 42794 274529
rect 660982 274033 661034 274085
rect 674710 274033 674762 274085
rect 42262 273737 42314 273789
rect 43126 273737 43178 273789
rect 282166 273737 282218 273789
rect 299446 273737 299498 273789
rect 319702 273737 319754 273789
rect 339766 273737 339818 273789
rect 403126 273515 403178 273567
rect 410422 273515 410474 273567
rect 64822 273441 64874 273493
rect 72598 273441 72650 273493
rect 437782 273441 437834 273493
rect 443542 273441 443594 273493
rect 100918 273367 100970 273419
rect 120790 273367 120842 273419
rect 207286 273367 207338 273419
rect 208438 273367 208490 273419
rect 645142 273367 645194 273419
rect 665206 273367 665258 273419
rect 256342 273293 256394 273345
rect 276406 273293 276458 273345
rect 664054 273293 664106 273345
rect 674710 273293 674762 273345
rect 66166 273219 66218 273271
rect 80566 273219 80618 273271
rect 308470 272257 308522 272309
rect 392662 272257 392714 272309
rect 297814 272183 297866 272235
rect 391126 272183 391178 272235
rect 283510 272109 283562 272161
rect 411958 272109 412010 272161
rect 64918 270925 64970 270977
rect 67606 270925 67658 270977
rect 378454 270703 378506 270755
rect 379510 270703 379562 270755
rect 67222 270629 67274 270681
rect 72118 270629 72170 270681
rect 112246 270629 112298 270681
rect 132982 270629 133034 270681
rect 137110 270629 137162 270681
rect 140470 270629 140522 270681
rect 158614 270629 158666 270681
rect 161206 270629 161258 270681
rect 162166 270629 162218 270681
rect 164086 270629 164138 270681
rect 165814 270629 165866 270681
rect 166966 270629 167018 270681
rect 172822 270629 172874 270681
rect 175606 270629 175658 270681
rect 176470 270629 176522 270681
rect 178486 270629 178538 270681
rect 180022 270629 180074 270681
rect 181366 270629 181418 270681
rect 183478 270629 183530 270681
rect 184246 270629 184298 270681
rect 184342 270629 184394 270681
rect 426934 270629 426986 270681
rect 427894 270629 427946 270681
rect 540406 270629 540458 270681
rect 72598 270555 72650 270607
rect 80662 270555 80714 270607
rect 108598 270555 108650 270607
rect 130006 270555 130058 270607
rect 130102 270555 130154 270607
rect 139894 270555 139946 270607
rect 105046 270481 105098 270533
rect 139318 270481 139370 270533
rect 174070 270481 174122 270533
rect 433078 270555 433130 270607
rect 521974 270555 522026 270607
rect 551062 270555 551114 270607
rect 179158 270481 179210 270533
rect 440566 270481 440618 270533
rect 508342 270481 508394 270533
rect 566518 270481 566570 270533
rect 101494 270407 101546 270459
rect 139702 270407 139754 270459
rect 164566 270407 164618 270459
rect 427990 270407 428042 270459
rect 429334 270407 429386 270459
rect 97942 270333 97994 270385
rect 132886 270333 132938 270385
rect 132982 270333 133034 270385
rect 139126 270333 139178 270385
rect 159766 270333 159818 270385
rect 424438 270333 424490 270385
rect 432310 270333 432362 270385
rect 432694 270407 432746 270459
rect 564214 270407 564266 270459
rect 94390 270259 94442 270311
rect 140182 270259 140234 270311
rect 163414 270259 163466 270311
rect 432406 270259 432458 270311
rect 567670 270333 567722 270385
rect 577270 270259 577322 270311
rect 89590 270185 89642 270237
rect 139798 270185 139850 270237
rect 157366 270185 157418 270237
rect 429238 270185 429290 270237
rect 432118 270185 432170 270237
rect 580822 270185 580874 270237
rect 84790 270111 84842 270163
rect 140374 270111 140426 270163
rect 152566 270111 152618 270163
rect 424246 270111 424298 270163
rect 424822 270111 424874 270163
rect 578422 270111 578474 270163
rect 80086 270037 80138 270089
rect 139414 270037 139466 270089
rect 150262 270037 150314 270089
rect 427318 270037 427370 270089
rect 427798 270037 427850 270089
rect 582070 270037 582122 270089
rect 75286 269963 75338 270015
rect 68182 269815 68234 269867
rect 133270 269815 133322 269867
rect 133558 269963 133610 270015
rect 140278 269963 140330 270015
rect 146710 269963 146762 270015
rect 426262 269963 426314 270015
rect 427126 269963 427178 270015
rect 585526 269963 585578 270015
rect 139510 269889 139562 269941
rect 425782 269889 425834 269941
rect 427222 269889 427274 269941
rect 589174 269889 589226 269941
rect 140086 269815 140138 269867
rect 141910 269815 141962 269867
rect 429910 269815 429962 269867
rect 431158 269815 431210 269867
rect 432694 269815 432746 269867
rect 434902 269815 434954 269867
rect 598678 269815 598730 269867
rect 132502 269741 132554 269793
rect 423190 269741 423242 269793
rect 429622 269741 429674 269793
rect 596278 269741 596330 269793
rect 134806 269667 134858 269719
rect 423478 269667 423530 269719
rect 429526 269667 429578 269719
rect 599830 269667 599882 269719
rect 127702 269593 127754 269645
rect 423382 269593 423434 269645
rect 426262 269593 426314 269645
rect 428950 269593 429002 269645
rect 429718 269593 429770 269645
rect 603382 269593 603434 269645
rect 121654 269519 121706 269571
rect 425974 269519 426026 269571
rect 426838 269519 426890 269571
rect 621238 269519 621290 269571
rect 128854 269445 128906 269497
rect 440086 269445 440138 269497
rect 459094 269445 459146 269497
rect 620086 269445 620138 269497
rect 114646 269371 114698 269423
rect 427510 269371 427562 269423
rect 429430 269371 429482 269423
rect 431158 269371 431210 269423
rect 432022 269371 432074 269423
rect 605782 269371 605834 269423
rect 109846 269297 109898 269349
rect 426454 269297 426506 269349
rect 429142 269297 429194 269349
rect 616438 269297 616490 269349
rect 102646 269223 102698 269275
rect 436822 269223 436874 269275
rect 452662 269223 452714 269275
rect 648694 269223 648746 269275
rect 115798 269149 115850 269201
rect 140566 269149 140618 269201
rect 166870 269149 166922 269201
rect 421654 269149 421706 269201
rect 427702 269149 427754 269201
rect 526102 269149 526154 269201
rect 119350 269075 119402 269127
rect 140758 269075 140810 269127
rect 171670 269075 171722 269127
rect 184342 269075 184394 269127
rect 184726 269075 184778 269127
rect 133270 269001 133322 269053
rect 140854 269001 140906 269053
rect 202582 269001 202634 269053
rect 204310 269001 204362 269053
rect 126454 268927 126506 268979
rect 140662 268927 140714 268979
rect 189526 268927 189578 268979
rect 418870 269001 418922 269053
rect 429046 269075 429098 269127
rect 469366 269075 469418 269127
rect 480886 269075 480938 269127
rect 489718 269075 489770 269127
rect 434614 269001 434666 269053
rect 470806 269001 470858 269053
rect 499702 269001 499754 269053
rect 509782 269001 509834 269053
rect 552214 269075 552266 269127
rect 130006 268853 130058 268905
rect 139606 268853 139658 268905
rect 132886 268779 132938 268831
rect 140950 268779 141002 268831
rect 188278 268779 188330 268831
rect 417622 268927 417674 268979
rect 418966 268927 419018 268979
rect 429046 268927 429098 268979
rect 430006 268927 430058 268979
rect 446422 268927 446474 268979
rect 212182 268853 212234 268905
rect 212950 268853 213002 268905
rect 219190 268853 219242 268905
rect 221494 268853 221546 268905
rect 225238 268853 225290 268905
rect 227350 268853 227402 268905
rect 210934 268779 210986 268831
rect 213046 268779 213098 268831
rect 222838 268779 222890 268831
rect 389878 268853 389930 268905
rect 389974 268853 390026 268905
rect 391702 268853 391754 268905
rect 397654 268853 397706 268905
rect 400726 268853 400778 268905
rect 401494 268853 401546 268905
rect 408310 268853 408362 268905
rect 426550 268853 426602 268905
rect 430198 268853 430250 268905
rect 227638 268779 227690 268831
rect 230134 268779 230186 268831
rect 234646 268779 234698 268831
rect 235894 268779 235946 268831
rect 252502 268779 252554 268831
rect 253366 268779 253418 268831
rect 259702 268779 259754 268831
rect 262006 268779 262058 268831
rect 266806 268779 266858 268831
rect 267766 268779 267818 268831
rect 274006 268779 274058 268831
rect 276406 268779 276458 268831
rect 298966 268779 299018 268831
rect 300310 268779 300362 268831
rect 300406 268779 300458 268831
rect 358486 268779 358538 268831
rect 364438 268779 364490 268831
rect 366646 268779 366698 268831
rect 377494 268779 377546 268831
rect 460822 268927 460874 268979
rect 459286 268853 459338 268905
rect 470806 268853 470858 268905
rect 509686 268927 509738 268979
rect 489718 268853 489770 268905
rect 533206 268853 533258 268905
rect 460822 268779 460874 268831
rect 122902 268705 122954 268757
rect 139990 268705 140042 268757
rect 295414 268705 295466 268757
rect 299542 268705 299594 268757
rect 300982 268705 301034 268757
rect 306070 268705 306122 268757
rect 342070 268705 342122 268757
rect 348790 268705 348842 268757
rect 364246 268705 364298 268757
rect 370294 268705 370346 268757
rect 376246 268705 376298 268757
rect 377206 268705 377258 268757
rect 378166 268705 378218 268757
rect 393910 268705 393962 268757
rect 147958 268631 148010 268683
rect 149686 268631 149738 268683
rect 226390 268631 226442 268683
rect 227446 268631 227498 268683
rect 276310 268631 276362 268683
rect 388726 268631 388778 268683
rect 190678 268557 190730 268609
rect 192886 268557 192938 268609
rect 310678 268557 310730 268609
rect 288214 268483 288266 268535
rect 299158 268483 299210 268535
rect 283414 268409 283466 268461
rect 288022 268409 288074 268461
rect 290614 268409 290666 268461
rect 307990 268483 308042 268535
rect 308182 268483 308234 268535
rect 387286 268557 387338 268609
rect 439126 268705 439178 268757
rect 439318 268705 439370 268757
rect 548758 268705 548810 268757
rect 407734 268631 407786 268683
rect 408982 268631 409034 268683
rect 417622 268631 417674 268683
rect 426262 268631 426314 268683
rect 429046 268631 429098 268683
rect 459286 268631 459338 268683
rect 408694 268557 408746 268609
rect 508246 268557 508298 268609
rect 286198 268335 286250 268387
rect 300406 268335 300458 268387
rect 281110 268261 281162 268313
rect 298774 268261 298826 268313
rect 144310 268187 144362 268239
rect 146518 268187 146570 268239
rect 288022 268187 288074 268239
rect 310678 268409 310730 268461
rect 389686 268483 389738 268535
rect 390550 268483 390602 268535
rect 400342 268483 400394 268535
rect 406582 268483 406634 268535
rect 501142 268483 501194 268535
rect 300598 268335 300650 268387
rect 302422 268335 302474 268387
rect 304918 268261 304970 268313
rect 315670 268335 315722 268387
rect 390358 268409 390410 268461
rect 391798 268409 391850 268461
rect 403606 268409 403658 268461
rect 425686 268409 425738 268461
rect 494038 268409 494090 268461
rect 499702 268409 499754 268461
rect 518902 268409 518954 268461
rect 348406 268261 348458 268313
rect 378166 268261 378218 268313
rect 389014 268335 389066 268387
rect 389878 268335 389930 268387
rect 398806 268335 398858 268387
rect 408598 268335 408650 268387
rect 418966 268335 419018 268387
rect 423286 268335 423338 268387
rect 486838 268335 486890 268387
rect 393334 268261 393386 268313
rect 424918 268261 424970 268313
rect 479734 268261 479786 268313
rect 335830 268187 335882 268239
rect 342070 268187 342122 268239
rect 301846 268113 301898 268165
rect 316726 268113 316778 268165
rect 333430 268113 333482 268165
rect 378934 268187 378986 268239
rect 388918 268187 388970 268239
rect 396502 268187 396554 268239
rect 408982 268187 409034 268239
rect 429046 268187 429098 268239
rect 368566 268113 368618 268165
rect 376726 268113 376778 268165
rect 301750 268039 301802 268091
rect 313270 268039 313322 268091
rect 332278 268039 332330 268091
rect 348118 268039 348170 268091
rect 348214 268039 348266 268091
rect 301366 267965 301418 268017
rect 309622 267965 309674 268017
rect 328726 267965 328778 268017
rect 151414 267891 151466 267943
rect 152566 267891 152618 267943
rect 339766 267965 339818 268017
rect 348406 267965 348458 268017
rect 347542 267891 347594 267943
rect 358390 268039 358442 268091
rect 380182 268113 380234 268165
rect 358486 267965 358538 268017
rect 378454 268039 378506 268091
rect 399574 268113 399626 268165
rect 418870 268113 418922 268165
rect 426550 268113 426602 268165
rect 440662 268113 440714 268165
rect 476182 268187 476234 268239
rect 377206 267965 377258 268017
rect 383350 268039 383402 268091
rect 399862 268039 399914 268091
rect 430486 268039 430538 268091
rect 378934 267965 378986 268017
rect 395062 267965 395114 268017
rect 440662 267965 440714 268017
rect 368566 267891 368618 267943
rect 326326 267817 326378 267869
rect 328054 267817 328106 267869
rect 339574 267817 339626 267869
rect 349270 267817 349322 267869
rect 365590 267817 365642 267869
rect 394582 267891 394634 267943
rect 401878 267891 401930 267943
rect 415510 267891 415562 267943
rect 521398 267891 521450 267943
rect 522262 267891 522314 267943
rect 376726 267817 376778 267869
rect 386998 267817 387050 267869
rect 508438 267817 508490 267869
rect 512758 267817 512810 267869
rect 139222 267743 139274 267795
rect 139702 267743 139754 267795
rect 247798 267743 247850 267795
rect 372502 267743 372554 267795
rect 372598 267743 372650 267795
rect 397750 267743 397802 267795
rect 402550 267743 402602 267795
rect 429814 267743 429866 267795
rect 622102 267743 622154 267795
rect 633142 267743 633194 267795
rect 244246 267669 244298 267721
rect 378550 267669 378602 267721
rect 379990 267669 380042 267721
rect 399382 267669 399434 267721
rect 402934 267669 402986 267721
rect 436918 267669 436970 267721
rect 240694 267595 240746 267647
rect 378358 267595 378410 267647
rect 215734 267521 215786 267573
rect 378742 267595 378794 267647
rect 397558 267595 397610 267647
rect 404086 267595 404138 267647
rect 454678 267595 454730 267647
rect 403318 267521 403370 267573
rect 404374 267521 404426 267573
rect 461878 267521 461930 267573
rect 208534 267447 208586 267499
rect 379990 267447 380042 267499
rect 380086 267447 380138 267499
rect 398998 267447 399050 267499
rect 404854 267447 404906 267499
rect 468982 267447 469034 267499
rect 204982 267373 205034 267425
rect 395542 267373 395594 267425
rect 354838 267299 354890 267351
rect 372598 267299 372650 267351
rect 378838 267299 378890 267351
rect 351286 267225 351338 267277
rect 378742 267225 378794 267277
rect 379798 267225 379850 267277
rect 336982 267151 337034 267203
rect 339766 267151 339818 267203
rect 352918 267151 352970 267203
rect 382198 267151 382250 267203
rect 383158 267225 383210 267277
rect 390646 267225 390698 267277
rect 390838 267299 390890 267351
rect 399094 267373 399146 267425
rect 402166 267373 402218 267425
rect 422614 267373 422666 267425
rect 424438 267373 424490 267425
rect 431638 267373 431690 267425
rect 397462 267299 397514 267351
rect 399958 267299 400010 267351
rect 423670 267299 423722 267351
rect 547510 267373 547562 267425
rect 480694 267299 480746 267351
rect 489814 267299 489866 267351
rect 398422 267225 398474 267277
rect 398806 267225 398858 267277
rect 407350 267225 407402 267277
rect 535702 267225 535754 267277
rect 536182 267225 536234 267277
rect 256918 267077 256970 267129
rect 277846 267077 277898 267129
rect 285622 267077 285674 267129
rect 367894 267077 367946 267129
rect 372502 267077 372554 267129
rect 182422 267003 182474 267055
rect 277942 267003 277994 267055
rect 282838 267003 282890 267055
rect 372694 267003 372746 267055
rect 382006 267077 382058 267129
rect 398806 267077 398858 267129
rect 382198 267003 382250 267055
rect 382294 267003 382346 267055
rect 393046 267003 393098 267055
rect 399094 267151 399146 267203
rect 600982 267151 601034 267203
rect 399190 267077 399242 267129
rect 604630 267077 604682 267129
rect 610486 267077 610538 267129
rect 621910 267077 621962 267129
rect 608182 267003 608234 267055
rect 610294 267003 610346 267055
rect 612022 267003 612074 267055
rect 235990 266929 236042 266981
rect 337366 266929 337418 266981
rect 348502 266929 348554 266981
rect 368566 266929 368618 266981
rect 378550 266929 378602 266981
rect 382582 266929 382634 266981
rect 382678 266929 382730 266981
rect 221590 266855 221642 266907
rect 360214 266855 360266 266907
rect 362038 266855 362090 266907
rect 378838 266855 378890 266907
rect 72118 266781 72170 266833
rect 83638 266781 83690 266833
rect 233494 266781 233546 266833
rect 256918 266781 256970 266833
rect 277846 266781 277898 266833
rect 229942 266707 229994 266759
rect 377206 266707 377258 266759
rect 378742 266781 378794 266833
rect 387862 266855 387914 266907
rect 398998 266929 399050 266981
rect 498262 266929 498314 266981
rect 498358 266929 498410 266981
rect 498550 266929 498602 266981
rect 611734 266929 611786 266981
rect 418966 266855 419018 266907
rect 460822 266855 460874 266907
rect 485206 266855 485258 266907
rect 495286 266855 495338 266907
rect 570262 266855 570314 266907
rect 610486 266855 610538 266907
rect 379222 266781 379274 266833
rect 398518 266781 398570 266833
rect 398806 266781 398858 266833
rect 480694 266781 480746 266833
rect 489814 266781 489866 266833
rect 535510 266781 535562 266833
rect 535606 266781 535658 266833
rect 590230 266781 590282 266833
rect 590518 266781 590570 266833
rect 610390 266781 610442 266833
rect 610678 266781 610730 266833
rect 626038 266781 626090 266833
rect 381238 266707 381290 266759
rect 382582 266707 382634 266759
rect 383638 266707 383690 266759
rect 383734 266707 383786 266759
rect 386326 266707 386378 266759
rect 393046 266707 393098 266759
rect 480790 266707 480842 266759
rect 489718 266707 489770 266759
rect 590134 266707 590186 266759
rect 590614 266707 590666 266759
rect 610294 266707 610346 266759
rect 612022 266707 612074 266759
rect 629590 266707 629642 266759
rect 66838 266633 66890 266685
rect 80566 266633 80618 266685
rect 135958 266633 136010 266685
rect 282262 266633 282314 266685
rect 289270 266633 289322 266685
rect 377494 266633 377546 266685
rect 378550 266633 378602 266685
rect 386710 266633 386762 266685
rect 418966 266633 419018 266685
rect 460822 266633 460874 266685
rect 535510 266633 535562 266685
rect 538486 266633 538538 266685
rect 561526 266633 561578 266685
rect 570262 266633 570314 266685
rect 125302 266559 125354 266611
rect 277846 266559 277898 266611
rect 286582 266559 286634 266611
rect 378646 266559 378698 266611
rect 378838 266559 378890 266611
rect 397462 266559 397514 266611
rect 397654 266559 397706 266611
rect 535798 266559 535850 266611
rect 535990 266559 536042 266611
rect 636694 266559 636746 266611
rect 194326 266485 194378 266537
rect 373078 266485 373130 266537
rect 374806 266485 374858 266537
rect 383446 266485 383498 266537
rect 201334 266411 201386 266463
rect 378070 266411 378122 266463
rect 378166 266411 378218 266463
rect 383350 266411 383402 266463
rect 385750 266485 385802 266537
rect 393430 266485 393482 266537
rect 535702 266485 535754 266537
rect 545686 266485 545738 266537
rect 640246 266485 640298 266537
rect 82486 266337 82538 266389
rect 282550 266337 282602 266389
rect 282646 266337 282698 266389
rect 383830 266411 383882 266463
rect 643894 266411 643946 266463
rect 383542 266337 383594 266389
rect 393430 266337 393482 266389
rect 398806 266337 398858 266389
rect 647446 266337 647498 266389
rect 254902 266263 254954 266315
rect 374806 266263 374858 266315
rect 374902 266263 374954 266315
rect 394870 266263 394922 266315
rect 408118 266263 408170 266315
rect 427702 266263 427754 266315
rect 480790 266263 480842 266315
rect 489718 266263 489770 266315
rect 498454 266263 498506 266315
rect 535414 266263 535466 266315
rect 541750 266263 541802 266315
rect 542806 266263 542858 266315
rect 258550 266189 258602 266241
rect 378550 266189 378602 266241
rect 262102 266115 262154 266167
rect 287926 266041 287978 266093
rect 378742 266041 378794 266093
rect 272758 265967 272810 266019
rect 348502 265967 348554 266019
rect 368566 265967 368618 266019
rect 378166 265967 378218 266019
rect 378838 265967 378890 266019
rect 286870 265893 286922 265945
rect 379414 266189 379466 266241
rect 399190 266189 399242 266241
rect 405142 266189 405194 266241
rect 430486 266189 430538 266241
rect 485206 266189 485258 266241
rect 495286 266189 495338 266241
rect 535702 266189 535754 266241
rect 545686 266189 545738 266241
rect 379030 266115 379082 266167
rect 383158 266115 383210 266167
rect 383350 266115 383402 266167
rect 388534 266115 388586 266167
rect 389014 266115 389066 266167
rect 392278 266115 392330 266167
rect 541462 266115 541514 266167
rect 542038 266115 542090 266167
rect 381622 266041 381674 266093
rect 622486 266041 622538 266093
rect 379126 265967 379178 266019
rect 383446 265967 383498 266019
rect 398518 265967 398570 266019
rect 597526 265967 597578 266019
rect 383062 265893 383114 265945
rect 386998 265893 387050 265945
rect 396694 265893 396746 265945
rect 265654 265819 265706 265871
rect 282742 265819 282794 265871
rect 394102 265819 394154 265871
rect 279958 265745 280010 265797
rect 378646 265745 378698 265797
rect 384214 265745 384266 265797
rect 398806 265745 398858 265797
rect 287158 265671 287210 265723
rect 392854 265671 392906 265723
rect 427510 265671 427562 265723
rect 438646 265671 438698 265723
rect 287926 265597 287978 265649
rect 328246 265597 328298 265649
rect 429334 265597 429386 265649
rect 327862 265523 327914 265575
rect 429430 265523 429482 265575
rect 287062 265449 287114 265501
rect 375190 265449 375242 265501
rect 286774 265375 286826 265427
rect 386902 265449 386954 265501
rect 375382 265375 375434 265427
rect 389590 265375 389642 265427
rect 389782 265375 389834 265427
rect 593878 265375 593930 265427
rect 329302 265301 329354 265353
rect 424822 265301 424874 265353
rect 294166 265227 294218 265279
rect 390742 265227 390794 265279
rect 405910 265227 405962 265279
rect 423286 265227 423338 265279
rect 301270 265153 301322 265205
rect 329878 265079 329930 265131
rect 374902 265079 374954 265131
rect 378070 265153 378122 265205
rect 378550 265153 378602 265205
rect 378646 265153 378698 265205
rect 389110 265153 389162 265205
rect 391894 265153 391946 265205
rect 394582 265153 394634 265205
rect 398902 265153 398954 265205
rect 283126 265005 283178 265057
rect 425590 265005 425642 265057
rect 429238 265005 429290 265057
rect 443446 265005 443498 265057
rect 251350 264931 251402 264983
rect 386038 264931 386090 264983
rect 421654 264931 421706 264983
rect 432502 264931 432554 264983
rect 271606 264857 271658 264909
rect 318262 264857 318314 264909
rect 325078 264857 325130 264909
rect 329398 264857 329450 264909
rect 329494 264857 329546 264909
rect 344374 264857 344426 264909
rect 359542 264857 359594 264909
rect 499894 264857 499946 264909
rect 267958 264783 268010 264835
rect 318070 264783 318122 264835
rect 264502 264709 264554 264761
rect 329206 264783 329258 264835
rect 339958 264783 340010 264835
rect 359926 264783 359978 264835
rect 506902 264783 506954 264835
rect 257302 264635 257354 264687
rect 318166 264635 318218 264687
rect 260854 264561 260906 264613
rect 333718 264709 333770 264761
rect 340342 264709 340394 264761
rect 360982 264709 361034 264761
rect 524950 264709 525002 264761
rect 318454 264635 318506 264687
rect 339574 264635 339626 264687
rect 360598 264635 360650 264687
rect 517750 264635 517802 264687
rect 318646 264561 318698 264613
rect 333718 264561 333770 264613
rect 253750 264487 253802 264539
rect 339286 264561 339338 264613
rect 361366 264561 361418 264613
rect 532054 264561 532106 264613
rect 335254 264487 335306 264539
rect 356182 264487 356234 264539
rect 361750 264487 361802 264539
rect 539158 264487 539210 264539
rect 283318 264413 283370 264465
rect 371446 264413 371498 264465
rect 374230 264413 374282 264465
rect 558262 264413 558314 264465
rect 250102 264339 250154 264391
rect 338902 264339 338954 264391
rect 42262 264265 42314 264317
rect 53302 264265 53354 264317
rect 246646 264265 246698 264317
rect 338518 264265 338570 264317
rect 338614 264265 338666 264317
rect 347350 264339 347402 264391
rect 362134 264339 362186 264391
rect 546358 264339 546410 264391
rect 243094 264191 243146 264243
rect 338134 264191 338186 264243
rect 341686 264265 341738 264317
rect 375382 264265 375434 264317
rect 568918 264265 568970 264317
rect 214486 264117 214538 264169
rect 335254 264117 335306 264169
rect 335350 264117 335402 264169
rect 338038 264117 338090 264169
rect 196726 264043 196778 264095
rect 312406 264043 312458 264095
rect 318454 264043 318506 264095
rect 339766 264191 339818 264243
rect 368662 264191 368714 264243
rect 374998 264191 375050 264243
rect 565366 264191 565418 264243
rect 200182 263969 200234 264021
rect 329494 263969 329546 264021
rect 329590 263969 329642 264021
rect 338230 263969 338282 264021
rect 207382 263895 207434 263947
rect 352150 264117 352202 264169
rect 375670 264117 375722 264169
rect 572470 264117 572522 264169
rect 340534 264043 340586 264095
rect 360022 264043 360074 264095
rect 376054 264043 376106 264095
rect 576118 264043 576170 264095
rect 338422 263969 338474 264021
rect 346486 263969 346538 264021
rect 347734 263969 347786 264021
rect 368470 263969 368522 264021
rect 376438 263969 376490 264021
rect 579670 263969 579722 264021
rect 338710 263895 338762 263947
rect 340726 263895 340778 263947
rect 377590 263895 377642 263947
rect 586774 263895 586826 263947
rect 203734 263821 203786 263873
rect 348502 263821 348554 263873
rect 352534 263821 352586 263873
rect 375094 263821 375146 263873
rect 376822 263821 376874 263873
rect 583126 263821 583178 263873
rect 239446 263747 239498 263799
rect 337750 263747 337802 263799
rect 337846 263747 337898 263799
rect 592726 263747 592778 263799
rect 228790 263673 228842 263725
rect 232342 263599 232394 263651
rect 314326 263599 314378 263651
rect 318070 263673 318122 263725
rect 330070 263599 330122 263651
rect 330166 263599 330218 263651
rect 339670 263673 339722 263725
rect 624790 263673 624842 263725
rect 42262 263525 42314 263577
rect 53398 263525 53450 263577
rect 275158 263525 275210 263577
rect 318454 263525 318506 263577
rect 318550 263525 318602 263577
rect 329590 263525 329642 263577
rect 329686 263525 329738 263577
rect 333238 263525 333290 263577
rect 334870 263525 334922 263577
rect 335350 263599 335402 263651
rect 628438 263599 628490 263651
rect 341110 263525 341162 263577
rect 318166 263451 318218 263503
rect 342550 263451 342602 263503
rect 285814 263377 285866 263429
rect 342838 263377 342890 263429
rect 278710 263303 278762 263355
rect 342166 263303 342218 263355
rect 282934 263229 282986 263281
rect 318166 263229 318218 263281
rect 319126 263229 319178 263281
rect 333142 263229 333194 263281
rect 333238 263229 333290 263281
rect 368566 263525 368618 263577
rect 383158 263525 383210 263577
rect 386806 263525 386858 263577
rect 423574 263525 423626 263577
rect 430390 263525 430442 263577
rect 535702 263525 535754 263577
rect 536182 263525 536234 263577
rect 359158 263451 359210 263503
rect 492790 263451 492842 263503
rect 358774 263377 358826 263429
rect 485590 263377 485642 263429
rect 358390 263303 358442 263355
rect 478582 263303 478634 263355
rect 358006 263229 358058 263281
rect 474934 263229 474986 263281
rect 289462 263155 289514 263207
rect 343318 263155 343370 263207
rect 357718 263155 357770 263207
rect 467830 263155 467882 263207
rect 124054 263007 124106 263059
rect 141142 263007 141194 263059
rect 149398 263007 149450 263059
rect 141142 262859 141194 262911
rect 149398 262859 149450 262911
rect 221686 262933 221738 262985
rect 221782 262933 221834 262985
rect 236182 263081 236234 263133
rect 262102 263081 262154 263133
rect 262294 263081 262346 263133
rect 236278 263007 236330 263059
rect 293014 263081 293066 263133
rect 343702 263081 343754 263133
rect 357334 263081 357386 263133
rect 460726 263081 460778 263133
rect 325462 263007 325514 263059
rect 328054 263007 328106 263059
rect 333526 263007 333578 263059
rect 333622 263007 333674 263059
rect 331510 262933 331562 262985
rect 368566 263007 368618 263059
rect 427798 263007 427850 263059
rect 318262 262859 318314 262911
rect 341494 262859 341546 262911
rect 429526 262933 429578 262985
rect 429622 262859 429674 262911
rect 296566 262785 296618 262837
rect 344086 262785 344138 262837
rect 356950 262785 357002 262837
rect 453526 262785 453578 262837
rect 286390 262711 286442 262763
rect 369046 262711 369098 262763
rect 383446 262711 383498 262763
rect 384022 262711 384074 262763
rect 426262 262711 426314 262763
rect 434902 262711 434954 262763
rect 300118 262637 300170 262689
rect 344758 262637 344810 262689
rect 355798 262637 355850 262689
rect 435670 262637 435722 262689
rect 303670 262563 303722 262615
rect 345142 262563 345194 262615
rect 355510 262563 355562 262615
rect 428566 262563 428618 262615
rect 310870 262489 310922 262541
rect 345910 262489 345962 262541
rect 355126 262489 355178 262541
rect 421462 262489 421514 262541
rect 426454 262489 426506 262541
rect 437494 262489 437546 262541
rect 307222 262415 307274 262467
rect 345526 262415 345578 262467
rect 354742 262415 354794 262467
rect 414358 262415 414410 262467
rect 312022 262341 312074 262393
rect 366838 262341 366890 262393
rect 383062 262341 383114 262393
rect 397654 262341 397706 262393
rect 42838 262267 42890 262319
rect 58966 262267 59018 262319
rect 314422 262267 314474 262319
rect 346294 262267 346346 262319
rect 353974 262267 354026 262319
rect 391798 262267 391850 262319
rect 314326 262193 314378 262245
rect 334102 262193 334154 262245
rect 301846 262119 301898 262171
rect 302038 262119 302090 262171
rect 321526 262119 321578 262171
rect 346966 262193 347018 262245
rect 353686 262193 353738 262245
rect 388918 262193 388970 262245
rect 337078 262119 337130 262171
rect 646294 262119 646346 262171
rect 256150 262045 256202 262097
rect 296950 262045 297002 262097
rect 310294 262045 310346 262097
rect 466582 262045 466634 262097
rect 249046 261971 249098 262023
rect 296566 261971 296618 262023
rect 311350 261971 311402 262023
rect 477334 261971 477386 262023
rect 231190 261897 231242 261949
rect 175222 261823 175274 261875
rect 234070 261823 234122 261875
rect 168022 261749 168074 261801
rect 233206 261749 233258 261801
rect 245398 261897 245450 261949
rect 296182 261897 296234 261949
rect 310102 261897 310154 261949
rect 473782 261897 473834 261949
rect 238294 261823 238346 261875
rect 295798 261823 295850 261875
rect 311638 261823 311690 261875
rect 484438 261823 484490 261875
rect 277078 261749 277130 261801
rect 312022 261749 312074 261801
rect 491638 261749 491690 261801
rect 303190 261675 303242 261727
rect 334582 261675 334634 261727
rect 373846 261675 373898 261727
rect 554614 261675 554666 261727
rect 303958 261601 304010 261653
rect 348886 261601 348938 261653
rect 353302 261601 353354 261653
rect 366262 261601 366314 261653
rect 374614 261601 374666 261653
rect 561814 261601 561866 261653
rect 185878 261527 185930 261579
rect 201622 261527 201674 261579
rect 206134 261527 206186 261579
rect 305014 261527 305066 261579
rect 312790 261527 312842 261579
rect 191926 261453 191978 261505
rect 288790 261453 288842 261505
rect 313558 261453 313610 261505
rect 326326 261527 326378 261579
rect 498838 261527 498890 261579
rect 80662 261379 80714 261431
rect 83542 261379 83594 261431
rect 199030 261379 199082 261431
rect 299926 261379 299978 261431
rect 193078 261305 193130 261357
rect 326038 261379 326090 261431
rect 505846 261453 505898 261505
rect 516502 261379 516554 261431
rect 195478 261231 195530 261283
rect 297334 261231 297386 261283
rect 302806 261231 302858 261283
rect 331030 261305 331082 261357
rect 354262 261305 354314 261357
rect 366166 261305 366218 261357
rect 366262 261305 366314 261357
rect 389302 261305 389354 261357
rect 424246 261305 424298 261357
rect 430870 261305 430922 261357
rect 314518 261231 314570 261283
rect 177622 261157 177674 261209
rect 288886 261157 288938 261209
rect 302614 261157 302666 261209
rect 323926 261157 323978 261209
rect 324118 261231 324170 261283
rect 523702 261231 523754 261283
rect 530902 261157 530954 261209
rect 181270 261083 181322 261135
rect 302422 261083 302474 261135
rect 314614 261083 314666 261135
rect 538006 261083 538058 261135
rect 170422 261009 170474 261061
rect 302518 261009 302570 261061
rect 313846 261009 313898 261061
rect 324118 261009 324170 261061
rect 326422 261009 326474 261061
rect 549814 261009 549866 261061
rect 279478 260935 279530 260987
rect 299446 260935 299498 260987
rect 312406 260935 312458 260987
rect 326326 260935 326378 260987
rect 326806 260935 326858 260987
rect 553462 260935 553514 260987
rect 149110 260861 149162 260913
rect 305494 260861 305546 260913
rect 305686 260861 305738 260913
rect 373558 260861 373610 260913
rect 380470 260861 380522 260913
rect 615382 260861 615434 260913
rect 138358 260713 138410 260765
rect 303574 260787 303626 260839
rect 341782 260787 341834 260839
rect 341878 260787 341930 260839
rect 574870 260787 574922 260839
rect 305590 260713 305642 260765
rect 305782 260713 305834 260765
rect 380758 260713 380810 260765
rect 380854 260713 380906 260765
rect 618838 260713 618890 260765
rect 131254 260639 131306 260691
rect 198742 260639 198794 260691
rect 279382 260639 279434 260691
rect 299446 260639 299498 260691
rect 299638 260639 299690 260691
rect 304726 260639 304778 260691
rect 218038 260565 218090 260617
rect 218710 260565 218762 260617
rect 218806 260565 218858 260617
rect 263254 260565 263306 260617
rect 297718 260565 297770 260617
rect 308758 260639 308810 260691
rect 313270 260639 313322 260691
rect 328630 260639 328682 260691
rect 571318 260639 571370 260691
rect 363190 260565 363242 260617
rect 373462 260565 373514 260617
rect 521974 260565 522026 260617
rect 270358 260491 270410 260543
rect 298006 260491 298058 260543
rect 310198 260491 310250 260543
rect 459478 260491 459530 260543
rect 277558 260417 277610 260469
rect 298390 260417 298442 260469
rect 309814 260417 309866 260469
rect 452374 260417 452426 260469
rect 216790 260343 216842 260395
rect 218806 260343 218858 260395
rect 220438 260343 220490 260395
rect 313174 260343 313226 260395
rect 313270 260343 313322 260395
rect 434518 260343 434570 260395
rect 213334 260269 213386 260321
rect 309046 260269 309098 260321
rect 309430 260269 309482 260321
rect 445270 260269 445322 260321
rect 269206 260195 269258 260247
rect 388246 260195 388298 260247
rect 403702 260195 403754 260247
rect 447670 260195 447722 260247
rect 156214 260121 156266 260173
rect 305398 260121 305450 260173
rect 308374 260121 308426 260173
rect 427414 260121 427466 260173
rect 431158 260121 431210 260173
rect 443254 260121 443306 260173
rect 145558 260047 145610 260099
rect 305302 260047 305354 260099
rect 307990 260047 308042 260099
rect 420214 260047 420266 260099
rect 426358 260047 426410 260099
rect 436054 260047 436106 260099
rect 307222 259973 307274 260025
rect 307606 259899 307658 259951
rect 405526 259973 405578 260025
rect 424918 259973 424970 260025
rect 432790 259973 432842 260025
rect 443158 259973 443210 260025
rect 306934 259825 306986 259877
rect 406006 259899 406058 259951
rect 306550 259751 306602 259803
rect 395254 259751 395306 259803
rect 306166 259677 306218 259729
rect 388150 259677 388202 259729
rect 402358 259677 402410 259729
rect 408790 259825 408842 259877
rect 427894 259825 427946 259877
rect 406294 259751 406346 259803
rect 425686 259751 425738 259803
rect 413110 259677 413162 259729
rect 304342 259603 304394 259655
rect 355990 259603 356042 259655
rect 356566 259603 356618 259655
rect 430006 259603 430058 259655
rect 286006 259529 286058 259581
rect 354262 259529 354314 259581
rect 354454 259529 354506 259581
rect 407158 259529 407210 259581
rect 286678 259455 286730 259507
rect 369430 259455 369482 259507
rect 377878 259455 377930 259507
rect 590326 259455 590378 259507
rect 286102 259381 286154 259433
rect 370870 259381 370922 259433
rect 378358 259381 378410 259433
rect 282454 259307 282506 259359
rect 369046 259307 369098 259359
rect 378262 259307 378314 259359
rect 379126 259307 379178 259359
rect 383638 259381 383690 259433
rect 385270 259381 385322 259433
rect 384886 259307 384938 259359
rect 389590 259307 389642 259359
rect 390070 259307 390122 259359
rect 284566 259233 284618 259285
rect 425014 259233 425066 259285
rect 305302 259159 305354 259211
rect 429814 259159 429866 259211
rect 305398 259085 305450 259137
rect 429718 259085 429770 259137
rect 302422 259011 302474 259063
rect 433846 259159 433898 259211
rect 440566 259159 440618 259211
rect 445654 259159 445706 259211
rect 430102 259085 430154 259137
rect 447862 259085 447914 259137
rect 447958 259085 448010 259137
rect 451894 259085 451946 259137
rect 435958 259011 436010 259063
rect 449398 259011 449450 259063
rect 305494 258937 305546 258989
rect 430486 258937 430538 258989
rect 433462 258937 433514 258989
rect 447958 258937 448010 258989
rect 302518 258863 302570 258915
rect 432694 258863 432746 258915
rect 288886 258789 288938 258841
rect 433462 258789 433514 258841
rect 443254 258789 443306 258841
rect 452950 258937 453002 258989
rect 282262 258715 282314 258767
rect 418774 258715 418826 258767
rect 418870 258715 418922 258767
rect 443062 258715 443114 258767
rect 443158 258715 443210 258767
rect 451126 258715 451178 258767
rect 277846 258641 277898 258693
rect 439702 258641 439754 258693
rect 277942 258567 277994 258619
rect 430102 258567 430154 258619
rect 430198 258567 430250 258619
rect 447094 258567 447146 258619
rect 234070 258493 234122 258545
rect 445270 258493 445322 258545
rect 233206 258419 233258 258471
rect 444502 258419 444554 258471
rect 201622 258345 201674 258397
rect 446710 258345 446762 258397
rect 161014 258271 161066 258323
rect 443734 258271 443786 258323
rect 153814 258197 153866 258249
rect 418870 258197 418922 258249
rect 143158 258123 143210 258175
rect 441526 258197 441578 258249
rect 423382 258123 423434 258175
rect 427990 258123 428042 258175
rect 428182 258123 428234 258175
rect 441238 258123 441290 258175
rect 83638 258049 83690 258101
rect 96310 258049 96362 258101
rect 118102 258049 118154 258101
rect 438838 258049 438890 258101
rect 106198 257975 106250 258027
rect 437110 257975 437162 258027
rect 437206 257975 437258 258027
rect 450358 257975 450410 258027
rect 99190 257901 99242 257953
rect 436438 257901 436490 257953
rect 110998 257827 111050 257879
rect 449590 257827 449642 257879
rect 103894 257753 103946 257805
rect 448918 257753 448970 257805
rect 455446 257753 455498 257805
rect 456790 257753 456842 257805
rect 460822 257753 460874 257805
rect 462838 257753 462890 257805
rect 469462 257753 469514 257805
rect 471094 257753 471146 257805
rect 480982 257753 481034 257805
rect 482998 257753 483050 257805
rect 486838 257753 486890 257805
rect 488950 257753 489002 257805
rect 492694 257753 492746 257805
rect 494806 257753 494858 257805
rect 495382 257753 495434 257805
rect 497302 257753 497354 257805
rect 501238 257753 501290 257805
rect 503158 257753 503210 257805
rect 507094 257753 507146 257805
rect 509206 257753 509258 257805
rect 509782 257753 509834 257805
rect 511606 257753 511658 257805
rect 512854 257753 512906 257805
rect 514006 257753 514058 257805
rect 527062 257753 527114 257805
rect 528214 257753 528266 257805
rect 533014 257753 533066 257805
rect 535318 257753 535370 257805
rect 541654 257753 541706 257805
rect 543670 257753 543722 257805
rect 282262 257679 282314 257731
rect 284374 257679 284426 257731
rect 305590 257679 305642 257731
rect 429046 257679 429098 257731
rect 430102 257679 430154 257731
rect 445942 257679 445994 257731
rect 512662 257679 512714 257731
rect 515158 257679 515210 257731
rect 527158 257679 527210 257731
rect 529462 257679 529514 257731
rect 309142 257605 309194 257657
rect 428278 257605 428330 257657
rect 428470 257605 428522 257657
rect 446326 257605 446378 257657
rect 325462 257235 325514 257287
rect 427606 257531 427658 257583
rect 430294 257531 430346 257583
rect 448534 257531 448586 257583
rect 331894 257457 331946 257509
rect 333622 257457 333674 257509
rect 334870 257457 334922 257509
rect 339670 257457 339722 257509
rect 331126 257383 331178 257435
rect 426838 257457 426890 257509
rect 426934 257457 426986 257509
rect 330742 257309 330794 257361
rect 427222 257383 427274 257435
rect 427894 257457 427946 257509
rect 444118 257457 444170 257509
rect 444886 257383 444938 257435
rect 351094 257309 351146 257361
rect 357430 257309 357482 257361
rect 358486 257309 358538 257361
rect 426454 257309 426506 257361
rect 333526 257235 333578 257287
rect 394486 257235 394538 257287
rect 401110 257235 401162 257287
rect 404758 257235 404810 257287
rect 406966 257235 407018 257287
rect 408694 257235 408746 257287
rect 409174 257235 409226 257287
rect 423670 257235 423722 257287
rect 425974 257235 426026 257287
rect 438934 257235 438986 257287
rect 333142 257161 333194 257213
rect 393718 257161 393770 257213
rect 427318 257161 427370 257213
rect 442678 257161 442730 257213
rect 331222 257087 331274 257139
rect 337846 257087 337898 257139
rect 350710 257087 350762 257139
rect 353590 257087 353642 257139
rect 360022 257087 360074 257139
rect 396310 257087 396362 257139
rect 418774 257087 418826 257139
rect 440854 257087 440906 257139
rect 346582 257013 346634 257065
rect 349942 257013 349994 257065
rect 378742 257013 378794 257065
rect 379222 257013 379274 257065
rect 383062 257013 383114 257065
rect 393046 257013 393098 257065
rect 423190 257013 423242 257065
rect 440470 257013 440522 257065
rect 342934 256939 342986 256991
rect 349558 256939 349610 256991
rect 351766 256939 351818 256991
rect 364342 256939 364394 256991
rect 368662 256939 368714 256991
rect 322294 256865 322346 256917
rect 327190 256865 327242 256917
rect 330934 256865 330986 256917
rect 282550 256791 282602 256843
rect 325654 256791 325706 256843
rect 329014 256791 329066 256843
rect 341878 256791 341930 256843
rect 366838 256865 366890 256917
rect 378454 256865 378506 256917
rect 358486 256791 358538 256843
rect 365590 256791 365642 256843
rect 285910 256717 285962 256769
rect 366838 256717 366890 256769
rect 367798 256791 367850 256843
rect 378550 256791 378602 256843
rect 378838 256939 378890 256991
rect 388726 256939 388778 256991
rect 423478 256939 423530 256991
rect 428662 256939 428714 256991
rect 428950 256939 429002 256991
rect 441910 256939 441962 256991
rect 425782 256865 425834 256917
rect 428182 256865 428234 256917
rect 429718 256865 429770 256917
rect 431254 256865 431306 256917
rect 395926 256791 395978 256843
rect 425878 256791 425930 256843
rect 437878 256791 437930 256843
rect 368374 256717 368426 256769
rect 368470 256717 368522 256769
rect 383158 256717 383210 256769
rect 286486 256643 286538 256695
rect 365878 256643 365930 256695
rect 367126 256643 367178 256695
rect 391606 256717 391658 256769
rect 452278 256717 452330 256769
rect 438262 256643 438314 256695
rect 285814 256569 285866 256621
rect 365590 256569 365642 256621
rect 285238 256495 285290 256547
rect 367510 256569 367562 256621
rect 367606 256569 367658 256621
rect 442294 256569 442346 256621
rect 285142 256421 285194 256473
rect 283606 256347 283658 256399
rect 300790 256347 300842 256399
rect 369814 256421 369866 256473
rect 371446 256421 371498 256473
rect 383638 256495 383690 256547
rect 383734 256495 383786 256547
rect 451510 256495 451562 256547
rect 378550 256421 378602 256473
rect 383062 256421 383114 256473
rect 393046 256421 393098 256473
rect 450070 256421 450122 256473
rect 310870 256347 310922 256399
rect 370198 256347 370250 256399
rect 370294 256347 370346 256399
rect 450742 256347 450794 256399
rect 640726 256347 640778 256399
rect 679702 256347 679754 256399
rect 310966 256273 311018 256325
rect 322390 256273 322442 256325
rect 322582 256273 322634 256325
rect 637654 256273 637706 256325
rect 288886 256199 288938 256251
rect 322486 256199 322538 256251
rect 322678 256199 322730 256251
rect 630742 256199 630794 256251
rect 300406 256125 300458 256177
rect 310390 256125 310442 256177
rect 282646 256051 282698 256103
rect 293110 256051 293162 256103
rect 293206 256051 293258 256103
rect 422422 256125 422474 256177
rect 495286 256125 495338 256177
rect 508438 256125 508490 256177
rect 310582 256051 310634 256103
rect 362806 256051 362858 256103
rect 285334 255977 285386 256029
rect 363190 255977 363242 256029
rect 259318 255903 259370 255955
rect 141142 255829 141194 255881
rect 60598 255533 60650 255585
rect 80662 255681 80714 255733
rect 106678 255681 106730 255733
rect 118102 255681 118154 255733
rect 138166 255681 138218 255733
rect 141142 255681 141194 255733
rect 178582 255755 178634 255807
rect 178678 255755 178730 255807
rect 218422 255755 218474 255807
rect 218806 255755 218858 255807
rect 284086 255903 284138 255955
rect 300406 255903 300458 255955
rect 300502 255903 300554 255955
rect 310582 255903 310634 255955
rect 310918 255903 310970 255955
rect 363958 255903 364010 255955
rect 421558 255903 421610 255955
rect 424438 255903 424490 255955
rect 288022 255829 288074 255881
rect 300694 255755 300746 255807
rect 300886 255829 300938 255881
rect 365398 255829 365450 255881
rect 423478 255829 423530 255881
rect 423862 255755 423914 255807
rect 218902 255681 218954 255733
rect 86710 255607 86762 255659
rect 106486 255607 106538 255659
rect 293110 255681 293162 255733
rect 300502 255681 300554 255733
rect 300790 255681 300842 255733
rect 541462 255755 541514 255807
rect 541846 255755 541898 255807
rect 259222 255607 259274 255659
rect 289462 255607 289514 255659
rect 322294 255607 322346 255659
rect 322390 255607 322442 255659
rect 324214 255607 324266 255659
rect 443542 255681 443594 255733
rect 443638 255681 443690 255733
rect 43606 255459 43658 255511
rect 60502 255459 60554 255511
rect 218902 255459 218954 255511
rect 288598 255533 288650 255585
rect 310774 255533 310826 255585
rect 310870 255533 310922 255585
rect 337270 255533 337322 255585
rect 423382 255607 423434 255659
rect 490966 255681 491018 255733
rect 501142 255681 501194 255733
rect 469366 255607 469418 255659
rect 538486 255607 538538 255659
rect 570166 255681 570218 255733
rect 590518 255681 590570 255733
rect 601942 255681 601994 255733
rect 622006 255681 622058 255733
rect 630646 255681 630698 255733
rect 570358 255607 570410 255659
rect 590326 255607 590378 255659
rect 630838 255607 630890 255659
rect 642262 255607 642314 255659
rect 662326 255607 662378 255659
rect 671062 255681 671114 255733
rect 286294 255459 286346 255511
rect 363574 255459 363626 255511
rect 469366 255459 469418 255511
rect 490966 255533 491018 255585
rect 301078 255385 301130 255437
rect 364246 255385 364298 255437
rect 283222 255311 283274 255363
rect 364630 255311 364682 255363
rect 284182 255237 284234 255289
rect 365014 255237 365066 255289
rect 518422 255237 518474 255289
rect 519862 255237 519914 255289
rect 286966 255163 287018 255215
rect 367990 255163 368042 255215
rect 287830 255089 287882 255141
rect 366454 255089 366506 255141
rect 283414 255015 283466 255067
rect 83542 254941 83594 254993
rect 112150 254941 112202 254993
rect 277078 254941 277130 254993
rect 293590 254941 293642 254993
rect 368662 255015 368714 255067
rect 388726 255015 388778 255067
rect 391510 255015 391562 255067
rect 319798 254941 319850 254993
rect 440758 254941 440810 254993
rect 65206 254867 65258 254919
rect 200278 254867 200330 254919
rect 288118 254867 288170 254919
rect 319894 254867 319946 254919
rect 321622 254867 321674 254919
rect 443638 254867 443690 254919
rect 295318 254793 295370 254845
rect 320854 254793 320906 254845
rect 322390 254793 322442 254845
rect 443542 254793 443594 254845
rect 316822 254719 316874 254771
rect 440662 254719 440714 254771
rect 285430 254645 285482 254697
rect 414358 254645 414410 254697
rect 285526 254571 285578 254623
rect 412150 254571 412202 254623
rect 282934 254497 282986 254549
rect 413974 254497 414026 254549
rect 283990 254423 284042 254475
rect 301078 254423 301130 254475
rect 310102 254423 310154 254475
rect 310966 254423 311018 254475
rect 316054 254423 316106 254475
rect 446422 254423 446474 254475
rect 318262 254349 318314 254401
rect 445366 254349 445418 254401
rect 317590 254275 317642 254327
rect 444310 254275 444362 254327
rect 284278 254201 284330 254253
rect 298294 254201 298346 254253
rect 315382 254201 315434 254253
rect 446422 254201 446474 254253
rect 287254 254127 287306 254179
rect 421366 254127 421418 254179
rect 287350 254053 287402 254105
rect 422038 254053 422090 254105
rect 284854 253979 284906 254031
rect 420214 253979 420266 254031
rect 287158 253905 287210 253957
rect 423190 253905 423242 253957
rect 285718 253831 285770 253883
rect 290998 253831 291050 253883
rect 298294 253831 298346 253883
rect 420598 253831 420650 253883
rect 288310 253757 288362 253809
rect 322486 253757 322538 253809
rect 322582 253757 322634 253809
rect 338326 253757 338378 253809
rect 351382 253757 351434 253809
rect 360790 253757 360842 253809
rect 285046 253683 285098 253735
rect 422806 253683 422858 253735
rect 284950 253609 285002 253661
rect 290902 253609 290954 253661
rect 290998 253609 291050 253661
rect 362422 253609 362474 253661
rect 204406 253535 204458 253587
rect 316726 253535 316778 253587
rect 322486 253535 322538 253587
rect 323062 253535 323114 253587
rect 338326 253535 338378 253587
rect 495286 253535 495338 253587
rect 287638 253461 287690 253513
rect 367222 253461 367274 253513
rect 288502 253387 288554 253439
rect 508342 253387 508394 253439
rect 674806 253387 674858 253439
rect 676822 253387 676874 253439
rect 287926 253313 287978 253365
rect 370582 253313 370634 253365
rect 283030 253239 283082 253291
rect 300886 253239 300938 253291
rect 282838 253165 282890 253217
rect 371254 253165 371306 253217
rect 418006 253165 418058 253217
rect 440278 253165 440330 253217
rect 140182 253091 140234 253143
rect 141526 253091 141578 253143
rect 287446 253091 287498 253143
rect 372406 253091 372458 253143
rect 416950 253091 417002 253143
rect 446422 253091 446474 253143
rect 287734 253017 287786 253069
rect 371638 253017 371690 253069
rect 423574 253017 423626 253069
rect 112150 252943 112202 252995
rect 142486 252943 142538 252995
rect 287542 252943 287594 252995
rect 372742 252943 372794 252995
rect 388438 252943 388490 252995
rect 392998 252943 393050 252995
rect 445366 252943 445418 252995
rect 96310 252869 96362 252921
rect 141142 252869 141194 252921
rect 287830 252869 287882 252921
rect 372022 252869 372074 252921
rect 416566 252869 416618 252921
rect 444982 252869 445034 252921
rect 446230 252869 446282 252921
rect 80854 252795 80906 252847
rect 146806 252795 146858 252847
rect 284374 252795 284426 252847
rect 411382 252795 411434 252847
rect 417286 252795 417338 252847
rect 67606 252721 67658 252773
rect 146902 252721 146954 252773
rect 45334 252647 45386 252699
rect 200374 252647 200426 252699
rect 45046 252573 45098 252625
rect 200182 252573 200234 252625
rect 45430 252499 45482 252551
rect 200566 252499 200618 252551
rect 44854 252425 44906 252477
rect 200470 252425 200522 252477
rect 45238 252351 45290 252403
rect 204502 252351 204554 252403
rect 45142 252277 45194 252329
rect 204694 252277 204746 252329
rect 44950 252203 45002 252255
rect 204886 252203 204938 252255
rect 44758 252129 44810 252181
rect 204790 252129 204842 252181
rect 44566 252055 44618 252107
rect 204598 252055 204650 252107
rect 44662 251981 44714 252033
rect 204214 251981 204266 252033
rect 675382 251167 675434 251219
rect 283318 251093 283370 251145
rect 283702 251093 283754 251145
rect 283126 250945 283178 250997
rect 283318 250945 283370 250997
rect 675382 250945 675434 250997
rect 282742 250797 282794 250849
rect 283126 250797 283178 250849
rect 139222 250723 139274 250775
rect 140182 250723 140234 250775
rect 42166 250575 42218 250627
rect 145366 250575 145418 250627
rect 182326 250575 182378 250627
rect 230134 250501 230186 250553
rect 282742 250501 282794 250553
rect 145366 250353 145418 250405
rect 141142 250279 141194 250331
rect 144406 250279 144458 250331
rect 139318 250205 139370 250257
rect 144310 250205 144362 250257
rect 674806 250205 674858 250257
rect 675286 250205 675338 250257
rect 139798 250131 139850 250183
rect 141334 250131 141386 250183
rect 139894 250057 139946 250109
rect 141238 250057 141290 250109
rect 44566 249983 44618 250035
rect 200086 249983 200138 250035
rect 218422 249095 218474 249147
rect 218806 249095 218858 249147
rect 541462 249095 541514 249147
rect 541846 249095 541898 249147
rect 282358 248873 282410 248925
rect 283894 248873 283946 248925
rect 288310 248355 288362 248407
rect 288118 248281 288170 248333
rect 288022 248133 288074 248185
rect 144022 247763 144074 247815
rect 191446 247763 191498 247815
rect 285622 247763 285674 247815
rect 145462 247689 145514 247741
rect 148246 247689 148298 247741
rect 286006 247689 286058 247741
rect 532918 247689 532970 247741
rect 533398 247689 533450 247741
rect 541558 247689 541610 247741
rect 541750 247689 541802 247741
rect 34582 247615 34634 247667
rect 42166 247615 42218 247667
rect 235894 247615 235946 247667
rect 282358 247615 282410 247667
rect 285622 247615 285674 247667
rect 285910 247615 285962 247667
rect 288310 247615 288362 247667
rect 182326 247541 182378 247593
rect 200758 247541 200810 247593
rect 674422 246727 674474 246779
rect 675190 246727 675242 246779
rect 282742 245247 282794 245299
rect 282742 245099 282794 245151
rect 283318 245099 283370 245151
rect 144118 244877 144170 244929
rect 148438 244877 148490 244929
rect 144022 244803 144074 244855
rect 197206 244803 197258 244855
rect 282166 244803 282218 244855
rect 282646 244803 282698 244855
rect 283798 244803 283850 244855
rect 284278 244803 284330 244855
rect 42070 244729 42122 244781
rect 42550 244729 42602 244781
rect 241654 244729 241706 244781
rect 282262 244729 282314 244781
rect 253366 244655 253418 244707
rect 284278 244655 284330 244707
rect 262006 244581 262058 244633
rect 282262 244581 282314 244633
rect 282454 244581 282506 244633
rect 282646 244581 282698 244633
rect 288310 244729 288362 244781
rect 267766 244507 267818 244559
rect 283030 244507 283082 244559
rect 37270 244433 37322 244485
rect 41782 244433 41834 244485
rect 144406 244433 144458 244485
rect 149590 244433 149642 244485
rect 276406 244433 276458 244485
rect 282454 244433 282506 244485
rect 288310 244507 288362 244559
rect 284278 243989 284330 244041
rect 139990 243619 140042 243671
rect 142198 243619 142250 243671
rect 674998 242953 675050 243005
rect 675382 242953 675434 243005
rect 674134 242361 674186 242413
rect 675382 242361 675434 242413
rect 41974 242287 42026 242339
rect 42742 242287 42794 242339
rect 43126 242065 43178 242117
rect 43510 242065 43562 242117
rect 37174 241991 37226 242043
rect 42646 241991 42698 242043
rect 144022 241991 144074 242043
rect 151126 241991 151178 242043
rect 288310 241991 288362 242043
rect 37366 241917 37418 241969
rect 43126 241917 43178 241969
rect 145750 241917 145802 241969
rect 148630 241917 148682 241969
rect 204214 241917 204266 241969
rect 207382 241917 207434 241969
rect 146806 241843 146858 241895
rect 152086 241843 152138 241895
rect 288310 241769 288362 241821
rect 674326 241695 674378 241747
rect 675478 241695 675530 241747
rect 42742 240733 42794 240785
rect 43222 240733 43274 240785
rect 41782 240585 41834 240637
rect 674902 240511 674954 240563
rect 675478 240511 675530 240563
rect 140182 240437 140234 240489
rect 141430 240437 141482 240489
rect 41782 240363 41834 240415
rect 288598 239623 288650 239675
rect 290518 239623 290570 239675
rect 366694 239623 366746 239675
rect 373942 239623 373994 239675
rect 381526 239623 381578 239675
rect 388918 239623 388970 239675
rect 396118 239623 396170 239675
rect 541654 239623 541706 239675
rect 288118 239549 288170 239601
rect 289414 239549 289466 239601
rect 288214 239475 288266 239527
rect 409270 239549 409322 239601
rect 409462 239549 409514 239601
rect 414550 239549 414602 239601
rect 437782 239549 437834 239601
rect 443734 239549 443786 239601
rect 443974 239549 444026 239601
rect 454006 239549 454058 239601
rect 291190 239475 291242 239527
rect 381526 239475 381578 239527
rect 401878 239475 401930 239527
rect 293110 239253 293162 239305
rect 401398 239401 401450 239453
rect 406390 239401 406442 239453
rect 406582 239475 406634 239527
rect 408886 239475 408938 239527
rect 410326 239475 410378 239527
rect 410998 239475 411050 239527
rect 411574 239475 411626 239527
rect 412054 239475 412106 239527
rect 445270 239475 445322 239527
rect 388918 239253 388970 239305
rect 401878 239253 401930 239305
rect 405334 239327 405386 239379
rect 410230 239327 410282 239379
rect 444406 239401 444458 239453
rect 411094 239327 411146 239379
rect 414070 239327 414122 239379
rect 444118 239327 444170 239379
rect 446326 239327 446378 239379
rect 447958 239327 448010 239379
rect 406582 239253 406634 239305
rect 407542 239253 407594 239305
rect 408886 239253 408938 239305
rect 412150 239253 412202 239305
rect 444310 239253 444362 239305
rect 140374 239179 140426 239231
rect 141142 239179 141194 239231
rect 288406 239179 288458 239231
rect 406294 239179 406346 239231
rect 408502 239179 408554 239231
rect 443542 239179 443594 239231
rect 149590 239105 149642 239157
rect 155350 239105 155402 239157
rect 391318 239105 391370 239157
rect 457942 239105 457994 239157
rect 144022 239031 144074 239083
rect 188566 239031 188618 239083
rect 325462 239031 325514 239083
rect 341590 239031 341642 239083
rect 345814 239031 345866 239083
rect 365494 239031 365546 239083
rect 391702 239031 391754 239083
rect 392662 239031 392714 239083
rect 397462 239031 397514 239083
rect 413686 239031 413738 239083
rect 413878 239031 413930 239083
rect 419638 239031 419690 239083
rect 146902 238957 146954 239009
rect 149782 238957 149834 239009
rect 218710 238957 218762 239009
rect 342742 238957 342794 239009
rect 344278 238957 344330 239009
rect 354742 238957 354794 239009
rect 354838 238957 354890 239009
rect 518422 238957 518474 239009
rect 227350 238883 227402 238935
rect 349366 238883 349418 238935
rect 350710 238883 350762 238935
rect 353206 238883 353258 238935
rect 283894 238809 283946 238861
rect 340150 238809 340202 238861
rect 342742 238809 342794 238861
rect 345334 238809 345386 238861
rect 346870 238809 346922 238861
rect 354454 238883 354506 238935
rect 354550 238883 354602 238935
rect 512950 238883 513002 238935
rect 140566 238735 140618 238787
rect 140950 238735 141002 238787
rect 289558 238735 289610 238787
rect 354358 238735 354410 238787
rect 354454 238735 354506 238787
rect 501238 238809 501290 238861
rect 283702 238661 283754 238713
rect 339478 238661 339530 238713
rect 346486 238661 346538 238713
rect 359158 238735 359210 238787
rect 507094 238735 507146 238787
rect 495478 238661 495530 238713
rect 285046 238587 285098 238639
rect 337174 238587 337226 238639
rect 337270 238587 337322 238639
rect 358486 238587 358538 238639
rect 360502 238587 360554 238639
rect 501334 238587 501386 238639
rect 42166 238513 42218 238565
rect 42358 238513 42410 238565
rect 287062 238513 287114 238565
rect 340534 238513 340586 238565
rect 346102 238513 346154 238565
rect 486838 238513 486890 238565
rect 42550 238439 42602 238491
rect 286582 238439 286634 238491
rect 339862 238439 339914 238491
rect 345718 238439 345770 238491
rect 481174 238439 481226 238491
rect 42358 238365 42410 238417
rect 286870 238365 286922 238417
rect 340918 238365 340970 238417
rect 341014 238365 341066 238417
rect 362134 238365 362186 238417
rect 390166 238365 390218 238417
rect 407830 238365 407882 238417
rect 408022 238365 408074 238417
rect 410998 238365 411050 238417
rect 411286 238365 411338 238417
rect 541462 238365 541514 238417
rect 286774 238291 286826 238343
rect 387286 238291 387338 238343
rect 392854 238291 392906 238343
rect 405910 238291 405962 238343
rect 406102 238291 406154 238343
rect 532918 238291 532970 238343
rect 286006 238217 286058 238269
rect 339094 238217 339146 238269
rect 344950 238217 345002 238269
rect 469462 238217 469514 238269
rect 285238 238143 285290 238195
rect 345622 238143 345674 238195
rect 402646 238143 402698 238195
rect 403126 238143 403178 238195
rect 403222 238143 403274 238195
rect 527254 238143 527306 238195
rect 305110 237995 305162 238047
rect 337174 238069 337226 238121
rect 341110 238069 341162 238121
rect 344662 238069 344714 238121
rect 345526 237995 345578 238047
rect 463702 238069 463754 238121
rect 365686 237995 365738 238047
rect 390166 237995 390218 238047
rect 393910 237995 393962 238047
rect 504022 237995 504074 238047
rect 288022 237921 288074 237973
rect 350710 237921 350762 237973
rect 350806 237921 350858 237973
rect 361462 237921 361514 237973
rect 366358 237921 366410 237973
rect 485494 237921 485546 237973
rect 288310 237847 288362 237899
rect 325558 237847 325610 237899
rect 325942 237847 325994 237899
rect 398902 237847 398954 237899
rect 282550 237773 282602 237825
rect 406006 237847 406058 237899
rect 408982 237847 409034 237899
rect 430582 237847 430634 237899
rect 435094 237847 435146 237899
rect 533014 237847 533066 237899
rect 399478 237773 399530 237825
rect 419062 237773 419114 237825
rect 436822 237773 436874 237825
rect 541558 237773 541610 237825
rect 42166 237699 42218 237751
rect 50422 237699 50474 237751
rect 287926 237699 287978 237751
rect 350806 237699 350858 237751
rect 350902 237699 350954 237751
rect 477814 237699 477866 237751
rect 350134 237625 350186 237677
rect 477430 237625 477482 237677
rect 140854 237551 140906 237603
rect 287350 237551 287402 237603
rect 331414 237551 331466 237603
rect 338518 237551 338570 237603
rect 351574 237551 351626 237603
rect 478198 237551 478250 237603
rect 334678 237477 334730 237529
rect 449398 237477 449450 237529
rect 140950 237329 141002 237381
rect 332086 237403 332138 237455
rect 446806 237403 446858 237455
rect 332470 237329 332522 237381
rect 447286 237329 447338 237381
rect 335446 237255 335498 237307
rect 450262 237255 450314 237307
rect 336118 237181 336170 237233
rect 450838 237181 450890 237233
rect 333238 237107 333290 237159
rect 448054 237107 448106 237159
rect 356278 237033 356330 237085
rect 358486 237033 358538 237085
rect 451798 237033 451850 237085
rect 287638 236959 287690 237011
rect 364726 236959 364778 237011
rect 398134 236959 398186 237011
rect 460822 236959 460874 237011
rect 285814 236885 285866 236937
rect 365302 236885 365354 236937
rect 397270 236885 397322 236937
rect 453814 236885 453866 236937
rect 284854 236811 284906 236863
rect 358102 236811 358154 236863
rect 398806 236811 398858 236863
rect 418966 236811 419018 236863
rect 419062 236811 419114 236863
rect 454966 236811 455018 236863
rect 285142 236737 285194 236789
rect 341014 236737 341066 236789
rect 341110 236737 341162 236789
rect 42166 236663 42218 236715
rect 43126 236663 43178 236715
rect 287734 236589 287786 236641
rect 351958 236663 352010 236715
rect 354742 236737 354794 236789
rect 455446 236737 455498 236789
rect 355510 236663 355562 236715
rect 398902 236663 398954 236715
rect 409078 236663 409130 236715
rect 409174 236663 409226 236715
rect 413878 236663 413930 236715
rect 144022 236515 144074 236567
rect 148822 236515 148874 236567
rect 287830 236515 287882 236567
rect 360598 236589 360650 236641
rect 398998 236589 399050 236641
rect 430294 236663 430346 236715
rect 433270 236663 433322 236715
rect 440182 236663 440234 236715
rect 418966 236589 419018 236641
rect 453430 236589 453482 236641
rect 338422 236515 338474 236567
rect 359254 236515 359306 236567
rect 389206 236515 389258 236567
rect 399190 236515 399242 236567
rect 400342 236515 400394 236567
rect 479638 236515 479690 236567
rect 287254 236441 287306 236493
rect 357430 236441 357482 236493
rect 397846 236441 397898 236493
rect 399958 236441 400010 236493
rect 400054 236441 400106 236493
rect 479254 236441 479306 236493
rect 287542 236367 287594 236419
rect 338230 236367 338282 236419
rect 338326 236367 338378 236419
rect 359638 236367 359690 236419
rect 360118 236367 360170 236419
rect 377302 236367 377354 236419
rect 398710 236367 398762 236419
rect 478870 236367 478922 236419
rect 296566 236293 296618 236345
rect 351958 236293 352010 236345
rect 287446 236219 287498 236271
rect 338326 236219 338378 236271
rect 345622 236219 345674 236271
rect 357046 236293 357098 236345
rect 396502 236293 396554 236345
rect 398902 236293 398954 236345
rect 478486 236293 478538 236345
rect 360310 236219 360362 236271
rect 360406 236219 360458 236271
rect 377110 236219 377162 236271
rect 397750 236219 397802 236271
rect 482614 236219 482666 236271
rect 140182 236145 140234 236197
rect 141238 236145 141290 236197
rect 287158 236145 287210 236197
rect 355222 236145 355274 236197
rect 390166 236145 390218 236197
rect 399478 236145 399530 236197
rect 399958 236145 400010 236197
rect 218806 236071 218858 236123
rect 298198 236071 298250 236123
rect 327286 236071 327338 236123
rect 353590 236071 353642 236123
rect 353782 236071 353834 236123
rect 400054 236071 400106 236123
rect 400246 236145 400298 236197
rect 482902 236145 482954 236197
rect 404470 236071 404522 236123
rect 404566 236071 404618 236123
rect 451990 236071 452042 236123
rect 452182 236071 452234 236123
rect 453526 236071 453578 236123
rect 453910 236071 453962 236123
rect 501142 236071 501194 236123
rect 204310 235997 204362 236049
rect 290134 235997 290186 236049
rect 324406 235997 324458 236049
rect 338230 235997 338282 236049
rect 338326 235997 338378 236049
rect 348886 235997 348938 236049
rect 354646 235997 354698 236049
rect 400342 235997 400394 236049
rect 401686 235997 401738 236049
rect 403798 235997 403850 236049
rect 403894 235997 403946 236049
rect 414838 235997 414890 236049
rect 414934 235997 414986 236049
rect 420310 235997 420362 236049
rect 420790 235997 420842 236049
rect 430678 235997 430730 236049
rect 434422 235997 434474 236049
rect 443638 235997 443690 236049
rect 444694 235997 444746 236049
rect 494998 235997 495050 236049
rect 209974 235923 210026 235975
rect 294166 235923 294218 235975
rect 325078 235923 325130 235975
rect 374998 235923 375050 235975
rect 375094 235923 375146 235975
rect 391510 235923 391562 235975
rect 398422 235923 398474 235975
rect 400246 235923 400298 235975
rect 400534 235923 400586 235975
rect 408790 235923 408842 235975
rect 408886 235923 408938 235975
rect 413014 235923 413066 235975
rect 413110 235923 413162 235975
rect 418486 235923 418538 235975
rect 418582 235923 418634 235975
rect 420406 235923 420458 235975
rect 425110 235923 425162 235975
rect 446326 235923 446378 235975
rect 446902 235923 446954 235975
rect 497878 235923 497930 235975
rect 285430 235849 285482 235901
rect 374326 235849 374378 235901
rect 374422 235849 374474 235901
rect 377206 235849 377258 235901
rect 395734 235849 395786 235901
rect 405430 235849 405482 235901
rect 285526 235775 285578 235827
rect 378838 235775 378890 235827
rect 389110 235775 389162 235827
rect 140086 235701 140138 235753
rect 141526 235701 141578 235753
rect 224566 235701 224618 235753
rect 302230 235701 302282 235753
rect 334294 235701 334346 235753
rect 284374 235627 284426 235679
rect 375094 235627 375146 235679
rect 375286 235627 375338 235679
rect 398806 235627 398858 235679
rect 338230 235553 338282 235605
rect 338710 235553 338762 235605
rect 338998 235553 339050 235605
rect 346774 235553 346826 235605
rect 357046 235553 357098 235605
rect 390166 235553 390218 235605
rect 399286 235775 399338 235827
rect 409462 235849 409514 235901
rect 411766 235849 411818 235901
rect 420502 235849 420554 235901
rect 420598 235849 420650 235901
rect 441526 235849 441578 235901
rect 443254 235849 443306 235901
rect 493750 235849 493802 235901
rect 406102 235775 406154 235827
rect 435574 235775 435626 235827
rect 441814 235775 441866 235827
rect 493558 235775 493610 235827
rect 399190 235701 399242 235753
rect 420598 235701 420650 235753
rect 420790 235701 420842 235753
rect 436438 235701 436490 235753
rect 440278 235701 440330 235753
rect 494806 235701 494858 235753
rect 412630 235627 412682 235679
rect 412726 235627 412778 235679
rect 414646 235627 414698 235679
rect 414838 235627 414890 235679
rect 420118 235627 420170 235679
rect 420886 235627 420938 235679
rect 437782 235627 437834 235679
rect 438838 235627 438890 235679
rect 494422 235627 494474 235679
rect 399190 235553 399242 235605
rect 399478 235553 399530 235605
rect 417622 235553 417674 235605
rect 424438 235553 424490 235605
rect 431350 235553 431402 235605
rect 439126 235553 439178 235605
rect 449782 235553 449834 235605
rect 449878 235553 449930 235605
rect 506902 235553 506954 235605
rect 312982 235479 313034 235531
rect 338326 235479 338378 235531
rect 353590 235479 353642 235531
rect 360118 235479 360170 235531
rect 42166 235405 42218 235457
rect 43030 235405 43082 235457
rect 311542 235405 311594 235457
rect 338614 235405 338666 235457
rect 338806 235405 338858 235457
rect 375286 235479 375338 235531
rect 377014 235405 377066 235457
rect 491734 235479 491786 235531
rect 382870 235405 382922 235457
rect 497686 235405 497738 235457
rect 309334 235331 309386 235383
rect 352150 235331 352202 235383
rect 356374 235331 356426 235383
rect 360118 235331 360170 235383
rect 360406 235331 360458 235383
rect 360694 235331 360746 235383
rect 328438 235257 328490 235309
rect 338134 235257 338186 235309
rect 338518 235257 338570 235309
rect 354838 235257 354890 235309
rect 355702 235257 355754 235309
rect 379510 235331 379562 235383
rect 379990 235331 380042 235383
rect 494710 235331 494762 235383
rect 317014 235183 317066 235235
rect 140182 235109 140234 235161
rect 141910 235109 141962 235161
rect 314038 235109 314090 235161
rect 338326 235109 338378 235161
rect 338422 235109 338474 235161
rect 344470 235109 344522 235161
rect 354934 235183 354986 235235
rect 379894 235257 379946 235309
rect 382198 235257 382250 235309
rect 496918 235257 496970 235309
rect 360694 235109 360746 235161
rect 360790 235109 360842 235161
rect 376822 235183 376874 235235
rect 379222 235183 379274 235235
rect 494038 235183 494090 235235
rect 376246 235109 376298 235161
rect 491062 235109 491114 235161
rect 311158 235035 311210 235087
rect 355030 235035 355082 235087
rect 357910 235035 357962 235087
rect 372790 235035 372842 235087
rect 372982 235035 373034 235087
rect 488854 235035 488906 235087
rect 318838 234961 318890 235013
rect 356854 234961 356906 235013
rect 357142 234961 357194 235013
rect 375382 234961 375434 235013
rect 321046 234887 321098 234939
rect 357718 234887 357770 234939
rect 359350 234887 359402 234939
rect 377686 234961 377738 235013
rect 378454 234961 378506 235013
rect 493270 234961 493322 235013
rect 375574 234887 375626 234939
rect 310006 234813 310058 234865
rect 338230 234813 338282 234865
rect 338326 234813 338378 234865
rect 359830 234813 359882 234865
rect 361174 234813 361226 234865
rect 378742 234813 378794 234865
rect 381430 234887 381482 234939
rect 496150 234887 496202 234939
rect 490294 234813 490346 234865
rect 318166 234739 318218 234791
rect 356086 234739 356138 234791
rect 358582 234739 358634 234791
rect 378070 234739 378122 234791
rect 380662 234739 380714 234791
rect 495478 234739 495530 234791
rect 42358 234665 42410 234717
rect 43510 234665 43562 234717
rect 317398 234665 317450 234717
rect 355894 234665 355946 234717
rect 377782 234665 377834 234717
rect 492502 234665 492554 234717
rect 311830 234443 311882 234495
rect 329878 234591 329930 234643
rect 344278 234517 344330 234569
rect 344470 234591 344522 234643
rect 378646 234591 378698 234643
rect 378838 234591 378890 234643
rect 390550 234591 390602 234643
rect 395734 234591 395786 234643
rect 408694 234591 408746 234643
rect 414742 234591 414794 234643
rect 415990 234591 416042 234643
rect 417718 234591 417770 234643
rect 419926 234591 419978 234643
rect 420022 234591 420074 234643
rect 443542 234591 443594 234643
rect 443638 234591 443690 234643
rect 446422 234591 446474 234643
rect 448438 234591 448490 234643
rect 498070 234591 498122 234643
rect 375958 234517 376010 234569
rect 396502 234517 396554 234569
rect 405046 234517 405098 234569
rect 408310 234517 408362 234569
rect 439126 234517 439178 234569
rect 442486 234517 442538 234569
rect 447478 234517 447530 234569
rect 451318 234517 451370 234569
rect 499702 234517 499754 234569
rect 329494 234443 329546 234495
rect 338998 234443 339050 234495
rect 342742 234443 342794 234495
rect 398134 234443 398186 234495
rect 399190 234443 399242 234495
rect 408790 234443 408842 234495
rect 408982 234443 409034 234495
rect 417430 234443 417482 234495
rect 417814 234443 417866 234495
rect 425878 234443 425930 234495
rect 426166 234443 426218 234495
rect 446134 234443 446186 234495
rect 446230 234443 446282 234495
rect 493942 234443 493994 234495
rect 312214 234369 312266 234421
rect 354742 234369 354794 234421
rect 310774 234295 310826 234347
rect 351670 234295 351722 234347
rect 353494 234295 353546 234347
rect 360982 234369 361034 234421
rect 361942 234369 361994 234421
rect 393430 234369 393482 234421
rect 393526 234369 393578 234421
rect 400246 234369 400298 234421
rect 400342 234369 400394 234421
rect 408022 234369 408074 234421
rect 408118 234369 408170 234421
rect 418870 234369 418922 234421
rect 355894 234295 355946 234347
rect 363478 234295 363530 234347
rect 365974 234295 366026 234347
rect 367990 234295 368042 234347
rect 368662 234295 368714 234347
rect 376246 234295 376298 234347
rect 388054 234295 388106 234347
rect 408406 234295 408458 234347
rect 424246 234369 424298 234421
rect 431926 234369 431978 234421
rect 452182 234369 452234 234421
rect 452854 234369 452906 234421
rect 499606 234369 499658 234421
rect 320374 234221 320426 234273
rect 359926 234221 359978 234273
rect 361558 234221 361610 234273
rect 376534 234221 376586 234273
rect 377206 234221 377258 234273
rect 397366 234221 397418 234273
rect 42454 234147 42506 234199
rect 323638 234147 323690 234199
rect 338518 234147 338570 234199
rect 338614 234147 338666 234199
rect 355126 234147 355178 234199
rect 362326 234147 362378 234199
rect 368662 234147 368714 234199
rect 374998 234147 375050 234199
rect 394582 234147 394634 234199
rect 397270 234147 397322 234199
rect 399286 234221 399338 234273
rect 399478 234221 399530 234273
rect 397558 234147 397610 234199
rect 404662 234147 404714 234199
rect 313750 234073 313802 234125
rect 327190 234073 327242 234125
rect 328726 234073 328778 234125
rect 346678 234073 346730 234125
rect 346774 234073 346826 234125
rect 352630 234073 352682 234125
rect 352726 234073 352778 234125
rect 362806 234073 362858 234125
rect 375958 234073 376010 234125
rect 395158 234073 395210 234125
rect 396886 234073 396938 234125
rect 405142 234073 405194 234125
rect 407062 234221 407114 234273
rect 410038 234221 410090 234273
rect 416758 234221 416810 234273
rect 418486 234221 418538 234273
rect 428086 234295 428138 234347
rect 431446 234295 431498 234347
rect 475606 234295 475658 234347
rect 422998 234221 423050 234273
rect 450550 234221 450602 234273
rect 450646 234221 450698 234273
rect 451894 234221 451946 234273
rect 405910 234147 405962 234199
rect 415318 234147 415370 234199
rect 415510 234147 415562 234199
rect 425398 234147 425450 234199
rect 425974 234147 426026 234199
rect 470038 234147 470090 234199
rect 42070 233999 42122 234051
rect 42454 233999 42506 234051
rect 43126 233999 43178 234051
rect 314422 233999 314474 234051
rect 327094 233999 327146 234051
rect 338326 233999 338378 234051
rect 351478 233999 351530 234051
rect 352342 233999 352394 234051
rect 398902 233999 398954 234051
rect 400150 233999 400202 234051
rect 408598 233999 408650 234051
rect 408886 234073 408938 234125
rect 410806 234073 410858 234125
rect 410902 234073 410954 234125
rect 426262 234073 426314 234125
rect 427414 234073 427466 234125
rect 471574 234073 471626 234125
rect 410134 233999 410186 234051
rect 410422 233999 410474 234051
rect 415222 233999 415274 234051
rect 416374 233999 416426 234051
rect 428470 233999 428522 234051
rect 428854 233999 428906 234051
rect 470614 233999 470666 234051
rect 322198 233925 322250 233977
rect 338422 233925 338474 233977
rect 338710 233925 338762 233977
rect 349174 233925 349226 233977
rect 356086 233925 356138 233977
rect 363574 233925 363626 233977
rect 319606 233851 319658 233903
rect 354454 233851 354506 233903
rect 364534 233851 364586 233903
rect 375094 233925 375146 233977
rect 378646 233925 378698 233977
rect 395254 233925 395306 233977
rect 400630 233925 400682 233977
rect 407926 233925 407978 233977
rect 411766 233925 411818 233977
rect 429910 233925 429962 233977
rect 430774 233925 430826 233977
rect 474838 233925 474890 233977
rect 374326 233851 374378 233903
rect 388342 233851 388394 233903
rect 394774 233851 394826 233903
rect 400534 233851 400586 233903
rect 400918 233851 400970 233903
rect 407158 233851 407210 233903
rect 407254 233851 407306 233903
rect 410038 233851 410090 233903
rect 319990 233777 320042 233829
rect 354262 233777 354314 233829
rect 357718 233777 357770 233829
rect 320662 233703 320714 233755
rect 308950 233629 309002 233681
rect 326902 233629 326954 233681
rect 321430 233555 321482 233607
rect 327094 233703 327146 233755
rect 327190 233629 327242 233681
rect 328726 233629 328778 233681
rect 328822 233629 328874 233681
rect 330454 233629 330506 233681
rect 338422 233703 338474 233755
rect 359542 233703 359594 233755
rect 360982 233777 361034 233829
rect 365110 233777 365162 233829
rect 365206 233777 365258 233829
rect 368662 233777 368714 233829
rect 366646 233703 366698 233755
rect 387670 233777 387722 233829
rect 393430 233777 393482 233829
rect 398902 233777 398954 233829
rect 399862 233777 399914 233829
rect 404566 233777 404618 233829
rect 404662 233777 404714 233829
rect 413782 233851 413834 233903
rect 413878 233851 413930 233903
rect 425110 233851 425162 233903
rect 425206 233851 425258 233903
rect 469366 233851 469418 233903
rect 410518 233777 410570 233829
rect 428374 233777 428426 233829
rect 428470 233777 428522 233829
rect 456118 233777 456170 233829
rect 348502 233629 348554 233681
rect 352630 233629 352682 233681
rect 367126 233629 367178 233681
rect 371158 233629 371210 233681
rect 371926 233629 371978 233681
rect 372310 233629 372362 233681
rect 376918 233703 376970 233755
rect 386902 233703 386954 233755
rect 396118 233703 396170 233755
rect 401878 233703 401930 233755
rect 401974 233703 402026 233755
rect 404950 233703 405002 233755
rect 405046 233703 405098 233755
rect 414742 233703 414794 233755
rect 392470 233629 392522 233681
rect 401206 233629 401258 233681
rect 401302 233629 401354 233681
rect 404086 233629 404138 233681
rect 405238 233629 405290 233681
rect 415510 233629 415562 233681
rect 415606 233629 415658 233681
rect 417526 233629 417578 233681
rect 308566 233481 308618 233533
rect 326806 233481 326858 233533
rect 351382 233555 351434 233607
rect 353110 233555 353162 233607
rect 398710 233555 398762 233607
rect 401686 233555 401738 233607
rect 405718 233555 405770 233607
rect 411766 233555 411818 233607
rect 429430 233703 429482 233755
rect 437398 233703 437450 233755
rect 475126 233703 475178 233755
rect 419926 233629 419978 233681
rect 426166 233629 426218 233681
rect 426262 233629 426314 233681
rect 428278 233629 428330 233681
rect 436630 233629 436682 233681
rect 466582 233629 466634 233681
rect 427798 233555 427850 233607
rect 428470 233555 428522 233607
rect 435190 233555 435242 233607
rect 437686 233555 437738 233607
rect 438070 233555 438122 233607
rect 440566 233555 440618 233607
rect 443542 233555 443594 233607
rect 446326 233555 446378 233607
rect 446518 233555 446570 233607
rect 446902 233555 446954 233607
rect 450550 233555 450602 233607
rect 467158 233555 467210 233607
rect 338326 233481 338378 233533
rect 338518 233481 338570 233533
rect 362710 233481 362762 233533
rect 362806 233481 362858 233533
rect 367606 233481 367658 233533
rect 368662 233481 368714 233533
rect 374710 233481 374762 233533
rect 378742 233481 378794 233533
rect 398422 233481 398474 233533
rect 402070 233481 402122 233533
rect 402934 233481 402986 233533
rect 322870 233407 322922 233459
rect 348598 233407 348650 233459
rect 356854 233407 356906 233459
rect 365110 233407 365162 233459
rect 365206 233407 365258 233459
rect 366454 233407 366506 233459
rect 144022 233333 144074 233385
rect 149206 233333 149258 233385
rect 286198 233333 286250 233385
rect 368566 233333 368618 233385
rect 368662 233333 368714 233385
rect 376918 233407 376970 233459
rect 377110 233407 377162 233459
rect 397750 233407 397802 233459
rect 397078 233333 397130 233385
rect 410422 233481 410474 233533
rect 413782 233481 413834 233533
rect 432502 233481 432554 233533
rect 436246 233481 436298 233533
rect 453622 233481 453674 233533
rect 403510 233407 403562 233459
rect 481846 233407 481898 233459
rect 404470 233333 404522 233385
rect 482230 233333 482282 233385
rect 142486 233259 142538 233311
rect 144118 233259 144170 233311
rect 168406 233259 168458 233311
rect 283126 233259 283178 233311
rect 372310 233259 372362 233311
rect 402646 233259 402698 233311
rect 402934 233259 402986 233311
rect 403030 233259 403082 233311
rect 403222 233259 403274 233311
rect 147190 233185 147242 233237
rect 283510 233185 283562 233237
rect 388726 233185 388778 233237
rect 399766 233185 399818 233237
rect 409366 233259 409418 233311
rect 409462 233259 409514 233311
rect 411862 233259 411914 233311
rect 411958 233259 412010 233311
rect 415414 233259 415466 233311
rect 415510 233259 415562 233311
rect 443542 233259 443594 233311
rect 444118 233259 444170 233311
rect 481462 233259 481514 233311
rect 283222 233111 283274 233163
rect 386518 233111 386570 233163
rect 402358 233111 402410 233163
rect 406678 233111 406730 233163
rect 407542 233111 407594 233163
rect 410230 233111 410282 233163
rect 421654 233111 421706 233163
rect 424150 233111 424202 233163
rect 440278 233111 440330 233163
rect 456406 233185 456458 233237
rect 456118 233111 456170 233163
rect 463414 233111 463466 233163
rect 286390 233037 286442 233089
rect 386134 233037 386186 233089
rect 401014 233037 401066 233089
rect 407062 233037 407114 233089
rect 407158 233037 407210 233089
rect 413974 233037 414026 233089
rect 414166 233037 414218 233089
rect 349078 232963 349130 233015
rect 414550 232963 414602 233015
rect 415030 232963 415082 233015
rect 417910 232963 417962 233015
rect 418966 233037 419018 233089
rect 443542 233037 443594 233089
rect 462358 233037 462410 233089
rect 470614 233037 470666 233089
rect 473014 233037 473066 233089
rect 443830 232963 443882 233015
rect 454582 232963 454634 233015
rect 336502 232889 336554 232941
rect 398710 232889 398762 232941
rect 398806 232889 398858 232941
rect 418966 232889 419018 232941
rect 419158 232889 419210 232941
rect 424534 232889 424586 232941
rect 424822 232889 424874 232941
rect 468982 232889 469034 232941
rect 348694 232815 348746 232867
rect 414646 232815 414698 232867
rect 414742 232815 414794 232867
rect 443638 232815 443690 232867
rect 443734 232815 443786 232867
rect 443830 232815 443882 232867
rect 455350 232815 455402 232867
rect 283414 232741 283466 232793
rect 363382 232741 363434 232793
rect 364822 232741 364874 232793
rect 374326 232741 374378 232793
rect 398710 232741 398762 232793
rect 413590 232741 413642 232793
rect 321814 232667 321866 232719
rect 409654 232667 409706 232719
rect 409750 232667 409802 232719
rect 413974 232667 414026 232719
rect 141142 232593 141194 232645
rect 141718 232593 141770 232645
rect 326998 232593 327050 232645
rect 399958 232593 400010 232645
rect 400054 232593 400106 232645
rect 443542 232741 443594 232793
rect 461590 232741 461642 232793
rect 414262 232667 414314 232719
rect 415030 232667 415082 232719
rect 415414 232667 415466 232719
rect 417142 232593 417194 232645
rect 424534 232667 424586 232719
rect 443638 232667 443690 232719
rect 461206 232667 461258 232719
rect 326230 232519 326282 232571
rect 417814 232519 417866 232571
rect 417910 232519 417962 232571
rect 421174 232519 421226 232571
rect 327670 232445 327722 232497
rect 391126 232445 391178 232497
rect 341590 232371 341642 232423
rect 418006 232445 418058 232497
rect 418294 232445 418346 232497
rect 423478 232519 423530 232571
rect 443830 232519 443882 232571
rect 453718 232519 453770 232571
rect 467350 232519 467402 232571
rect 391414 232371 391466 232423
rect 418390 232371 418442 232423
rect 463798 232445 463850 232497
rect 423478 232371 423530 232423
rect 423766 232371 423818 232423
rect 443542 232371 443594 232423
rect 444406 232371 444458 232423
rect 453334 232371 453386 232423
rect 453430 232371 453482 232423
rect 467830 232371 467882 232423
rect 337654 232297 337706 232349
rect 428758 232297 428810 232349
rect 429238 232297 429290 232349
rect 473398 232297 473450 232349
rect 335830 232223 335882 232275
rect 426262 232223 426314 232275
rect 426646 232223 426698 232275
rect 470806 232223 470858 232275
rect 324790 232149 324842 232201
rect 391222 232149 391274 232201
rect 324022 232075 324074 232127
rect 417238 232149 417290 232201
rect 420310 232149 420362 232201
rect 462742 232149 462794 232201
rect 398806 232075 398858 232127
rect 419638 232075 419690 232127
rect 421174 232075 421226 232127
rect 421846 232075 421898 232127
rect 422614 232075 422666 232127
rect 466774 232075 466826 232127
rect 323254 232001 323306 232053
rect 419254 232001 419306 232053
rect 420406 232001 420458 232053
rect 464566 232001 464618 232053
rect 475126 232001 475178 232053
rect 505750 232001 505802 232053
rect 335062 231927 335114 231979
rect 431830 231927 431882 231979
rect 432214 231927 432266 231979
rect 476278 231927 476330 231979
rect 322486 231853 322538 231905
rect 398806 231853 398858 231905
rect 399958 231853 400010 231905
rect 408886 231853 408938 231905
rect 411190 231853 411242 231905
rect 419158 231853 419210 231905
rect 419350 231853 419402 231905
rect 464950 231853 465002 231905
rect 466582 231853 466634 231905
rect 504982 231853 505034 231905
rect 333622 231779 333674 231831
rect 436054 231779 436106 231831
rect 437686 231779 437738 231831
rect 503542 231779 503594 231831
rect 285910 231705 285962 231757
rect 363670 231705 363722 231757
rect 397942 231705 397994 231757
rect 403894 231705 403946 231757
rect 403990 231705 404042 231757
rect 405238 231705 405290 231757
rect 406198 231705 406250 231757
rect 286102 231631 286154 231683
rect 361174 231631 361226 231683
rect 394678 231631 394730 231683
rect 336886 231557 336938 231609
rect 404278 231557 404330 231609
rect 406774 231631 406826 231683
rect 406966 231557 407018 231609
rect 410134 231631 410186 231683
rect 418102 231631 418154 231683
rect 419062 231705 419114 231757
rect 454198 231705 454250 231757
rect 458326 231631 458378 231683
rect 420502 231557 420554 231609
rect 422038 231557 422090 231609
rect 428566 231557 428618 231609
rect 430678 231557 430730 231609
rect 439510 231557 439562 231609
rect 439606 231557 439658 231609
rect 458614 231557 458666 231609
rect 286678 231483 286730 231535
rect 362614 231483 362666 231535
rect 363766 231483 363818 231535
rect 375478 231483 375530 231535
rect 386518 231483 386570 231535
rect 411766 231483 411818 231535
rect 413494 231483 413546 231535
rect 421174 231483 421226 231535
rect 421654 231483 421706 231535
rect 427606 231483 427658 231535
rect 284566 231409 284618 231461
rect 353398 231409 353450 231461
rect 362998 231409 363050 231461
rect 375862 231409 375914 231461
rect 391414 231409 391466 231461
rect 403606 231409 403658 231461
rect 403702 231409 403754 231461
rect 423382 231409 423434 231461
rect 426358 231409 426410 231461
rect 460150 231483 460202 231535
rect 431350 231409 431402 231461
rect 468598 231409 468650 231461
rect 351286 231335 351338 231387
rect 372694 231335 372746 231387
rect 391606 231335 391658 231387
rect 413782 231335 413834 231387
rect 413974 231335 414026 231387
rect 338038 231261 338090 231313
rect 391222 231261 391274 231313
rect 349750 231187 349802 231239
rect 373750 231187 373802 231239
rect 384790 231187 384842 231239
rect 414454 231261 414506 231313
rect 417622 231261 417674 231313
rect 420214 231261 420266 231313
rect 282646 231113 282698 231165
rect 362998 231113 363050 231165
rect 391126 231113 391178 231165
rect 417046 231187 417098 231239
rect 417718 231187 417770 231239
rect 422038 231261 422090 231313
rect 422230 231335 422282 231387
rect 426454 231335 426506 231387
rect 428182 231335 428234 231387
rect 472246 231335 472298 231387
rect 426358 231261 426410 231313
rect 426646 231261 426698 231313
rect 470422 231261 470474 231313
rect 420598 231187 420650 231239
rect 439414 231187 439466 231239
rect 439510 231187 439562 231239
rect 465622 231187 465674 231239
rect 393046 231113 393098 231165
rect 431926 231113 431978 231165
rect 432022 231113 432074 231165
rect 439222 231113 439274 231165
rect 286966 231039 287018 231091
rect 364054 231039 364106 231091
rect 390934 231039 390986 231091
rect 403702 231039 403754 231091
rect 403894 231039 403946 231091
rect 419062 231039 419114 231091
rect 421558 231039 421610 231091
rect 345622 230965 345674 231017
rect 355990 230965 356042 231017
rect 356758 230965 356810 231017
rect 427318 230965 427370 231017
rect 353206 230891 353258 230943
rect 365494 230891 365546 230943
rect 389878 230891 389930 230943
rect 345910 230817 345962 230869
rect 364438 230817 364490 230869
rect 392086 230817 392138 230869
rect 403702 230817 403754 230869
rect 409174 230891 409226 230943
rect 427798 230891 427850 230943
rect 427990 231039 428042 231091
rect 428950 231039 429002 231091
rect 429622 231039 429674 231091
rect 473782 231113 473834 231165
rect 428566 230965 428618 231017
rect 439510 230965 439562 231017
rect 466006 231039 466058 231091
rect 440278 230965 440330 231017
rect 468214 230965 468266 231017
rect 439702 230891 439754 230943
rect 474070 230891 474122 230943
rect 426070 230817 426122 230869
rect 430006 230817 430058 230869
rect 431926 230817 431978 230869
rect 432598 230817 432650 230869
rect 476662 230817 476714 230869
rect 389494 230743 389546 230795
rect 403606 230743 403658 230795
rect 387670 230669 387722 230721
rect 403318 230669 403370 230721
rect 409078 230743 409130 230795
rect 155350 230595 155402 230647
rect 156886 230595 156938 230647
rect 391702 230595 391754 230647
rect 403894 230669 403946 230721
rect 426166 230743 426218 230795
rect 426454 230743 426506 230795
rect 466390 230743 466442 230795
rect 409750 230669 409802 230721
rect 414070 230669 414122 230721
rect 415318 230669 415370 230721
rect 419350 230669 419402 230721
rect 427030 230669 427082 230721
rect 471190 230669 471242 230721
rect 403606 230595 403658 230647
rect 423958 230595 424010 230647
rect 383638 230521 383690 230573
rect 425782 230521 425834 230573
rect 456118 230595 456170 230647
rect 144022 230447 144074 230499
rect 194326 230447 194378 230499
rect 360310 230447 360362 230499
rect 379126 230447 379178 230499
rect 140278 230373 140330 230425
rect 141046 230373 141098 230425
rect 147190 230373 147242 230425
rect 207862 230373 207914 230425
rect 285718 230373 285770 230425
rect 369526 230373 369578 230425
rect 371062 230373 371114 230425
rect 372598 230373 372650 230425
rect 395350 230373 395402 230425
rect 402742 230373 402794 230425
rect 403510 230373 403562 230425
rect 403702 230447 403754 230499
rect 409174 230447 409226 230499
rect 409366 230447 409418 230499
rect 417430 230447 417482 230499
rect 417526 230447 417578 230499
rect 427606 230521 427658 230573
rect 457942 230521 457994 230573
rect 430582 230447 430634 230499
rect 440758 230447 440810 230499
rect 410134 230373 410186 230425
rect 411862 230373 411914 230425
rect 428086 230373 428138 230425
rect 428470 230373 428522 230425
rect 439222 230373 439274 230425
rect 439510 230373 439562 230425
rect 442774 230373 442826 230425
rect 149782 230299 149834 230351
rect 207766 230299 207818 230351
rect 283990 230299 284042 230351
rect 357814 230299 357866 230351
rect 152086 230225 152138 230277
rect 208150 230225 208202 230277
rect 283318 230225 283370 230277
rect 367414 230299 367466 230351
rect 367606 230299 367658 230351
rect 370294 230299 370346 230351
rect 370390 230299 370442 230351
rect 372214 230299 372266 230351
rect 393526 230299 393578 230351
rect 402262 230299 402314 230351
rect 402358 230299 402410 230351
rect 404182 230299 404234 230351
rect 404278 230299 404330 230351
rect 446326 230447 446378 230499
rect 465238 230447 465290 230499
rect 443254 230373 443306 230425
rect 495190 230373 495242 230425
rect 495286 230373 495338 230425
rect 500950 230373 501002 230425
rect 451702 230299 451754 230351
rect 451894 230299 451946 230351
rect 463126 230299 463178 230351
rect 166966 230151 167018 230203
rect 212470 230151 212522 230203
rect 285334 230151 285386 230203
rect 368854 230225 368906 230277
rect 370774 230225 370826 230277
rect 373270 230225 373322 230277
rect 373654 230225 373706 230277
rect 382870 230225 382922 230277
rect 387286 230225 387338 230277
rect 398518 230225 398570 230277
rect 399094 230225 399146 230277
rect 404950 230225 405002 230277
rect 367510 230151 367562 230203
rect 369430 230151 369482 230203
rect 369622 230151 369674 230203
rect 372502 230151 372554 230203
rect 373750 230151 373802 230203
rect 382486 230151 382538 230203
rect 398710 230151 398762 230203
rect 400246 230151 400298 230203
rect 400438 230151 400490 230203
rect 404182 230151 404234 230203
rect 404374 230151 404426 230203
rect 413494 230225 413546 230277
rect 413590 230225 413642 230277
rect 427990 230225 428042 230277
rect 428758 230225 428810 230277
rect 429334 230225 429386 230277
rect 431062 230225 431114 230277
rect 436918 230225 436970 230277
rect 437014 230225 437066 230277
rect 443062 230225 443114 230277
rect 405238 230151 405290 230203
rect 419158 230151 419210 230203
rect 425590 230151 425642 230203
rect 439126 230151 439178 230203
rect 161206 230077 161258 230129
rect 212086 230077 212138 230129
rect 352342 230077 352394 230129
rect 152566 230003 152618 230055
rect 211702 230003 211754 230055
rect 351958 230003 352010 230055
rect 146518 229929 146570 229981
rect 211030 229929 211082 229981
rect 350134 229929 350186 229981
rect 140758 229855 140810 229907
rect 209494 229855 209546 229907
rect 349750 229855 349802 229907
rect 140662 229781 140714 229833
rect 209878 229781 209930 229833
rect 348982 229781 349034 229833
rect 140950 229707 141002 229759
rect 208822 229707 208874 229759
rect 348694 229707 348746 229759
rect 140470 229633 140522 229685
rect 209110 229633 209162 229685
rect 348310 229633 348362 229685
rect 432598 229633 432650 229685
rect 140374 229485 140426 229537
rect 210646 229559 210698 229611
rect 347926 229559 347978 229611
rect 368086 229559 368138 229611
rect 368182 229559 368234 229611
rect 373270 229559 373322 229611
rect 373366 229559 373418 229611
rect 432406 229559 432458 229611
rect 141142 229485 141194 229537
rect 210262 229485 210314 229537
rect 350518 229485 350570 229537
rect 354070 229485 354122 229537
rect 354166 229485 354218 229537
rect 358390 229485 358442 229537
rect 358486 229485 358538 229537
rect 432310 229485 432362 229537
rect 434806 230077 434858 230129
rect 440182 230151 440234 230203
rect 501718 230225 501770 230277
rect 483862 230151 483914 230203
rect 495190 230151 495242 230203
rect 505366 230151 505418 230203
rect 454678 230077 454730 230129
rect 501334 230077 501386 230129
rect 439798 230003 439850 230055
rect 507574 230003 507626 230055
rect 438838 229929 438890 229981
rect 439030 229929 439082 229981
rect 447862 229929 447914 229981
rect 452086 229929 452138 229981
rect 480406 229929 480458 229981
rect 494422 229929 494474 229981
rect 507190 229929 507242 229981
rect 439894 229855 439946 229907
rect 439990 229855 440042 229907
rect 445942 229855 445994 229907
rect 446422 229855 446474 229907
rect 502774 229855 502826 229907
rect 443638 229781 443690 229833
rect 436054 229707 436106 229759
rect 445558 229781 445610 229833
rect 510550 229781 510602 229833
rect 448342 229707 448394 229759
rect 453622 229707 453674 229759
rect 504694 229707 504746 229759
rect 444502 229633 444554 229685
rect 447478 229633 447530 229685
rect 459286 229633 459338 229685
rect 501142 229633 501194 229685
rect 514582 229633 514634 229685
rect 445846 229559 445898 229611
rect 445942 229559 445994 229611
rect 447670 229559 447722 229611
rect 511606 229559 511658 229611
rect 633814 229559 633866 229611
rect 649846 229559 649898 229611
rect 446902 229485 446954 229537
rect 447478 229485 447530 229537
rect 449110 229485 449162 229537
rect 512374 229485 512426 229537
rect 633142 229485 633194 229537
rect 649558 229485 649610 229537
rect 663958 229485 664010 229537
rect 674422 229485 674474 229537
rect 139990 229411 140042 229463
rect 140566 229411 140618 229463
rect 215062 229411 215114 229463
rect 282838 229411 282890 229463
rect 370198 229411 370250 229463
rect 370390 229411 370442 229463
rect 374038 229411 374090 229463
rect 375190 229411 375242 229463
rect 382774 229411 382826 229463
rect 398326 229411 398378 229463
rect 405334 229411 405386 229463
rect 406390 229411 406442 229463
rect 413014 229411 413066 229463
rect 413110 229411 413162 229463
rect 427606 229411 427658 229463
rect 428182 229411 428234 229463
rect 433078 229411 433130 229463
rect 433654 229411 433706 229463
rect 479446 229411 479498 229463
rect 494806 229411 494858 229463
rect 507958 229411 508010 229463
rect 632758 229411 632810 229463
rect 649462 229411 649514 229463
rect 211318 229337 211370 229389
rect 347158 229337 347210 229389
rect 449494 229337 449546 229389
rect 451990 229337 452042 229389
rect 513814 229337 513866 229389
rect 632374 229337 632426 229389
rect 650422 229337 650474 229389
rect 141238 229263 141290 229315
rect 213910 229263 213962 229315
rect 347542 229263 347594 229315
rect 358486 229263 358538 229315
rect 358582 229263 358634 229315
rect 367894 229263 367946 229315
rect 139990 229189 140042 229241
rect 141430 229189 141482 229241
rect 214678 229189 214730 229241
rect 284182 229189 284234 229241
rect 356278 229189 356330 229241
rect 215446 229115 215498 229167
rect 282934 229115 282986 229167
rect 366646 229189 366698 229241
rect 144310 229041 144362 229093
rect 215734 229041 215786 229093
rect 282262 229041 282314 229093
rect 358198 229115 358250 229167
rect 358774 229115 358826 229167
rect 368182 229115 368234 229167
rect 417622 229263 417674 229315
rect 456118 229263 456170 229315
rect 463030 229263 463082 229315
rect 463126 229263 463178 229315
rect 513142 229263 513194 229315
rect 631990 229263 632042 229315
rect 650230 229263 650282 229315
rect 369430 229189 369482 229241
rect 373654 229189 373706 229241
rect 376726 229189 376778 229241
rect 370294 229115 370346 229167
rect 381046 229115 381098 229167
rect 148726 228967 148778 229019
rect 288694 228967 288746 229019
rect 318838 228967 318890 229019
rect 346486 228967 346538 229019
rect 372694 229041 372746 229093
rect 381718 229041 381770 229093
rect 382774 229189 382826 229241
rect 382870 229115 382922 229167
rect 477526 229115 477578 229167
rect 479446 229189 479498 229241
rect 502102 229189 502154 229241
rect 631606 229189 631658 229241
rect 650134 229189 650186 229241
rect 489910 229115 489962 229167
rect 493558 229115 493610 229167
rect 508726 229115 508778 229167
rect 631318 229115 631370 229167
rect 649942 229115 649994 229167
rect 491446 229041 491498 229093
rect 493942 229041 493994 229093
rect 510934 229041 510986 229093
rect 633526 229041 633578 229093
rect 649750 229041 649802 229093
rect 357814 228967 357866 229019
rect 367798 228967 367850 229019
rect 367894 228967 367946 229019
rect 380278 228967 380330 229019
rect 380566 228967 380618 229019
rect 169846 228893 169898 228945
rect 212854 228893 212906 228945
rect 284086 228893 284138 228945
rect 350326 228893 350378 228945
rect 178486 228819 178538 228871
rect 213238 228819 213290 228871
rect 286294 228819 286346 228871
rect 368470 228893 368522 228945
rect 370198 228893 370250 228945
rect 350518 228819 350570 228871
rect 184246 228745 184298 228797
rect 213526 228745 213578 228797
rect 286486 228745 286538 228797
rect 366262 228745 366314 228797
rect 204598 228671 204650 228723
rect 205846 228671 205898 228723
rect 192886 228597 192938 228649
rect 214294 228671 214346 228723
rect 285622 228671 285674 228723
rect 365878 228671 365930 228723
rect 366454 228819 366506 228871
rect 380662 228819 380714 228871
rect 367990 228745 368042 228797
rect 374422 228745 374474 228797
rect 376054 228745 376106 228797
rect 380566 228745 380618 228797
rect 349366 228597 349418 228649
rect 360982 228597 361034 228649
rect 361078 228597 361130 228649
rect 368374 228597 368426 228649
rect 370006 228671 370058 228723
rect 374806 228671 374858 228723
rect 384310 228819 384362 228871
rect 397462 228893 397514 228945
rect 397654 228893 397706 228945
rect 405622 228893 405674 228945
rect 410614 228893 410666 228945
rect 414262 228893 414314 228945
rect 414838 228893 414890 228945
rect 427894 228893 427946 228945
rect 427990 228893 428042 228945
rect 451318 228893 451370 228945
rect 452278 228893 452330 228945
rect 457558 228893 457610 228945
rect 477526 228967 477578 229019
rect 489238 228967 489290 229019
rect 497878 228967 497930 229019
rect 511318 228967 511370 229019
rect 541366 228967 541418 229019
rect 650902 228967 650954 229019
rect 490678 228893 490730 228945
rect 494998 228893 495050 228945
rect 510166 228893 510218 228945
rect 669526 228893 669578 228945
rect 674710 228893 674762 228945
rect 394294 228819 394346 228871
rect 393910 228745 393962 228797
rect 403222 228745 403274 228797
rect 403990 228819 404042 228871
rect 417526 228745 417578 228797
rect 388726 228671 388778 228723
rect 394198 228671 394250 228723
rect 398134 228671 398186 228723
rect 398326 228671 398378 228723
rect 412246 228671 412298 228723
rect 413686 228671 413738 228723
rect 418582 228671 418634 228723
rect 418774 228819 418826 228871
rect 456790 228819 456842 228871
rect 498070 228819 498122 228871
rect 511990 228819 512042 228871
rect 419158 228745 419210 228797
rect 456118 228745 456170 228797
rect 493750 228745 493802 228797
rect 509398 228745 509450 228797
rect 453142 228671 453194 228723
rect 432214 228597 432266 228649
rect 432406 228597 432458 228649
rect 434902 228597 434954 228649
rect 282742 228523 282794 228575
rect 352630 228523 352682 228575
rect 356278 228523 356330 228575
rect 367030 228523 367082 228575
rect 368950 228523 369002 228575
rect 372886 228523 372938 228575
rect 375382 228523 375434 228575
rect 378838 228523 378890 228575
rect 382870 228523 382922 228575
rect 403030 228523 403082 228575
rect 403222 228523 403274 228575
rect 410614 228523 410666 228575
rect 283606 228449 283658 228501
rect 361846 228449 361898 228501
rect 372790 228449 372842 228501
rect 378454 228449 378506 228501
rect 346102 228375 346154 228427
rect 394198 228449 394250 228501
rect 403318 228449 403370 228501
rect 411286 228449 411338 228501
rect 390262 228375 390314 228427
rect 399382 228375 399434 228427
rect 409654 228375 409706 228427
rect 420022 228523 420074 228575
rect 426262 228523 426314 228575
rect 450550 228597 450602 228649
rect 499606 228597 499658 228649
rect 514198 228597 514250 228649
rect 438934 228523 438986 228575
rect 475990 228523 476042 228575
rect 411478 228449 411530 228501
rect 434902 228449 434954 228501
rect 434998 228449 435050 228501
rect 439030 228449 439082 228501
rect 440086 228449 440138 228501
rect 452758 228449 452810 228501
rect 459286 228449 459338 228501
rect 509110 228449 509162 228501
rect 411574 228375 411626 228427
rect 416566 228375 416618 228427
rect 418582 228375 418634 228427
rect 204694 228301 204746 228353
rect 205078 228301 205130 228353
rect 206614 228301 206666 228353
rect 284278 228301 284330 228353
rect 346774 228301 346826 228353
rect 358390 228301 358442 228353
rect 350326 228227 350378 228279
rect 368086 228301 368138 228353
rect 368182 228301 368234 228353
rect 382102 228301 382154 228353
rect 395062 228301 395114 228353
rect 399094 228301 399146 228353
rect 402934 228301 402986 228353
rect 418774 228301 418826 228353
rect 423478 228375 423530 228427
rect 435958 228375 436010 228427
rect 428182 228301 428234 228353
rect 428662 228301 428714 228353
rect 472630 228375 472682 228427
rect 439126 228301 439178 228353
rect 469654 228301 469706 228353
rect 360022 228227 360074 228279
rect 411382 228227 411434 228279
rect 411670 228227 411722 228279
rect 423094 228227 423146 228279
rect 431734 228227 431786 228279
rect 438934 228227 438986 228279
rect 439222 228227 439274 228279
rect 471862 228227 471914 228279
rect 499702 228227 499754 228279
rect 513526 228227 513578 228279
rect 360790 228153 360842 228205
rect 360886 228153 360938 228205
rect 431158 228153 431210 228205
rect 432598 228153 432650 228205
rect 447190 228153 447242 228205
rect 447382 228153 447434 228205
rect 474454 228153 474506 228205
rect 283798 228079 283850 228131
rect 357814 228079 357866 228131
rect 358582 228079 358634 228131
rect 434998 228079 435050 228131
rect 440758 228079 440810 228131
rect 459766 228079 459818 228131
rect 354934 228005 354986 228057
rect 360886 228005 360938 228057
rect 360982 228005 361034 228057
rect 414838 228005 414890 228057
rect 414934 228005 414986 228057
rect 423286 228005 423338 228057
rect 431830 228005 431882 228057
rect 435766 228005 435818 228057
rect 435862 228005 435914 228057
rect 440854 228005 440906 228057
rect 352054 227931 352106 227983
rect 358486 227931 358538 227983
rect 358678 227931 358730 227983
rect 369238 227931 369290 227983
rect 378646 227931 378698 227983
rect 435190 227931 435242 227983
rect 351574 227857 351626 227909
rect 432118 227857 432170 227909
rect 432310 227857 432362 227909
rect 440566 227931 440618 227983
rect 449782 228005 449834 228057
rect 459382 228005 459434 228057
rect 477046 227931 477098 227983
rect 351190 227783 351242 227835
rect 432886 227783 432938 227835
rect 204502 227709 204554 227761
rect 206902 227709 206954 227761
rect 207766 227709 207818 227761
rect 242038 227709 242090 227761
rect 350902 227709 350954 227761
rect 432310 227709 432362 227761
rect 434038 227709 434090 227761
rect 435574 227709 435626 227761
rect 144118 227635 144170 227687
rect 149398 227635 149450 227687
rect 204982 227635 205034 227687
rect 207286 227635 207338 227687
rect 207862 227635 207914 227687
rect 293398 227635 293450 227687
rect 139990 227561 140042 227613
rect 140278 227561 140330 227613
rect 144022 227561 144074 227613
rect 177046 227561 177098 227613
rect 199990 227561 200042 227613
rect 204790 227561 204842 227613
rect 206230 227561 206282 227613
rect 221878 227561 221930 227613
rect 242038 227561 242090 227613
rect 358966 227635 359018 227687
rect 359158 227635 359210 227687
rect 432022 227635 432074 227687
rect 432982 227635 433034 227687
rect 441142 227857 441194 227909
rect 447382 227857 447434 227909
rect 447478 227857 447530 227909
rect 475222 227857 475274 227909
rect 669622 227857 669674 227909
rect 674422 227857 674474 227909
rect 435766 227783 435818 227835
rect 449782 227783 449834 227835
rect 435766 227635 435818 227687
rect 502486 227709 502538 227761
rect 437494 227635 437546 227687
rect 506134 227635 506186 227687
rect 506902 227635 506954 227687
rect 512758 227635 512810 227687
rect 200086 227487 200138 227539
rect 208150 227487 208202 227539
rect 221782 227487 221834 227539
rect 242038 227339 242090 227391
rect 357526 227561 357578 227613
rect 360022 227487 360074 227539
rect 360598 227487 360650 227539
rect 378646 227561 378698 227613
rect 386902 227561 386954 227613
rect 398902 227561 398954 227613
rect 399094 227561 399146 227613
rect 408118 227561 408170 227613
rect 415990 227561 416042 227613
rect 423190 227561 423242 227613
rect 430390 227561 430442 227613
rect 435862 227561 435914 227613
rect 435958 227561 436010 227613
rect 461974 227561 462026 227613
rect 501046 227561 501098 227613
rect 539638 227561 539690 227613
rect 541366 227561 541418 227613
rect 384022 227487 384074 227539
rect 391606 227487 391658 227539
rect 403222 227487 403274 227539
rect 409654 227487 409706 227539
rect 329206 227413 329258 227465
rect 348214 227413 348266 227465
rect 348502 227413 348554 227465
rect 418582 227487 418634 227539
rect 418678 227487 418730 227539
rect 432790 227487 432842 227539
rect 432886 227487 432938 227539
rect 441334 227487 441386 227539
rect 441430 227487 441482 227539
rect 455734 227487 455786 227539
rect 346678 227339 346730 227391
rect 418102 227413 418154 227465
rect 418774 227413 418826 227465
rect 431830 227413 431882 227465
rect 432118 227413 432170 227465
rect 440662 227413 440714 227465
rect 409942 227339 409994 227391
rect 422902 227339 422954 227391
rect 423382 227339 423434 227391
rect 430678 227339 430730 227391
rect 432310 227339 432362 227391
rect 442102 227339 442154 227391
rect 344278 227265 344330 227317
rect 326806 227191 326858 227243
rect 409846 227191 409898 227243
rect 315958 227117 316010 227169
rect 414646 227191 414698 227243
rect 414838 227265 414890 227317
rect 422806 227265 422858 227317
rect 423478 227265 423530 227317
rect 431446 227265 431498 227317
rect 432214 227265 432266 227317
rect 442870 227265 442922 227317
rect 434710 227191 434762 227243
rect 434902 227191 434954 227243
rect 527158 227339 527210 227391
rect 443062 227191 443114 227243
rect 450166 227191 450218 227243
rect 410038 227117 410090 227169
rect 422998 227117 423050 227169
rect 423286 227117 423338 227169
rect 446614 227117 446666 227169
rect 316630 227043 316682 227095
rect 422614 227043 422666 227095
rect 423382 227043 423434 227095
rect 429622 227043 429674 227095
rect 439030 227043 439082 227095
rect 458998 227043 459050 227095
rect 315190 226969 315242 227021
rect 423286 226969 423338 227021
rect 432790 226969 432842 227021
rect 437494 226969 437546 227021
rect 437590 226969 437642 227021
rect 464182 226969 464234 227021
rect 333910 226895 333962 226947
rect 429526 226895 429578 226947
rect 432118 226895 432170 226947
rect 443062 226895 443114 226947
rect 326614 226821 326666 226873
rect 418774 226821 418826 226873
rect 418870 226821 418922 226873
rect 429046 226821 429098 226873
rect 348214 226747 348266 226799
rect 317782 226673 317834 226725
rect 418678 226673 418730 226725
rect 419062 226747 419114 226799
rect 438166 226821 438218 226873
rect 429718 226747 429770 226799
rect 446710 226747 446762 226799
rect 318454 226599 318506 226651
rect 418870 226599 418922 226651
rect 307126 226525 307178 226577
rect 426070 226599 426122 226651
rect 419734 226525 419786 226577
rect 428470 226599 428522 226651
rect 429334 226673 429386 226725
rect 452374 226673 452426 226725
rect 433750 226599 433802 226651
rect 435382 226599 435434 226651
rect 439318 226599 439370 226651
rect 426262 226525 426314 226577
rect 319222 226451 319274 226503
rect 418870 226451 418922 226503
rect 419158 226451 419210 226503
rect 420790 226451 420842 226503
rect 422998 226451 423050 226503
rect 305590 226377 305642 226429
rect 409942 226377 409994 226429
rect 307798 226303 307850 226355
rect 427030 226377 427082 226429
rect 304150 226229 304202 226281
rect 410038 226229 410090 226281
rect 306358 226155 306410 226207
rect 427702 226303 427754 226355
rect 428374 226451 428426 226503
rect 428854 226303 428906 226355
rect 410326 226229 410378 226281
rect 426454 226229 426506 226281
rect 410614 226155 410666 226207
rect 412150 226155 412202 226207
rect 413206 226155 413258 226207
rect 435862 226303 435914 226355
rect 429238 226229 429290 226281
rect 429718 226229 429770 226281
rect 431830 226229 431882 226281
rect 438934 226229 438986 226281
rect 527062 226525 527114 226577
rect 460534 226229 460586 226281
rect 429526 226155 429578 226207
rect 448726 226155 448778 226207
rect 304918 226081 304970 226133
rect 418678 226081 418730 226133
rect 418774 226081 418826 226133
rect 425302 226081 425354 226133
rect 425398 226081 425450 226133
rect 439030 226081 439082 226133
rect 439318 226081 439370 226133
rect 484054 226081 484106 226133
rect 359830 226007 359882 226059
rect 413206 226007 413258 226059
rect 355030 225933 355082 225985
rect 418870 226007 418922 226059
rect 358774 225859 358826 225911
rect 418870 225859 418922 225911
rect 434326 225933 434378 225985
rect 434998 226007 435050 226059
rect 454294 226007 454346 226059
rect 436246 225933 436298 225985
rect 362422 225785 362474 225837
rect 436534 225859 436586 225911
rect 419446 225785 419498 225837
rect 419734 225785 419786 225837
rect 420118 225785 420170 225837
rect 425878 225785 425930 225837
rect 426262 225785 426314 225837
rect 427414 225785 427466 225837
rect 427510 225785 427562 225837
rect 432502 225785 432554 225837
rect 352150 225711 352202 225763
rect 410326 225711 410378 225763
rect 410422 225711 410474 225763
rect 420886 225711 420938 225763
rect 362326 225637 362378 225689
rect 411286 225637 411338 225689
rect 411382 225637 411434 225689
rect 415606 225637 415658 225689
rect 417238 225637 417290 225689
rect 418870 225637 418922 225689
rect 419062 225637 419114 225689
rect 419254 225637 419306 225689
rect 437302 225711 437354 225763
rect 351670 225563 351722 225615
rect 418774 225563 418826 225615
rect 429622 225637 429674 225689
rect 437782 225711 437834 225763
rect 457174 225711 457226 225763
rect 512662 225711 512714 225763
rect 360694 225489 360746 225541
rect 418966 225489 419018 225541
rect 420694 225489 420746 225541
rect 420982 225563 421034 225615
rect 424822 225563 424874 225615
rect 426358 225563 426410 225615
rect 521398 225563 521450 225615
rect 433654 225489 433706 225541
rect 433750 225489 433802 225541
rect 443926 225489 443978 225541
rect 354742 225415 354794 225467
rect 420790 225415 420842 225467
rect 425206 225415 425258 225467
rect 354838 225341 354890 225393
rect 420118 225341 420170 225393
rect 355126 225267 355178 225319
rect 420214 225267 420266 225319
rect 365110 225193 365162 225245
rect 421462 225341 421514 225393
rect 422902 225341 422954 225393
rect 427798 225415 427850 225467
rect 427894 225415 427946 225467
rect 445078 225415 445130 225467
rect 426262 225341 426314 225393
rect 489718 225341 489770 225393
rect 363574 225119 363626 225171
rect 421846 225267 421898 225319
rect 423574 225267 423626 225319
rect 431062 225267 431114 225319
rect 431542 225267 431594 225319
rect 433078 225267 433130 225319
rect 438934 225267 438986 225319
rect 442102 225267 442154 225319
rect 420502 225193 420554 225245
rect 435478 225193 435530 225245
rect 366742 225045 366794 225097
rect 420310 225045 420362 225097
rect 363478 224971 363530 225023
rect 422230 225119 422282 225171
rect 423094 225119 423146 225171
rect 448150 225119 448202 225171
rect 420598 225045 420650 225097
rect 434038 225045 434090 225097
rect 421942 224971 421994 225023
rect 435094 224971 435146 225023
rect 368374 224897 368426 224949
rect 381334 224897 381386 224949
rect 395158 224897 395210 224949
rect 444694 224971 444746 225023
rect 436438 224897 436490 224949
rect 449110 224897 449162 224949
rect 359926 224823 359978 224875
rect 374998 224823 375050 224875
rect 395254 224823 395306 224875
rect 443158 224823 443210 224875
rect 394582 224749 394634 224801
rect 441334 224749 441386 224801
rect 144022 224675 144074 224727
rect 174166 224675 174218 224727
rect 348886 224675 348938 224727
rect 424438 224675 424490 224727
rect 395830 224601 395882 224653
rect 405718 224601 405770 224653
rect 417718 224601 417770 224653
rect 418006 224601 418058 224653
rect 418102 224601 418154 224653
rect 424054 224601 424106 224653
rect 374998 224527 375050 224579
rect 420790 224527 420842 224579
rect 420886 224527 420938 224579
rect 425782 224675 425834 224727
rect 426550 224675 426602 224727
rect 426166 224601 426218 224653
rect 432118 224675 432170 224727
rect 432598 224675 432650 224727
rect 452470 224675 452522 224727
rect 430390 224601 430442 224653
rect 433462 224601 433514 224653
rect 426646 224527 426698 224579
rect 427318 224527 427370 224579
rect 428182 224527 428234 224579
rect 429046 224527 429098 224579
rect 438070 224527 438122 224579
rect 354262 224453 354314 224505
rect 438742 224453 438794 224505
rect 354454 224379 354506 224431
rect 421078 224379 421130 224431
rect 422326 224379 422378 224431
rect 436918 224379 436970 224431
rect 351382 224305 351434 224357
rect 439126 224305 439178 224357
rect 325846 224157 325898 224209
rect 338326 224157 338378 224209
rect 364630 224231 364682 224283
rect 391894 224231 391946 224283
rect 444310 224231 444362 224283
rect 351478 224157 351530 224209
rect 328054 224009 328106 224061
rect 363862 224083 363914 224135
rect 364342 224083 364394 224135
rect 396022 224157 396074 224209
rect 405430 224157 405482 224209
rect 405718 224157 405770 224209
rect 439510 224157 439562 224209
rect 348598 224009 348650 224061
rect 364630 224009 364682 224061
rect 378550 224009 378602 224061
rect 395830 224083 395882 224135
rect 395926 224083 395978 224135
rect 417718 224083 417770 224135
rect 427318 224083 427370 224135
rect 418102 224009 418154 224061
rect 427606 224009 427658 224061
rect 207382 223935 207434 223987
rect 379318 223935 379370 223987
rect 403222 223935 403274 223987
rect 405142 223935 405194 223987
rect 406102 223935 406154 223987
rect 418006 223935 418058 223987
rect 418198 223935 418250 223987
rect 418486 223935 418538 223987
rect 442486 224083 442538 224135
rect 428182 224009 428234 224061
rect 440278 224009 440330 224061
rect 204310 223787 204362 223839
rect 330454 223861 330506 223913
rect 363862 223861 363914 223913
rect 364342 223861 364394 223913
rect 396022 223861 396074 223913
rect 405430 223861 405482 223913
rect 418102 223861 418154 223913
rect 427606 223861 427658 223913
rect 207670 223787 207722 223839
rect 330262 223787 330314 223839
rect 338326 223787 338378 223839
rect 364246 223787 364298 223839
rect 378550 223787 378602 223839
rect 379318 223787 379370 223839
rect 379414 223787 379466 223839
rect 417910 223787 417962 223839
rect 418006 223787 418058 223839
rect 441718 223787 441770 223839
rect 443590 223787 443642 223839
rect 445078 223787 445130 223839
rect 451798 223787 451850 223839
rect 452038 223787 452090 223839
rect 483862 223787 483914 223839
rect 503206 223787 503258 223839
rect 204502 223195 204554 223247
rect 204502 223047 204554 223099
rect 204982 223047 205034 223099
rect 204886 222825 204938 222877
rect 641014 222381 641066 222433
rect 649654 222381 649706 222433
rect 144022 221789 144074 221841
rect 171286 221789 171338 221841
rect 199990 221789 200042 221841
rect 200086 221789 200138 221841
rect 141526 221715 141578 221767
rect 198742 221715 198794 221767
rect 641302 221345 641354 221397
rect 650326 221345 650378 221397
rect 42358 221049 42410 221101
rect 45718 221049 45770 221101
rect 641302 220753 641354 220805
rect 650038 220753 650090 220805
rect 42358 220309 42410 220361
rect 45814 220309 45866 220361
rect 42358 219421 42410 219473
rect 45526 219421 45578 219473
rect 144118 218977 144170 219029
rect 149590 218977 149642 219029
rect 144022 218903 144074 218955
rect 165526 218903 165578 218955
rect 141910 218829 141962 218881
rect 199030 218829 199082 218881
rect 142198 218755 142250 218807
rect 198742 218755 198794 218807
rect 140854 218681 140906 218733
rect 198838 218681 198890 218733
rect 149686 218607 149738 218659
rect 198934 218607 198986 218659
rect 155446 218533 155498 218585
rect 198742 218533 198794 218585
rect 144022 218015 144074 218067
rect 159766 218015 159818 218067
rect 141334 215943 141386 215995
rect 199030 215943 199082 215995
rect 141718 215869 141770 215921
rect 198934 215869 198986 215921
rect 164086 215795 164138 215847
rect 198742 215795 198794 215847
rect 175606 215721 175658 215773
rect 198838 215721 198890 215773
rect 181366 215647 181418 215699
rect 198742 215647 198794 215699
rect 187126 215573 187178 215625
rect 198838 215573 198890 215625
rect 144022 213205 144074 213257
rect 154006 213205 154058 213257
rect 146518 213131 146570 213183
rect 148342 213131 148394 213183
rect 139990 213057 140042 213109
rect 198742 213057 198794 213109
rect 144022 210245 144074 210297
rect 185686 210245 185738 210297
rect 639766 210245 639818 210297
rect 679702 210245 679754 210297
rect 144022 207359 144074 207411
rect 148054 207359 148106 207411
rect 204598 207359 204650 207411
rect 204886 207359 204938 207411
rect 674518 205731 674570 205783
rect 675478 205731 675530 205783
rect 146806 205139 146858 205191
rect 156886 205139 156938 205191
rect 675094 204991 675146 205043
rect 675190 204991 675242 205043
rect 675478 204991 675530 205043
rect 674998 204769 675050 204821
rect 146806 204473 146858 204525
rect 182806 204473 182858 204525
rect 42358 204325 42410 204377
rect 44566 204325 44618 204377
rect 144982 201587 145034 201639
rect 179926 201587 179978 201639
rect 200662 201513 200714 201565
rect 200950 201513 201002 201565
rect 42070 201291 42122 201343
rect 42934 201291 42986 201343
rect 674422 201291 674474 201343
rect 675382 201291 675434 201343
rect 37366 200773 37418 200825
rect 41782 200773 41834 200825
rect 42742 198849 42794 198901
rect 43318 198849 43370 198901
rect 42838 198775 42890 198827
rect 43222 198775 43274 198827
rect 144982 198775 145034 198827
rect 162646 198775 162698 198827
rect 144406 198701 144458 198753
rect 197302 198701 197354 198753
rect 41878 198183 41930 198235
rect 42358 198183 42410 198235
rect 674806 197591 674858 197643
rect 675382 197591 675434 197643
rect 41974 197443 42026 197495
rect 42454 197443 42506 197495
rect 41782 197369 41834 197421
rect 41782 197147 41834 197199
rect 674134 196999 674186 197051
rect 675478 196999 675530 197051
rect 674710 196555 674762 196607
rect 675382 196555 675434 196607
rect 639574 195815 639626 195867
rect 639958 195815 640010 195867
rect 42166 195297 42218 195349
rect 42358 195297 42410 195349
rect 42358 195149 42410 195201
rect 43222 195149 43274 195201
rect 42070 194483 42122 194535
rect 47638 194483 47690 194535
rect 42070 193447 42122 193499
rect 43318 193447 43370 193499
rect 144598 193077 144650 193129
rect 148534 193077 148586 193129
rect 146806 193003 146858 193055
rect 191542 193003 191594 193055
rect 42166 192189 42218 192241
rect 43030 192189 43082 192241
rect 42070 191449 42122 191501
rect 42358 191449 42410 191501
rect 42166 191005 42218 191057
rect 43126 191005 43178 191057
rect 144310 190117 144362 190169
rect 188662 190117 188714 190169
rect 42262 189229 42314 189281
rect 42646 189229 42698 189281
rect 42166 187823 42218 187875
rect 42742 187823 42794 187875
rect 146806 187231 146858 187283
rect 185782 187231 185834 187283
rect 200758 187231 200810 187283
rect 201046 187231 201098 187283
rect 42166 187083 42218 187135
rect 42646 187083 42698 187135
rect 42070 186639 42122 186691
rect 42454 186639 42506 186691
rect 146806 184419 146858 184471
rect 180022 184419 180074 184471
rect 146614 184345 146666 184397
rect 182902 184345 182954 184397
rect 655318 184345 655370 184397
rect 674422 184345 674474 184397
rect 661174 183901 661226 183953
rect 674710 183901 674762 183953
rect 144982 182865 145034 182917
rect 146518 182865 146570 182917
rect 666742 182865 666794 182917
rect 674422 182865 674474 182917
rect 144694 181533 144746 181585
rect 148918 181533 148970 181585
rect 146806 181459 146858 181511
rect 168502 181459 168554 181511
rect 200662 181459 200714 181511
rect 200854 181459 200906 181511
rect 144886 181311 144938 181363
rect 146806 181311 146858 181363
rect 144022 178573 144074 178625
rect 177142 178573 177194 178625
rect 144982 175761 145034 175813
rect 149014 175761 149066 175813
rect 144982 172801 145034 172853
rect 149302 172801 149354 172853
rect 144982 169915 145034 169967
rect 151222 169915 151274 169967
rect 144982 167843 145034 167895
rect 156982 167843 157034 167895
rect 641494 167177 641546 167229
rect 674710 167177 674762 167229
rect 144982 167029 145034 167081
rect 149494 167029 149546 167081
rect 144982 164217 145034 164269
rect 149686 164217 149738 164269
rect 642166 164217 642218 164269
rect 674710 164217 674762 164269
rect 144022 164143 144074 164195
rect 194422 164143 194474 164195
rect 642070 164143 642122 164195
rect 674614 164143 674666 164195
rect 675190 163033 675242 163085
rect 676918 163033 676970 163085
rect 675094 162071 675146 162123
rect 676822 162071 676874 162123
rect 144310 161405 144362 161457
rect 148150 161405 148202 161457
rect 144982 161331 145034 161383
rect 171382 161331 171434 161383
rect 144214 161257 144266 161309
rect 174262 161257 174314 161309
rect 144502 161109 144554 161161
rect 144886 161109 144938 161161
rect 675670 160961 675722 161013
rect 674422 160739 674474 160791
rect 675382 160739 675434 160791
rect 675670 159999 675722 160051
rect 144310 158445 144362 158497
rect 147958 158445 148010 158497
rect 674902 157039 674954 157091
rect 675094 157039 675146 157091
rect 674806 156891 674858 156943
rect 675478 156891 675530 156943
rect 144310 156003 144362 156055
rect 149110 156003 149162 156055
rect 144502 155559 144554 155611
rect 165622 155559 165674 155611
rect 144502 152747 144554 152799
rect 159862 152747 159914 152799
rect 144310 152673 144362 152725
rect 202966 152673 203018 152725
rect 674230 152599 674282 152651
rect 675382 152599 675434 152651
rect 674038 152007 674090 152059
rect 675478 152007 675530 152059
rect 674518 151489 674570 151541
rect 675382 151489 675434 151541
rect 144310 149861 144362 149913
rect 154102 149861 154154 149913
rect 144502 149787 144554 149839
rect 203062 149787 203114 149839
rect 640150 149787 640202 149839
rect 643606 149787 643658 149839
rect 144214 149047 144266 149099
rect 144502 149047 144554 149099
rect 144502 147123 144554 147175
rect 144214 147049 144266 147101
rect 147862 147049 147914 147101
rect 144310 146975 144362 147027
rect 162742 146975 162794 147027
rect 144214 146901 144266 146953
rect 144502 146901 144554 146953
rect 163030 146901 163082 146953
rect 144310 144089 144362 144141
rect 147766 144089 147818 144141
rect 144502 144015 144554 144067
rect 162838 144015 162890 144067
rect 642166 142535 642218 142587
rect 674326 142609 674378 142661
rect 679702 142609 679754 142661
rect 144502 142239 144554 142291
rect 157078 142239 157130 142291
rect 144310 141129 144362 141181
rect 203158 141129 203210 141181
rect 143926 139427 143978 139479
rect 144214 139427 144266 139479
rect 655222 138539 655274 138591
rect 674710 138539 674762 138591
rect 144214 138391 144266 138443
rect 151318 138391 151370 138443
rect 655126 138391 655178 138443
rect 674422 138391 674474 138443
rect 144310 138317 144362 138369
rect 162934 138317 162986 138369
rect 144406 138243 144458 138295
rect 144502 138243 144554 138295
rect 203254 138243 203306 138295
rect 143926 138021 143978 138073
rect 144310 138021 144362 138073
rect 144406 138021 144458 138073
rect 655414 135579 655466 135631
rect 674710 135579 674762 135631
rect 144214 135505 144266 135557
rect 144118 135431 144170 135483
rect 197398 135431 197450 135483
rect 203350 135357 203402 135409
rect 640726 135357 640778 135409
rect 674710 135357 674762 135409
rect 144022 132619 144074 132671
rect 147670 132619 147722 132671
rect 144214 132545 144266 132597
rect 194518 132545 194570 132597
rect 144118 132471 144170 132523
rect 204982 132471 205034 132523
rect 643606 132471 643658 132523
rect 674422 132471 674474 132523
rect 144118 129659 144170 129711
rect 191638 129659 191690 129711
rect 144214 129585 144266 129637
rect 203446 129585 203498 129637
rect 144118 126773 144170 126825
rect 188758 126773 188810 126825
rect 144214 126699 144266 126751
rect 203542 126699 203594 126751
rect 200854 126625 200906 126677
rect 201046 126625 201098 126677
rect 144214 124035 144266 124087
rect 185878 124035 185930 124087
rect 144022 123961 144074 124013
rect 203734 123961 203786 124013
rect 144118 123887 144170 123939
rect 203638 123887 203690 123939
rect 642070 121223 642122 121275
rect 674710 121223 674762 121275
rect 642166 121149 642218 121201
rect 674806 121149 674858 121201
rect 641398 121075 641450 121127
rect 674614 121075 674666 121127
rect 144214 121001 144266 121053
rect 203830 121001 203882 121053
rect 200470 120927 200522 120979
rect 200758 120927 200810 120979
rect 200854 120927 200906 120979
rect 201046 120927 201098 120979
rect 674902 119521 674954 119573
rect 675094 119521 675146 119573
rect 674134 118485 674186 118537
rect 675286 118485 675338 118537
rect 144214 118263 144266 118315
rect 180118 118263 180170 118315
rect 144118 118189 144170 118241
rect 182998 118189 183050 118241
rect 144022 118115 144074 118167
rect 203926 118115 203978 118167
rect 144214 115303 144266 115355
rect 168598 115303 168650 115355
rect 144118 115229 144170 115281
rect 204022 115229 204074 115281
rect 674902 114785 674954 114837
rect 675094 114785 675146 114837
rect 674134 114119 674186 114171
rect 675382 114119 675434 114171
rect 674230 113601 674282 113653
rect 675190 113601 675242 113653
rect 674518 113305 674570 113357
rect 675094 113305 675146 113357
rect 144214 112417 144266 112469
rect 204118 112417 204170 112469
rect 144118 112343 144170 112395
rect 204886 112343 204938 112395
rect 674422 111159 674474 111211
rect 675382 111159 675434 111211
rect 144214 109605 144266 109657
rect 174358 109605 174410 109657
rect 144022 109531 144074 109583
rect 177238 109531 177290 109583
rect 144118 109457 144170 109509
rect 204214 109457 204266 109509
rect 674806 107533 674858 107585
rect 675382 107533 675434 107585
rect 674038 106867 674090 106919
rect 675478 106867 675530 106919
rect 144214 106571 144266 106623
rect 171478 106571 171530 106623
rect 200470 106497 200522 106549
rect 200662 106497 200714 106549
rect 674614 106349 674666 106401
rect 675382 106349 675434 106401
rect 674326 105165 674378 105217
rect 675382 105165 675434 105217
rect 144118 103833 144170 103885
rect 165718 103833 165770 103885
rect 144214 103759 144266 103811
rect 202774 103759 202826 103811
rect 144022 103685 144074 103737
rect 202870 103685 202922 103737
rect 144214 100799 144266 100851
rect 202678 100799 202730 100851
rect 652534 100799 652586 100851
rect 668182 100799 668234 100851
rect 144214 97913 144266 97965
rect 202582 97913 202634 97965
rect 204982 96507 205034 96559
rect 204886 96285 204938 96337
rect 663286 96433 663338 96485
rect 665206 96433 665258 96485
rect 144118 95101 144170 95153
rect 202198 95101 202250 95153
rect 144214 95027 144266 95079
rect 201814 95027 201866 95079
rect 197206 94953 197258 95005
rect 198742 94953 198794 95005
rect 191446 94879 191498 94931
rect 198934 94879 198986 94931
rect 144214 93547 144266 93599
rect 149782 93547 149834 93599
rect 635254 92807 635306 92859
rect 662518 92807 662570 92859
rect 635062 92733 635114 92785
rect 663094 92733 663146 92785
rect 641014 92659 641066 92711
rect 659830 92659 659882 92711
rect 635350 92585 635402 92637
rect 658870 92585 658922 92637
rect 634966 92511 635018 92563
rect 658294 92511 658346 92563
rect 635446 92437 635498 92489
rect 659350 92437 659402 92489
rect 635158 92363 635210 92415
rect 661174 92363 661226 92415
rect 634006 92289 634058 92341
rect 660694 92289 660746 92341
rect 640726 92215 640778 92267
rect 661750 92215 661802 92267
rect 152662 92141 152714 92193
rect 198838 92141 198890 92193
rect 640822 92141 640874 92193
rect 657526 92141 657578 92193
rect 151126 92067 151178 92119
rect 198742 92067 198794 92119
rect 156886 91993 156938 92045
rect 199030 91993 199082 92045
rect 188566 91919 188618 91971
rect 199126 91919 199178 91971
rect 185686 91845 185738 91897
rect 198838 91845 198890 91897
rect 182806 91771 182858 91823
rect 198934 91771 198986 91823
rect 144214 90587 144266 90639
rect 160246 90587 160298 90639
rect 144214 89255 144266 89307
rect 163126 89255 163178 89307
rect 168406 89181 168458 89233
rect 198934 89181 198986 89233
rect 174166 89107 174218 89159
rect 199030 89107 199082 89159
rect 177046 89033 177098 89085
rect 198838 89033 198890 89085
rect 179926 88959 179978 89011
rect 198742 88959 198794 89011
rect 194326 88885 194378 88937
rect 199222 88885 199274 88937
rect 635542 87775 635594 87827
rect 652534 87775 652586 87827
rect 144214 87035 144266 87087
rect 144118 86517 144170 86569
rect 163222 86517 163274 86569
rect 202582 86517 202634 86569
rect 204886 86517 204938 86569
rect 144214 86443 144266 86495
rect 202390 86443 202442 86495
rect 640918 86443 640970 86495
rect 652630 86443 652682 86495
rect 144118 86369 144170 86421
rect 151222 86369 151274 86421
rect 199222 86369 199274 86421
rect 200854 86369 200906 86421
rect 201046 86369 201098 86421
rect 154006 86295 154058 86347
rect 199126 86295 199178 86347
rect 202198 86295 202250 86347
rect 202582 86295 202634 86347
rect 159766 86221 159818 86273
rect 198934 86221 198986 86273
rect 162646 86147 162698 86199
rect 199030 86147 199082 86199
rect 165526 86073 165578 86125
rect 198742 86073 198794 86125
rect 171286 85999 171338 86051
rect 198838 85999 198890 86051
rect 146902 83779 146954 83831
rect 163606 83779 163658 83831
rect 641110 83705 641162 83757
rect 653590 83705 653642 83757
rect 144118 83631 144170 83683
rect 163318 83631 163370 83683
rect 635638 83631 635690 83683
rect 653686 83631 653738 83683
rect 635734 83557 635786 83609
rect 653494 83557 653546 83609
rect 146902 83483 146954 83535
rect 148726 83483 148778 83535
rect 197302 83483 197354 83535
rect 200758 83483 200810 83535
rect 194422 83409 194474 83461
rect 199510 83409 199562 83461
rect 191542 83335 191594 83387
rect 198838 83335 198890 83387
rect 188662 83261 188714 83313
rect 198934 83261 198986 83313
rect 156982 83187 157034 83239
rect 198742 83187 198794 83239
rect 146998 82151 147050 82203
rect 160054 82151 160106 82203
rect 640630 81041 640682 81093
rect 663286 81041 663338 81093
rect 641302 80893 641354 80945
rect 663478 80893 663530 80945
rect 635926 80745 635978 80797
rect 662422 80819 662474 80871
rect 641206 80745 641258 80797
rect 653686 80745 653738 80797
rect 144118 80671 144170 80723
rect 162646 80671 162698 80723
rect 201814 80671 201866 80723
rect 202102 80671 202154 80723
rect 635830 80671 635882 80723
rect 640630 80671 640682 80723
rect 641398 80671 641450 80723
rect 653590 80671 653642 80723
rect 168502 80597 168554 80649
rect 198934 80597 198986 80649
rect 177142 80523 177194 80575
rect 199030 80523 199082 80575
rect 180022 80449 180074 80501
rect 198838 80449 198890 80501
rect 185782 80375 185834 80427
rect 198742 80375 198794 80427
rect 182902 80227 182954 80279
rect 198742 80227 198794 80279
rect 144214 78599 144266 78651
rect 144118 77859 144170 77911
rect 163414 77859 163466 77911
rect 144214 77785 144266 77837
rect 163510 77785 163562 77837
rect 144118 77711 144170 77763
rect 149110 77711 149162 77763
rect 199126 77711 199178 77763
rect 641494 77711 641546 77763
rect 657526 77711 657578 77763
rect 149014 77637 149066 77689
rect 198742 77637 198794 77689
rect 642166 77637 642218 77689
rect 663766 77637 663818 77689
rect 149782 77563 149834 77615
rect 198934 77563 198986 77615
rect 165622 77489 165674 77541
rect 199030 77489 199082 77541
rect 171382 77415 171434 77467
rect 198838 77415 198890 77467
rect 174262 77341 174314 77393
rect 198742 77341 198794 77393
rect 144214 77267 144266 77319
rect 155542 77267 155594 77319
rect 641590 76897 641642 76949
rect 659638 76897 659690 76949
rect 636310 76749 636362 76801
rect 658294 76823 658346 76875
rect 641686 76749 641738 76801
rect 658870 76749 658922 76801
rect 636022 76675 636074 76727
rect 656950 76675 657002 76727
rect 636214 76601 636266 76653
rect 660694 76601 660746 76653
rect 636118 76527 636170 76579
rect 661174 76527 661226 76579
rect 634774 76453 634826 76505
rect 661750 76453 661802 76505
rect 634870 76379 634922 76431
rect 660118 76379 660170 76431
rect 636406 76305 636458 76357
rect 662518 76305 662570 76357
rect 144214 75343 144266 75395
rect 159766 75343 159818 75395
rect 144022 75195 144074 75247
rect 144214 75195 144266 75247
rect 143926 74973 143978 75025
rect 144118 74973 144170 75025
rect 146902 74899 146954 74951
rect 151126 74899 151178 74951
rect 154102 74825 154154 74877
rect 198934 74825 198986 74877
rect 157078 74751 157130 74803
rect 199126 74751 199178 74803
rect 160246 74677 160298 74729
rect 199030 74677 199082 74729
rect 159862 74603 159914 74655
rect 198742 74603 198794 74655
rect 163030 74529 163082 74581
rect 198838 74529 198890 74581
rect 143926 73715 143978 73767
rect 159958 73715 160010 73767
rect 143926 72013 143978 72065
rect 160150 72013 160202 72065
rect 197398 71939 197450 71991
rect 200758 71939 200810 71991
rect 194518 71865 194570 71917
rect 199606 71865 199658 71917
rect 191638 71791 191690 71843
rect 198838 71791 198890 71843
rect 188758 71717 188810 71769
rect 198934 71717 198986 71769
rect 151318 71643 151370 71695
rect 198742 71643 198794 71695
rect 146902 70015 146954 70067
rect 159862 70015 159914 70067
rect 147478 69053 147530 69105
rect 199030 69053 199082 69105
rect 168598 68979 168650 69031
rect 199126 68979 199178 69031
rect 180118 68905 180170 68957
rect 198934 68905 198986 68957
rect 185878 68831 185930 68883
rect 198838 68831 198890 68883
rect 182998 68757 183050 68809
rect 198742 68757 198794 68809
rect 143926 66907 143978 66959
rect 160246 66907 160298 66959
rect 143926 66759 143978 66811
rect 160342 66759 160394 66811
rect 200854 66315 200906 66367
rect 143830 66241 143882 66293
rect 167062 66241 167114 66293
rect 201046 66241 201098 66293
rect 147382 66167 147434 66219
rect 199126 66167 199178 66219
rect 147286 66093 147338 66145
rect 199222 66093 199274 66145
rect 165718 66019 165770 66071
rect 199030 66019 199082 66071
rect 171478 65945 171530 65997
rect 198838 65945 198890 65997
rect 174358 65871 174410 65923
rect 198742 65871 198794 65923
rect 177238 65797 177290 65849
rect 198934 65797 198986 65849
rect 152662 65353 152714 65405
rect 155158 65353 155210 65405
rect 146902 64095 146954 64147
rect 160438 64095 160490 64147
rect 143926 63355 143978 63407
rect 164278 63355 164330 63407
rect 146998 63281 147050 63333
rect 199126 63281 199178 63333
rect 151126 63207 151178 63259
rect 199030 63207 199082 63259
rect 155542 63133 155594 63185
rect 198934 63133 198986 63185
rect 160054 63059 160106 63111
rect 198838 63059 198890 63111
rect 163606 62985 163658 63037
rect 198742 62985 198794 63037
rect 202006 61505 202058 61557
rect 203062 61505 203114 61557
rect 202294 61431 202346 61483
rect 202966 61431 203018 61483
rect 202198 61357 202250 61409
rect 203350 61357 203402 61409
rect 202486 61283 202538 61335
rect 203254 61283 203306 61335
rect 203254 60839 203306 60891
rect 203734 60839 203786 60891
rect 146902 60617 146954 60669
rect 160534 60617 160586 60669
rect 146998 60543 147050 60595
rect 138166 60469 138218 60521
rect 159094 60469 159146 60521
rect 198934 60395 198986 60447
rect 640150 60395 640202 60447
rect 663574 60395 663626 60447
rect 164278 60321 164330 60373
rect 198838 60321 198890 60373
rect 167062 60247 167114 60299
rect 198742 60247 198794 60299
rect 204022 59063 204074 59115
rect 204982 59063 205034 59115
rect 204790 58915 204842 58967
rect 204982 58915 205034 58967
rect 204118 57287 204170 57339
rect 204502 57287 204554 57339
rect 204214 56251 204266 56303
rect 204694 56251 204746 56303
rect 204982 54771 205034 54823
rect 639574 54623 639626 54675
rect 639958 54623 640010 54675
rect 205942 54179 205994 54231
rect 201046 54105 201098 54157
rect 215158 54179 215210 54231
rect 632278 54179 632330 54231
rect 634966 54179 635018 54231
rect 206326 54105 206378 54157
rect 214966 54105 215018 54157
rect 633718 54105 633770 54157
rect 636214 54105 636266 54157
rect 200662 54031 200714 54083
rect 214774 54031 214826 54083
rect 633334 54031 633386 54083
rect 636022 54031 636074 54083
rect 201142 53957 201194 54009
rect 204982 53883 205034 53935
rect 206134 53883 206186 53935
rect 199702 53809 199754 53861
rect 206326 53809 206378 53861
rect 632566 53957 632618 54009
rect 635830 53957 635882 54009
rect 631894 53883 631946 53935
rect 635446 53883 635498 53935
rect 201430 53735 201482 53787
rect 201238 53661 201290 53713
rect 629302 53809 629354 53861
rect 634774 53809 634826 53861
rect 630358 53735 630410 53787
rect 635254 53735 635306 53787
rect 630070 53661 630122 53713
rect 635158 53661 635210 53713
rect 204310 53587 204362 53639
rect 207478 53587 207530 53639
rect 207574 53587 207626 53639
rect 209734 53587 209786 53639
rect 210742 53587 210794 53639
rect 211558 53587 211610 53639
rect 211942 53587 211994 53639
rect 213430 53587 213482 53639
rect 214150 53587 214202 53639
rect 214774 53587 214826 53639
rect 215638 53587 215690 53639
rect 631510 53587 631562 53639
rect 635638 53587 635690 53639
rect 199798 53513 199850 53565
rect 210070 53513 210122 53565
rect 631126 53513 631178 53565
rect 635926 53513 635978 53565
rect 163510 53439 163562 53491
rect 212854 53439 212906 53491
rect 627766 53439 627818 53491
rect 635734 53439 635786 53491
rect 202102 53365 202154 53417
rect 204310 53365 204362 53417
rect 204502 53365 204554 53417
rect 206326 53365 206378 53417
rect 206518 53365 206570 53417
rect 211222 53365 211274 53417
rect 160438 53291 160490 53343
rect 210262 53291 210314 53343
rect 204118 53217 204170 53269
rect 204502 53217 204554 53269
rect 204598 53217 204650 53269
rect 205558 53217 205610 53269
rect 206902 53217 206954 53269
rect 215830 53217 215882 53269
rect 160342 53143 160394 53195
rect 210646 53143 210698 53195
rect 204406 53069 204458 53121
rect 205270 53069 205322 53121
rect 205846 53069 205898 53121
rect 227926 53069 227978 53121
rect 160246 52995 160298 53047
rect 211030 52995 211082 53047
rect 163414 52921 163466 52973
rect 213238 52921 213290 52973
rect 160150 52847 160202 52899
rect 211702 52847 211754 52899
rect 163318 52773 163370 52825
rect 213910 52773 213962 52825
rect 159958 52699 160010 52751
rect 212086 52699 212138 52751
rect 160534 52625 160586 52677
rect 209878 52625 209930 52677
rect 159958 52551 160010 52603
rect 211414 52551 211466 52603
rect 162646 52477 162698 52529
rect 213622 52477 213674 52529
rect 162934 52403 162986 52455
rect 222550 52403 222602 52455
rect 163222 52329 163274 52381
rect 218710 52329 218762 52381
rect 162838 52255 162890 52307
rect 223510 52255 223562 52307
rect 163126 52181 163178 52233
rect 221302 52181 221354 52233
rect 162742 52107 162794 52159
rect 224278 52107 224330 52159
rect 204694 52033 204746 52085
rect 205174 52033 205226 52085
rect 205366 52033 205418 52085
rect 634102 52033 634154 52085
rect 159958 51959 160010 52011
rect 212470 51959 212522 52011
rect 212662 51959 212714 52011
rect 639766 51959 639818 52011
rect 204790 51885 204842 51937
rect 205078 51885 205130 51937
rect 206038 51885 206090 51937
rect 639670 51885 639722 51937
rect 205942 51811 205994 51863
rect 210838 51811 210890 51863
rect 204502 51663 204554 51715
rect 212278 51663 212330 51715
rect 204598 51589 204650 51641
rect 213046 51589 213098 51641
rect 202966 51515 203018 51567
rect 215254 51515 215306 51567
rect 145558 51367 145610 51419
rect 238006 51367 238058 51419
rect 145750 51293 145802 51345
rect 237142 51293 237194 51345
rect 143926 51219 143978 51271
rect 145558 51219 145610 51271
rect 145846 51219 145898 51271
rect 236374 51219 236426 51271
rect 146422 51145 146474 51197
rect 237526 51145 237578 51197
rect 144406 51071 144458 51123
rect 234550 51071 234602 51123
rect 144598 50997 144650 51049
rect 234166 50997 234218 51049
rect 144790 50923 144842 50975
rect 234934 50923 234986 50975
rect 145942 50849 145994 50901
rect 235798 50849 235850 50901
rect 146038 50775 146090 50827
rect 235318 50775 235370 50827
rect 145174 50701 145226 50753
rect 230902 50701 230954 50753
rect 145270 50627 145322 50679
rect 232726 50627 232778 50679
rect 146518 50553 146570 50605
rect 232342 50553 232394 50605
rect 146614 50479 146666 50531
rect 230998 50479 231050 50531
rect 146710 50405 146762 50457
rect 233110 50405 233162 50457
rect 146806 50331 146858 50383
rect 231382 50331 231434 50383
rect 145558 50257 145610 50309
rect 227542 50257 227594 50309
rect 144694 50183 144746 50235
rect 228790 50183 228842 50235
rect 144886 50109 144938 50161
rect 228694 50109 228746 50161
rect 144982 50035 145034 50087
rect 229174 50035 229226 50087
rect 145078 49961 145130 50013
rect 230134 49961 230186 50013
rect 144118 49887 144170 49939
rect 226966 49887 227018 49939
rect 144022 49813 144074 49865
rect 226102 49813 226154 49865
rect 144310 49739 144362 49791
rect 225718 49739 225770 49791
rect 146134 49665 146186 49717
rect 241942 49665 241994 49717
rect 145366 49591 145418 49643
rect 239734 49591 239786 49643
rect 144502 49517 144554 49569
rect 226486 49517 226538 49569
rect 146230 49443 146282 49495
rect 241174 49443 241226 49495
rect 145462 49295 145514 49347
rect 238966 49295 239018 49347
rect 146326 49221 146378 49273
rect 240790 49221 240842 49273
rect 145654 49147 145706 49199
rect 237622 49147 237674 49199
rect 202582 48925 202634 48977
rect 214294 48925 214346 48977
rect 216310 48925 216362 48977
rect 264886 48925 264938 48977
rect 627190 48925 627242 48977
rect 636118 48925 636170 48977
rect 202678 48851 202730 48903
rect 215062 48851 215114 48903
rect 215158 48851 215210 48903
rect 226582 48851 226634 48903
rect 202774 48777 202826 48829
rect 215446 48777 215498 48829
rect 204694 48629 204746 48681
rect 208918 48629 208970 48681
rect 204502 48555 204554 48607
rect 217654 48555 217706 48607
rect 203830 48481 203882 48533
rect 216886 48481 216938 48533
rect 203734 48407 203786 48459
rect 209302 48407 209354 48459
rect 235414 48407 235466 48459
rect 217270 48333 217322 48385
rect 628918 48259 628970 48311
rect 663382 48259 663434 48311
rect 147670 48185 147722 48237
rect 201622 48185 201674 48237
rect 203446 48185 203498 48237
rect 211606 48185 211658 48237
rect 147574 48111 147626 48163
rect 216118 48185 216170 48237
rect 216022 48111 216074 48163
rect 639382 48111 639434 48163
rect 202390 48037 202442 48089
rect 216502 48037 216554 48089
rect 216598 48037 216650 48089
rect 224758 48037 224810 48089
rect 148150 47963 148202 48015
rect 230518 47963 230570 48015
rect 203350 47889 203402 47941
rect 203254 47815 203306 47867
rect 208726 47815 208778 47867
rect 208918 47889 208970 47941
rect 221686 47889 221738 47941
rect 211606 47815 211658 47867
rect 219094 47815 219146 47867
rect 219478 47741 219530 47793
rect 148534 47667 148586 47719
rect 231958 47667 232010 47719
rect 627958 47667 628010 47719
rect 663190 47667 663242 47719
rect 148918 47593 148970 47645
rect 229750 47593 229802 47645
rect 208726 47519 208778 47571
rect 219862 47519 219914 47571
rect 201622 47445 201674 47497
rect 208342 47445 208394 47497
rect 148342 47371 148394 47423
rect 209302 47371 209354 47423
rect 209398 47371 209450 47423
rect 233590 47371 233642 47423
rect 149494 46779 149546 46831
rect 209398 46779 209450 46831
rect 149686 46705 149738 46757
rect 217846 46853 217898 46905
rect 639958 46853 640010 46905
rect 233302 46779 233354 46831
rect 209686 46705 209738 46757
rect 215158 46705 215210 46757
rect 215254 46705 215306 46757
rect 223126 46705 223178 46757
rect 149302 46631 149354 46683
rect 161302 46631 161354 46683
rect 181366 46631 181418 46683
rect 221782 46631 221834 46683
rect 202486 46557 202538 46609
rect 147862 46483 147914 46535
rect 202294 46409 202346 46461
rect 147958 46335 148010 46387
rect 207862 46335 207914 46387
rect 202006 46261 202058 46313
rect 207958 46261 208010 46313
rect 208534 46557 208586 46609
rect 216598 46557 216650 46609
rect 216694 46557 216746 46609
rect 639862 46557 639914 46609
rect 208342 46483 208394 46535
rect 220918 46483 220970 46535
rect 221782 46483 221834 46535
rect 228310 46483 228362 46535
rect 222166 46409 222218 46461
rect 224662 46335 224714 46387
rect 225334 46261 225386 46313
rect 147766 46187 147818 46239
rect 223894 46187 223946 46239
rect 202198 46113 202250 46165
rect 222070 46113 222122 46165
rect 205174 45151 205226 45203
rect 403126 45151 403178 45203
rect 206998 45077 207050 45129
rect 408886 45077 408938 45129
rect 207382 45003 207434 45055
rect 406294 45003 406346 45055
rect 208054 44929 208106 44981
rect 446518 44929 446570 44981
rect 209206 44855 209258 44907
rect 499990 44855 500042 44907
rect 205270 44781 205322 44833
rect 508246 44781 508298 44833
rect 209590 44707 209642 44759
rect 523894 44707 523946 44759
rect 205558 44633 205610 44685
rect 521206 44633 521258 44685
rect 613462 44633 613514 44685
rect 635542 44633 635594 44685
rect 508246 43227 508298 43279
rect 520342 43153 520394 43205
rect 206614 42339 206666 42391
rect 310102 42339 310154 42391
rect 201334 42117 201386 42169
rect 405238 42117 405290 42169
rect 207670 42043 207722 42095
rect 460054 42043 460106 42095
rect 459190 41969 459242 42021
rect 463702 41969 463754 42021
rect 403126 41895 403178 41947
rect 514870 41747 514922 41799
rect 208438 41673 208490 41725
rect 499990 40341 500042 40393
rect 512566 40267 512618 40319
rect 446518 37381 446570 37433
rect 459190 37381 459242 37433
<< metal2 >>
rect 447766 1005723 447818 1005729
rect 447766 1005665 447818 1005671
rect 95062 1005575 95114 1005581
rect 95062 1005517 95114 1005523
rect 437206 1005575 437258 1005581
rect 437206 1005517 437258 1005523
rect 93622 1005501 93674 1005507
rect 93622 1005443 93674 1005449
rect 92566 1005353 92618 1005359
rect 92566 1005295 92618 1005301
rect 92374 1005279 92426 1005285
rect 92374 1005221 92426 1005227
rect 61846 999433 61898 999439
rect 61846 999375 61898 999381
rect 74710 999433 74762 999439
rect 74710 999375 74762 999381
rect 45142 985521 45194 985527
rect 45142 985463 45194 985469
rect 45046 985225 45098 985231
rect 45046 985167 45098 985173
rect 44950 985151 45002 985157
rect 44950 985093 45002 985099
rect 44854 985077 44906 985083
rect 44854 985019 44906 985025
rect 42550 985003 42602 985009
rect 42550 984945 42602 984951
rect 41794 968771 41822 969252
rect 41780 968762 41836 968771
rect 41780 968697 41836 968706
rect 41794 967143 41822 967402
rect 42562 967323 42590 984945
rect 44758 983819 44810 983825
rect 44758 983761 44810 983767
rect 44566 983745 44618 983751
rect 44566 983687 44618 983693
rect 42166 967317 42218 967323
rect 42166 967259 42218 967265
rect 42550 967317 42602 967323
rect 42550 967259 42602 967265
rect 41780 967134 41836 967143
rect 41780 967069 41836 967078
rect 42178 966736 42206 967259
rect 41794 965071 41822 965552
rect 41780 965062 41836 965071
rect 41780 964997 41836 965006
rect 41794 964035 41822 964368
rect 41780 964026 41836 964035
rect 41780 963961 41836 963970
rect 41794 963443 41822 963702
rect 41780 963434 41836 963443
rect 41780 963369 41836 963378
rect 41794 962851 41822 963081
rect 41780 962842 41836 962851
rect 41780 962777 41836 962786
rect 41890 962259 41918 962518
rect 41876 962250 41932 962259
rect 41876 962185 41932 962194
rect 42356 962250 42412 962259
rect 42356 962185 42412 962194
rect 42068 961806 42124 961815
rect 42068 961741 42124 961750
rect 42082 961260 42110 961741
rect 42370 961033 42398 962185
rect 42166 961027 42218 961033
rect 42166 960969 42218 960975
rect 42358 961027 42410 961033
rect 42358 960969 42410 960975
rect 42178 960594 42206 960969
rect 41794 959743 41822 960045
rect 41780 959734 41836 959743
rect 41780 959669 41836 959678
rect 41890 959151 41918 959410
rect 41876 959142 41932 959151
rect 41876 959077 41932 959086
rect 42082 958411 42110 958744
rect 42068 958402 42124 958411
rect 42068 958337 42124 958346
rect 42178 957819 42206 958226
rect 42164 957810 42220 957819
rect 42164 957745 42220 957754
rect 42178 956191 42206 956376
rect 42358 956217 42410 956223
rect 42164 956182 42220 956191
rect 42358 956159 42410 956165
rect 42164 956117 42220 956126
rect 42082 955261 42110 955710
rect 42070 955255 42122 955261
rect 42070 955197 42122 955203
rect 42178 954669 42206 955077
rect 42166 954663 42218 954669
rect 42166 954605 42218 954611
rect 42262 907525 42314 907531
rect 42260 907490 42262 907499
rect 42314 907490 42316 907499
rect 42260 907425 42316 907434
rect 42370 906759 42398 956159
rect 42934 955255 42986 955261
rect 42934 955197 42986 955203
rect 42646 908117 42698 908123
rect 42644 908082 42646 908091
rect 42698 908082 42700 908091
rect 42644 908017 42700 908026
rect 42356 906750 42412 906759
rect 42356 906685 42412 906694
rect 40340 905418 40396 905427
rect 40340 905353 40396 905362
rect 40052 901422 40108 901431
rect 40052 901357 40108 901366
rect 40066 872677 40094 901357
rect 40054 872671 40106 872677
rect 40054 872613 40106 872619
rect 39958 869859 40010 869865
rect 39958 869801 40010 869807
rect 39970 852549 39998 869801
rect 39958 852543 40010 852549
rect 39958 852485 40010 852491
rect 40054 852395 40106 852401
rect 40054 852337 40106 852343
rect 40066 846703 40094 852337
rect 40054 846697 40106 846703
rect 40054 846639 40106 846645
rect 40150 846697 40202 846703
rect 40150 846639 40202 846645
rect 40162 842675 40190 846639
rect 40148 842666 40204 842675
rect 40148 842601 40204 842610
rect 39956 827570 40012 827579
rect 39956 827505 40012 827514
rect 39970 826649 39998 827505
rect 39958 826643 40010 826649
rect 39958 826585 40010 826591
rect 40150 826643 40202 826649
rect 40150 826585 40202 826591
rect 40162 819439 40190 826585
rect 40354 820771 40382 905353
rect 42646 904861 42698 904867
rect 42644 904826 42646 904835
rect 42698 904826 42700 904835
rect 42644 904761 42700 904770
rect 42946 897731 42974 955197
rect 43030 954663 43082 954669
rect 43030 954605 43082 954611
rect 43042 901135 43070 954605
rect 43124 907194 43180 907203
rect 43124 907129 43180 907138
rect 43028 901126 43084 901135
rect 43028 901061 43084 901070
rect 42932 897722 42988 897731
rect 42932 897657 42988 897666
rect 42356 891210 42412 891219
rect 42356 891145 42412 891154
rect 42370 889739 42398 891145
rect 42356 889730 42412 889739
rect 42356 889665 42358 889674
rect 42410 889665 42412 889674
rect 42358 889633 42410 889639
rect 43138 887371 43166 907129
rect 43220 904234 43276 904243
rect 43220 904169 43276 904178
rect 43234 901579 43262 904169
rect 44578 903355 44606 983687
rect 44662 983671 44714 983677
rect 44662 983613 44714 983619
rect 44674 904867 44702 983613
rect 44662 904861 44714 904867
rect 44662 904803 44714 904809
rect 44770 904243 44798 983761
rect 44756 904234 44812 904243
rect 44756 904169 44812 904178
rect 44564 903346 44620 903355
rect 44564 903281 44620 903290
rect 43220 901570 43276 901579
rect 43220 901505 43276 901514
rect 44566 889691 44618 889697
rect 44566 889633 44618 889639
rect 43124 887362 43180 887371
rect 43124 887297 43180 887306
rect 40438 872671 40490 872677
rect 40438 872613 40490 872619
rect 40450 869865 40478 872613
rect 40438 869859 40490 869865
rect 40438 869801 40490 869807
rect 40820 852730 40876 852739
rect 40820 852665 40876 852674
rect 40340 820762 40396 820771
rect 40340 820697 40396 820706
rect 40834 819587 40862 852665
rect 42358 823905 42410 823911
rect 42356 823870 42358 823879
rect 42410 823870 42412 823879
rect 42356 823805 42412 823814
rect 42452 822686 42508 822695
rect 42452 822621 42508 822630
rect 42358 822277 42410 822283
rect 42356 822242 42358 822251
rect 42410 822242 42412 822251
rect 42356 822177 42412 822186
rect 42466 821913 42494 822621
rect 42454 821907 42506 821913
rect 42454 821849 42506 821855
rect 43220 821206 43276 821215
rect 43220 821141 43276 821150
rect 40820 819578 40876 819587
rect 40820 819513 40876 819522
rect 40148 819430 40204 819439
rect 40148 819365 40204 819374
rect 40162 817917 40190 819365
rect 42356 817950 42412 817959
rect 40150 817911 40202 817917
rect 42356 817885 42412 817894
rect 40150 817853 40202 817859
rect 40244 816766 40300 816775
rect 40244 816701 40300 816710
rect 37268 815878 37324 815887
rect 37268 815813 37324 815822
rect 37282 802123 37310 815813
rect 37364 812770 37420 812779
rect 37364 812705 37420 812714
rect 37268 802114 37324 802123
rect 37268 802049 37324 802058
rect 37378 801975 37406 812705
rect 40258 803487 40286 816701
rect 41972 814398 42028 814407
rect 41972 814333 42028 814342
rect 41876 813658 41932 813667
rect 41876 813593 41932 813602
rect 41684 811142 41740 811151
rect 41684 811077 41740 811086
rect 40246 803481 40298 803487
rect 40246 803423 40298 803429
rect 37364 801966 37420 801975
rect 37364 801901 37420 801910
rect 41698 800495 41726 811077
rect 41780 809662 41836 809671
rect 41780 809597 41836 809606
rect 41684 800486 41740 800495
rect 41684 800421 41740 800430
rect 41794 800347 41822 809597
rect 41780 800338 41836 800347
rect 41780 800273 41836 800282
rect 41890 800231 41918 813593
rect 41986 802451 42014 814333
rect 42068 809218 42124 809227
rect 42068 809153 42124 809162
rect 41974 802445 42026 802451
rect 41974 802387 42026 802393
rect 42082 800347 42110 809153
rect 42164 808330 42220 808339
rect 42164 808265 42220 808274
rect 42068 800338 42124 800347
rect 42068 800273 42124 800282
rect 41878 800225 41930 800231
rect 41878 800167 41930 800173
rect 42178 800176 42206 808265
rect 42260 805222 42316 805231
rect 42260 805157 42262 805166
rect 42314 805157 42316 805166
rect 42262 805125 42314 805131
rect 42370 804468 42398 817885
rect 42452 815286 42508 815295
rect 42452 815221 42508 815230
rect 42274 804440 42398 804468
rect 42274 800305 42302 804440
rect 42466 803635 42494 815221
rect 43124 812326 43180 812335
rect 43124 812261 43180 812270
rect 43138 810536 43166 812261
rect 43042 810508 43166 810536
rect 42932 807294 42988 807303
rect 42932 807229 42988 807238
rect 42946 804172 42974 807229
rect 42754 804144 42974 804172
rect 42454 803629 42506 803635
rect 42454 803571 42506 803577
rect 42454 803481 42506 803487
rect 42454 803423 42506 803429
rect 42262 800299 42314 800305
rect 42262 800241 42314 800247
rect 42178 800148 42302 800176
rect 42274 800051 42302 800148
rect 42260 800042 42316 800051
rect 42260 799977 42316 799986
rect 41878 799781 41930 799787
rect 41878 799723 41930 799729
rect 41890 799422 41918 799723
rect 42466 798085 42494 803423
rect 42166 798079 42218 798085
rect 42166 798021 42218 798027
rect 42454 798079 42506 798085
rect 42454 798021 42506 798027
rect 42178 797605 42206 798021
rect 42452 797970 42508 797979
rect 42452 797905 42508 797914
rect 42070 797339 42122 797345
rect 42070 797281 42122 797287
rect 42082 796980 42110 797281
rect 42166 796303 42218 796309
rect 42166 796245 42218 796251
rect 42178 795765 42206 796245
rect 42166 795045 42218 795051
rect 42166 794987 42218 794993
rect 42178 794569 42206 794987
rect 41780 794270 41836 794279
rect 41780 794205 41836 794214
rect 41794 793946 41822 794205
rect 42466 793867 42494 797905
rect 42754 795051 42782 804144
rect 43042 803876 43070 810508
rect 43124 810402 43180 810411
rect 43124 810337 43180 810346
rect 42850 803848 43070 803876
rect 42742 795045 42794 795051
rect 42742 794987 42794 794993
rect 42740 794862 42796 794871
rect 42740 794797 42796 794806
rect 42166 793861 42218 793867
rect 42166 793803 42218 793809
rect 42454 793861 42506 793867
rect 42454 793803 42506 793809
rect 42178 793280 42206 793803
rect 42166 793195 42218 793201
rect 42166 793137 42218 793143
rect 42178 792729 42206 793137
rect 42260 792198 42316 792207
rect 42260 792133 42316 792142
rect 41794 791171 41822 791430
rect 41780 791162 41836 791171
rect 41780 791097 41836 791106
rect 42164 791014 42220 791023
rect 42164 790949 42220 790958
rect 42178 790797 42206 790949
rect 42274 790260 42302 792133
rect 42754 792059 42782 794797
rect 42740 792050 42796 792059
rect 42740 791985 42796 791994
rect 42452 791902 42508 791911
rect 42452 791837 42508 791846
rect 42192 790232 42302 790260
rect 42262 790087 42314 790093
rect 42262 790029 42314 790035
rect 42166 789939 42218 789945
rect 42166 789881 42218 789887
rect 42178 789580 42206 789881
rect 42274 788971 42302 790029
rect 42192 788943 42302 788971
rect 42262 788903 42314 788909
rect 42262 788845 42314 788851
rect 42274 788410 42302 788845
rect 42192 788382 42302 788410
rect 42166 787053 42218 787059
rect 42166 786995 42218 787001
rect 42178 786546 42206 786995
rect 42466 786467 42494 791837
rect 42740 791754 42796 791763
rect 42740 791689 42796 791698
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42454 786461 42506 786467
rect 42454 786403 42506 786409
rect 42178 785921 42206 786403
rect 42754 785653 42782 791689
rect 42850 790093 42878 803848
rect 42934 803629 42986 803635
rect 42934 803571 42986 803577
rect 42838 790087 42890 790093
rect 42838 790029 42890 790035
rect 42946 788909 42974 803571
rect 43030 802445 43082 802451
rect 43030 802387 43082 802393
rect 43042 793201 43070 802387
rect 43138 796309 43166 810337
rect 43126 796303 43178 796309
rect 43126 796245 43178 796251
rect 43126 796155 43178 796161
rect 43126 796097 43178 796103
rect 43030 793195 43082 793201
rect 43030 793137 43082 793143
rect 43138 792165 43166 796097
rect 43126 792159 43178 792165
rect 43126 792101 43178 792107
rect 43124 792050 43180 792059
rect 43030 792011 43082 792017
rect 43124 791985 43180 791994
rect 43030 791953 43082 791959
rect 42934 788903 42986 788909
rect 42934 788845 42986 788851
rect 43042 787059 43070 791953
rect 43138 789945 43166 791985
rect 43126 789939 43178 789945
rect 43126 789881 43178 789887
rect 43030 787053 43082 787059
rect 43030 786995 43082 787001
rect 42070 785647 42122 785653
rect 42070 785589 42122 785595
rect 42742 785647 42794 785653
rect 42742 785589 42794 785595
rect 42082 785288 42110 785589
rect 42740 780506 42796 780515
rect 42740 780441 42742 780450
rect 42794 780441 42796 780450
rect 42742 780409 42794 780415
rect 42454 779949 42506 779955
rect 42452 779914 42454 779923
rect 42506 779914 42508 779923
rect 42452 779849 42508 779858
rect 42742 778913 42794 778919
rect 42740 778878 42742 778887
rect 42794 778878 42796 778887
rect 42740 778813 42796 778822
rect 43234 777259 43262 821141
rect 43318 817911 43370 817917
rect 43318 817853 43370 817859
rect 43220 777250 43276 777259
rect 43220 777185 43276 777194
rect 43220 776510 43276 776519
rect 43330 776496 43358 817853
rect 43510 800891 43562 800897
rect 43510 800833 43562 800839
rect 43414 800299 43466 800305
rect 43414 800241 43466 800247
rect 43426 796161 43454 800241
rect 43522 797345 43550 800833
rect 43510 797339 43562 797345
rect 43510 797281 43562 797287
rect 43414 796155 43466 796161
rect 43414 796097 43466 796103
rect 43606 792159 43658 792165
rect 43606 792101 43658 792107
rect 43618 792017 43646 792101
rect 43606 792011 43658 792017
rect 43606 791953 43658 791959
rect 43412 777990 43468 777999
rect 43412 777925 43468 777934
rect 43276 776468 43358 776496
rect 43220 776445 43276 776454
rect 42836 774882 42892 774891
rect 42836 774817 42892 774826
rect 38804 773550 38860 773559
rect 38804 773485 38860 773494
rect 35924 772662 35980 772671
rect 35924 772597 35980 772606
rect 35938 760239 35966 772597
rect 37364 769554 37420 769563
rect 37364 769489 37420 769498
rect 35924 760230 35980 760239
rect 35924 760165 35980 760174
rect 37378 759647 37406 769489
rect 37364 759638 37420 759647
rect 37364 759573 37420 759582
rect 38818 758611 38846 773485
rect 41972 771182 42028 771191
rect 41972 771117 42028 771126
rect 41780 770442 41836 770451
rect 41780 770377 41836 770386
rect 38804 758602 38860 758611
rect 38804 758537 38860 758546
rect 41794 757015 41822 770377
rect 41876 767926 41932 767935
rect 41876 767861 41932 767870
rect 41890 757089 41918 767861
rect 41986 757163 42014 771117
rect 42452 769110 42508 769119
rect 42452 769045 42508 769054
rect 42164 766002 42220 766011
rect 42164 765937 42220 765946
rect 42068 765262 42124 765271
rect 42068 765197 42124 765206
rect 41974 757157 42026 757163
rect 41974 757099 42026 757105
rect 41878 757083 41930 757089
rect 41878 757025 41930 757031
rect 42082 757015 42110 765197
rect 42178 757131 42206 765937
rect 42466 757311 42494 769045
rect 42740 764596 42796 764605
rect 42740 764531 42796 764540
rect 42454 757305 42506 757311
rect 42454 757247 42506 757253
rect 42164 757122 42220 757131
rect 42164 757057 42220 757066
rect 41782 757009 41834 757015
rect 41782 756951 41834 756957
rect 42070 757009 42122 757015
rect 42070 756951 42122 756957
rect 41782 756787 41834 756793
rect 41782 756729 41834 756735
rect 41794 756245 41822 756729
rect 41876 754902 41932 754911
rect 41876 754837 41932 754846
rect 41890 754430 41918 754837
rect 42452 754310 42508 754319
rect 42452 754245 42508 754254
rect 42166 754123 42218 754129
rect 42166 754065 42218 754071
rect 42178 753764 42206 754065
rect 42070 753087 42122 753093
rect 42070 753029 42122 753035
rect 42082 752580 42110 753029
rect 42070 751829 42122 751835
rect 42070 751771 42122 751777
rect 42082 751396 42110 751771
rect 42070 751163 42122 751169
rect 42070 751105 42122 751111
rect 42082 750730 42110 751105
rect 42166 750423 42218 750429
rect 42166 750365 42218 750371
rect 42178 750064 42206 750365
rect 42070 749979 42122 749985
rect 42070 749921 42122 749927
rect 42082 749546 42110 749921
rect 42262 748943 42314 748949
rect 42262 748885 42314 748891
rect 41780 748686 41836 748695
rect 41780 748621 41836 748630
rect 41794 748214 41822 748621
rect 41986 747363 42014 747622
rect 42166 747463 42218 747469
rect 42166 747405 42218 747411
rect 41972 747354 42028 747363
rect 41972 747289 42028 747298
rect 42178 747030 42206 747405
rect 42274 746415 42302 748885
rect 42466 747469 42494 754245
rect 42754 751835 42782 764531
rect 42850 751951 42878 774817
rect 42932 772514 42988 772523
rect 42932 772449 42988 772458
rect 42946 767172 42974 772449
rect 43124 767778 43180 767787
rect 43124 767713 43180 767722
rect 42946 767144 43070 767172
rect 42932 767038 42988 767047
rect 42932 766973 42988 766982
rect 42946 758125 42974 766973
rect 42934 758119 42986 758125
rect 42934 758061 42986 758067
rect 42934 757971 42986 757977
rect 42934 757913 42986 757919
rect 42946 754129 42974 757913
rect 42934 754123 42986 754129
rect 42934 754065 42986 754071
rect 42934 753975 42986 753981
rect 42934 753917 42986 753923
rect 42836 751942 42892 751951
rect 42946 751909 42974 753917
rect 42836 751877 42892 751886
rect 42934 751903 42986 751909
rect 42934 751845 42986 751851
rect 42742 751829 42794 751835
rect 42742 751771 42794 751777
rect 42838 751829 42890 751835
rect 42838 751771 42890 751777
rect 42740 751646 42796 751655
rect 42740 751581 42796 751590
rect 42454 747463 42506 747469
rect 42454 747405 42506 747411
rect 42192 746387 42302 746415
rect 42070 746131 42122 746137
rect 42070 746073 42122 746079
rect 42082 745772 42110 746073
rect 42166 745687 42218 745693
rect 42166 745629 42218 745635
rect 42178 745180 42206 745629
rect 42754 743843 42782 751581
rect 42850 751169 42878 751771
rect 42934 751755 42986 751761
rect 42934 751697 42986 751703
rect 42838 751163 42890 751169
rect 42838 751105 42890 751111
rect 42838 751015 42890 751021
rect 42838 750957 42890 750963
rect 42850 748949 42878 750957
rect 42946 749985 42974 751697
rect 42934 749979 42986 749985
rect 42934 749921 42986 749927
rect 42838 748943 42890 748949
rect 42838 748885 42890 748891
rect 42836 747206 42892 747215
rect 42836 747141 42892 747150
rect 42166 743837 42218 743843
rect 42166 743779 42218 743785
rect 42742 743837 42794 743843
rect 42742 743779 42794 743785
rect 42178 743365 42206 743779
rect 42850 743103 42878 747141
rect 42932 746910 42988 746919
rect 42932 746845 42988 746854
rect 42070 743097 42122 743103
rect 42070 743039 42122 743045
rect 42838 743097 42890 743103
rect 42838 743039 42890 743045
rect 42082 742738 42110 743039
rect 42946 742437 42974 746845
rect 43042 745693 43070 767144
rect 43138 753093 43166 767713
rect 43234 761867 43262 776445
rect 43220 761858 43276 761867
rect 43220 761793 43276 761802
rect 43222 758119 43274 758125
rect 43222 758061 43274 758067
rect 43234 753981 43262 758061
rect 43318 757009 43370 757015
rect 43318 756951 43370 756957
rect 43222 753975 43274 753981
rect 43222 753917 43274 753923
rect 43330 753112 43358 756951
rect 43126 753087 43178 753093
rect 43126 753029 43178 753035
rect 43234 753084 43358 753112
rect 43234 752964 43262 753084
rect 43138 752936 43262 752964
rect 43138 750429 43166 752936
rect 43126 750423 43178 750429
rect 43126 750365 43178 750371
rect 43126 750275 43178 750281
rect 43126 750217 43178 750223
rect 43138 746137 43166 750217
rect 43126 746131 43178 746137
rect 43126 746073 43178 746079
rect 43030 745687 43082 745693
rect 43030 745629 43082 745635
rect 42166 742431 42218 742437
rect 42166 742373 42218 742379
rect 42934 742431 42986 742437
rect 42934 742373 42986 742379
rect 42178 742072 42206 742373
rect 42644 737290 42700 737299
rect 42644 737225 42646 737234
rect 42698 737225 42700 737234
rect 42646 737193 42698 737199
rect 42358 736733 42410 736739
rect 42356 736698 42358 736707
rect 42410 736698 42412 736707
rect 42356 736633 42412 736642
rect 42356 735514 42412 735523
rect 42356 735449 42358 735458
rect 42410 735449 42412 735458
rect 42358 735417 42410 735423
rect 43220 734922 43276 734931
rect 43220 734857 43276 734866
rect 42932 731666 42988 731675
rect 42932 731601 42988 731610
rect 40244 730334 40300 730343
rect 40244 730269 40300 730278
rect 40258 715057 40286 730269
rect 41588 728854 41644 728863
rect 41588 728789 41644 728798
rect 41492 727226 41548 727235
rect 41492 727161 41548 727170
rect 40246 715051 40298 715057
rect 40246 714993 40298 714999
rect 41506 714095 41534 727161
rect 41602 714169 41630 728789
rect 41780 727966 41836 727975
rect 41780 727901 41836 727910
rect 41684 725894 41740 725903
rect 41684 725829 41740 725838
rect 41590 714163 41642 714169
rect 41590 714105 41642 714111
rect 41698 714095 41726 725829
rect 41794 716135 41822 727901
rect 42068 724710 42124 724719
rect 42068 724645 42124 724654
rect 41972 723230 42028 723239
rect 41972 723165 42028 723174
rect 41780 716126 41836 716135
rect 41780 716061 41836 716070
rect 41878 715051 41930 715057
rect 41878 714993 41930 714999
rect 41494 714089 41546 714095
rect 41494 714031 41546 714037
rect 41686 714089 41738 714095
rect 41890 714063 41918 714993
rect 41686 714031 41738 714037
rect 41876 714054 41932 714063
rect 41876 713989 41932 713998
rect 41986 713873 42014 723165
rect 42082 713915 42110 724645
rect 42164 724118 42220 724127
rect 42164 724053 42220 724062
rect 42178 717888 42206 724053
rect 42260 719974 42316 719983
rect 42260 719909 42316 719918
rect 42274 718799 42302 719909
rect 42260 718790 42316 718799
rect 42260 718725 42262 718734
rect 42314 718725 42316 718734
rect 42262 718693 42314 718699
rect 42178 717860 42398 717888
rect 42068 713906 42124 713915
rect 41974 713867 42026 713873
rect 42068 713841 42124 713850
rect 41974 713809 42026 713815
rect 41782 713571 41834 713577
rect 41782 713513 41834 713519
rect 41794 713064 41822 713513
rect 42068 711686 42124 711695
rect 42068 711621 42124 711630
rect 42082 711214 42110 711621
rect 42166 710907 42218 710913
rect 42166 710849 42218 710855
rect 42178 710548 42206 710849
rect 42370 709951 42398 717860
rect 42946 711843 42974 731601
rect 43028 723082 43084 723091
rect 43028 723017 43084 723026
rect 42932 711834 42988 711843
rect 42932 711769 42988 711778
rect 43042 711695 43070 723017
rect 43126 717123 43178 717129
rect 43126 717065 43178 717071
rect 43028 711686 43084 711695
rect 43028 711621 43084 711630
rect 43138 711505 43166 717065
rect 42934 711499 42986 711505
rect 42934 711441 42986 711447
rect 43126 711499 43178 711505
rect 43126 711441 43178 711447
rect 42946 711357 42974 711441
rect 42934 711351 42986 711357
rect 42934 711293 42986 711299
rect 43124 711242 43180 711251
rect 43124 711177 43180 711186
rect 42836 711094 42892 711103
rect 42836 711029 42892 711038
rect 42166 709945 42218 709951
rect 42166 709887 42218 709893
rect 42358 709945 42410 709951
rect 42358 709887 42410 709893
rect 42178 709364 42206 709887
rect 42068 708578 42124 708587
rect 42068 708513 42124 708522
rect 42082 708180 42110 708513
rect 42166 707947 42218 707953
rect 42166 707889 42218 707895
rect 42178 707514 42206 707889
rect 42164 707394 42220 707403
rect 42164 707329 42220 707338
rect 42178 706881 42206 707329
rect 41972 706506 42028 706515
rect 41972 706441 42028 706450
rect 42550 706467 42602 706473
rect 41986 706330 42014 706441
rect 42550 706409 42602 706415
rect 42262 705653 42314 705659
rect 42262 705595 42314 705601
rect 41794 704739 41822 705041
rect 41780 704730 41836 704739
rect 41780 704665 41836 704674
rect 42082 704147 42110 704406
rect 42068 704138 42124 704147
rect 42068 704073 42124 704082
rect 42274 703859 42302 705595
rect 42192 703831 42302 703859
rect 42070 703729 42122 703735
rect 42070 703671 42122 703677
rect 42260 703694 42316 703703
rect 42082 703222 42110 703671
rect 42260 703629 42316 703638
rect 42166 702915 42218 702921
rect 42166 702857 42218 702863
rect 42178 702556 42206 702857
rect 42166 702323 42218 702329
rect 42166 702265 42218 702271
rect 42178 702005 42206 702265
rect 42274 700891 42302 703629
rect 42562 702329 42590 706409
rect 42850 703735 42878 711029
rect 43028 707838 43084 707847
rect 43028 707773 43084 707782
rect 42934 707281 42986 707287
rect 42934 707223 42986 707229
rect 42838 703729 42890 703735
rect 42838 703671 42890 703677
rect 42836 703546 42892 703555
rect 42836 703481 42892 703490
rect 42550 702323 42602 702329
rect 42550 702265 42602 702271
rect 42260 700882 42316 700891
rect 42260 700817 42316 700826
rect 42070 700621 42122 700627
rect 42070 700563 42122 700569
rect 42260 700586 42316 700595
rect 42082 700188 42110 700563
rect 42260 700521 42316 700530
rect 42166 700103 42218 700109
rect 42166 700045 42218 700051
rect 42178 699522 42206 700045
rect 42274 699388 42302 700521
rect 42850 700109 42878 703481
rect 42946 702921 42974 707223
rect 42934 702915 42986 702921
rect 42934 702857 42986 702863
rect 43042 700627 43070 707773
rect 43138 705659 43166 711177
rect 43126 705653 43178 705659
rect 43126 705595 43178 705601
rect 43030 700621 43082 700627
rect 43030 700563 43082 700569
rect 42838 700103 42890 700109
rect 42838 700045 42890 700051
rect 42358 699881 42410 699887
rect 42358 699823 42410 699829
rect 42178 699360 42302 699388
rect 42178 698856 42206 699360
rect 42370 693491 42398 699823
rect 42644 694074 42700 694083
rect 42644 694009 42646 694018
rect 42698 694009 42700 694018
rect 42646 693977 42698 693983
rect 42356 693482 42412 693491
rect 42356 693417 42412 693426
rect 41396 692742 41452 692751
rect 41396 692677 41452 692686
rect 40244 687118 40300 687127
rect 40244 687053 40300 687062
rect 40258 672211 40286 687053
rect 41410 674843 41438 692677
rect 42646 692481 42698 692487
rect 42644 692446 42646 692455
rect 42698 692446 42700 692455
rect 42644 692381 42700 692390
rect 43234 690827 43262 734857
rect 43426 734043 43454 777925
rect 43510 757305 43562 757311
rect 43510 757247 43562 757253
rect 43522 750281 43550 757247
rect 43702 757157 43754 757163
rect 43702 757099 43754 757105
rect 43606 757083 43658 757089
rect 43606 757025 43658 757031
rect 43618 751021 43646 757025
rect 43714 751761 43742 757099
rect 43702 751755 43754 751761
rect 43702 751697 43754 751703
rect 43606 751015 43658 751021
rect 43606 750957 43658 750963
rect 43510 750275 43562 750281
rect 43510 750217 43562 750223
rect 43412 734034 43468 734043
rect 43412 733969 43468 733978
rect 43510 714163 43562 714169
rect 43510 714105 43562 714111
rect 43318 713867 43370 713873
rect 43318 713809 43370 713815
rect 43330 711579 43358 713809
rect 43318 711573 43370 711579
rect 43318 711515 43370 711521
rect 43414 711425 43466 711431
rect 43414 711367 43466 711373
rect 43426 710913 43454 711367
rect 43414 710907 43466 710913
rect 43414 710849 43466 710855
rect 43522 706473 43550 714105
rect 43606 714089 43658 714095
rect 43606 714031 43658 714037
rect 43618 707287 43646 714031
rect 43702 711277 43754 711283
rect 43702 711219 43754 711225
rect 43714 707953 43742 711219
rect 43702 707947 43754 707953
rect 43702 707889 43754 707895
rect 43606 707281 43658 707287
rect 43606 707223 43658 707229
rect 43510 706467 43562 706473
rect 43510 706409 43562 706415
rect 43412 691706 43468 691715
rect 43412 691641 43468 691650
rect 43220 690818 43276 690827
rect 43220 690753 43276 690762
rect 41588 688302 41644 688311
rect 41588 688237 41644 688246
rect 41396 674834 41452 674843
rect 41396 674769 41452 674778
rect 41602 674579 41630 688237
rect 41684 685638 41740 685647
rect 41684 685573 41740 685582
rect 41590 674573 41642 674579
rect 41590 674515 41642 674521
rect 40246 672205 40298 672211
rect 40246 672147 40298 672153
rect 41014 672205 41066 672211
rect 41014 672147 41066 672153
rect 41026 670995 41054 672147
rect 41698 672063 41726 685573
rect 41780 684010 41836 684019
rect 41780 683945 41836 683954
rect 41686 672057 41738 672063
rect 41686 671999 41738 672005
rect 41012 670986 41068 670995
rect 41012 670921 41068 670930
rect 41794 670657 41822 683945
rect 41876 681494 41932 681503
rect 41876 681429 41932 681438
rect 41890 670805 41918 681429
rect 41972 680902 42028 680911
rect 41972 680837 42028 680846
rect 41878 670799 41930 670805
rect 41878 670741 41930 670747
rect 41986 670657 42014 680837
rect 42260 680014 42316 680023
rect 42260 679949 42316 679958
rect 42274 671989 42302 679949
rect 43124 678238 43180 678247
rect 43124 678173 43180 678182
rect 42356 677202 42412 677211
rect 42356 677137 42412 677146
rect 42370 675731 42398 677137
rect 42356 675722 42412 675731
rect 42356 675657 42358 675666
rect 42410 675657 42412 675666
rect 42358 675625 42410 675631
rect 43138 674672 43166 678173
rect 43042 674644 43166 674672
rect 42646 672057 42698 672063
rect 42646 671999 42698 672005
rect 42262 671983 42314 671989
rect 42262 671925 42314 671931
rect 42454 671983 42506 671989
rect 42454 671925 42506 671931
rect 41782 670651 41834 670657
rect 41782 670593 41834 670599
rect 41974 670651 42026 670657
rect 41974 670593 42026 670599
rect 41782 670355 41834 670361
rect 41782 670297 41834 670303
rect 41794 669848 41822 670297
rect 42466 669251 42494 671925
rect 42658 670995 42686 671999
rect 43042 670995 43070 674644
rect 43126 674573 43178 674579
rect 43126 674515 43178 674521
rect 42644 670986 42700 670995
rect 42644 670921 42700 670930
rect 43028 670986 43084 670995
rect 43028 670921 43084 670930
rect 43138 670879 43166 674515
rect 43318 671391 43370 671397
rect 43318 671333 43370 671339
rect 43126 670873 43178 670879
rect 43126 670815 43178 670821
rect 43222 670799 43274 670805
rect 43222 670741 43274 670747
rect 42934 670651 42986 670657
rect 42934 670593 42986 670599
rect 42454 669245 42506 669251
rect 42454 669187 42506 669193
rect 42838 668949 42890 668955
rect 42548 668914 42604 668923
rect 42838 668891 42890 668897
rect 42548 668849 42604 668858
rect 41780 668470 41836 668479
rect 41780 668405 41836 668414
rect 41794 667998 41822 668405
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42178 667361 42206 667855
rect 42166 666729 42218 666735
rect 42166 666671 42218 666677
rect 42178 666148 42206 666671
rect 42164 665362 42220 665371
rect 42164 665297 42220 665306
rect 42178 664964 42206 665297
rect 42166 664879 42218 664885
rect 42166 664821 42218 664827
rect 42178 664298 42206 664821
rect 42166 664213 42218 664219
rect 42166 664155 42218 664161
rect 42178 664016 42206 664155
rect 42082 663988 42206 664016
rect 42082 663706 42110 663988
rect 42562 663553 42590 668849
rect 42850 664885 42878 668891
rect 42946 666735 42974 670593
rect 43234 668456 43262 670741
rect 43042 668428 43262 668456
rect 42934 666729 42986 666735
rect 42934 666671 42986 666677
rect 42932 666546 42988 666555
rect 42932 666481 42988 666490
rect 42838 664879 42890 664885
rect 42838 664821 42890 664827
rect 42838 664731 42890 664737
rect 42838 664673 42890 664679
rect 42550 663547 42602 663553
rect 42550 663489 42602 663495
rect 42548 663438 42604 663447
rect 42166 663399 42218 663405
rect 42548 663373 42604 663382
rect 42166 663341 42218 663347
rect 42178 663114 42206 663341
rect 42262 662437 42314 662443
rect 42262 662379 42314 662385
rect 41794 661375 41822 661856
rect 41780 661366 41836 661375
rect 41780 661301 41836 661310
rect 41890 661079 41918 661190
rect 42166 661105 42218 661111
rect 41876 661070 41932 661079
rect 42166 661047 42218 661053
rect 41876 661005 41932 661014
rect 42178 660908 42206 661047
rect 42082 660880 42206 660908
rect 42082 660672 42110 660880
rect 42274 660020 42302 662379
rect 42192 659992 42302 660020
rect 42166 659699 42218 659705
rect 42166 659641 42218 659647
rect 42178 659340 42206 659641
rect 42562 659113 42590 663373
rect 42850 661111 42878 664673
rect 42838 661105 42890 661111
rect 42838 661047 42890 661053
rect 42836 660922 42892 660931
rect 42836 660857 42892 660866
rect 42070 659107 42122 659113
rect 42070 659049 42122 659055
rect 42550 659107 42602 659113
rect 42550 659049 42602 659055
rect 42082 658822 42110 659049
rect 42082 656819 42110 656972
rect 42850 656893 42878 660857
rect 42946 659705 42974 666481
rect 43042 662443 43070 668428
rect 43124 668322 43180 668331
rect 43124 668257 43180 668266
rect 43138 664219 43166 668257
rect 43330 667919 43358 671333
rect 43318 667913 43370 667919
rect 43318 667855 43370 667861
rect 43126 664213 43178 664219
rect 43126 664155 43178 664161
rect 43126 664065 43178 664071
rect 43126 664007 43178 664013
rect 43030 662437 43082 662443
rect 43030 662379 43082 662385
rect 42934 659699 42986 659705
rect 42934 659641 42986 659647
rect 42166 656887 42218 656893
rect 42166 656829 42218 656835
rect 42838 656887 42890 656893
rect 42838 656829 42890 656835
rect 42070 656813 42122 656819
rect 42070 656755 42122 656761
rect 42178 656306 42206 656829
rect 43138 656819 43166 664007
rect 43126 656813 43178 656819
rect 43126 656755 43178 656761
rect 42838 656739 42890 656745
rect 42838 656681 42890 656687
rect 41780 656186 41836 656195
rect 41780 656121 41836 656130
rect 41794 655677 41822 656121
rect 42850 650867 42878 656681
rect 42836 650858 42892 650867
rect 42836 650793 42892 650802
rect 42452 649822 42508 649831
rect 42452 649757 42454 649766
rect 42506 649757 42508 649766
rect 42454 649725 42506 649731
rect 42454 649561 42506 649567
rect 42452 649526 42454 649535
rect 42506 649526 42508 649535
rect 42452 649461 42508 649470
rect 43220 648490 43276 648499
rect 43220 648425 43276 648434
rect 42548 645530 42604 645539
rect 42604 645488 42686 645516
rect 42548 645465 42604 645474
rect 40052 643902 40108 643911
rect 40052 643837 40108 643846
rect 40066 627885 40094 643837
rect 41684 642422 41740 642431
rect 41684 642357 41740 642366
rect 41492 641682 41548 641691
rect 41492 641617 41548 641626
rect 40054 627879 40106 627885
rect 40054 627821 40106 627827
rect 41206 627879 41258 627885
rect 41206 627821 41258 627827
rect 41218 627779 41246 627821
rect 41204 627770 41260 627779
rect 41506 627737 41534 641617
rect 41698 627811 41726 642357
rect 41780 640794 41836 640803
rect 41780 640729 41836 640738
rect 41686 627805 41738 627811
rect 41686 627747 41738 627753
rect 41204 627705 41260 627714
rect 41494 627731 41546 627737
rect 41494 627673 41546 627679
rect 41794 627441 41822 640729
rect 41876 639462 41932 639471
rect 41876 639397 41932 639406
rect 41890 627483 41918 639397
rect 42068 636798 42124 636807
rect 42068 636733 42124 636742
rect 41972 636354 42028 636363
rect 41972 636289 42028 636298
rect 41986 627631 42014 636289
rect 41972 627622 42028 627631
rect 41972 627557 42028 627566
rect 41876 627474 41932 627483
rect 41782 627435 41834 627441
rect 42082 627441 42110 636733
rect 42658 635919 42686 645488
rect 42932 638426 42988 638435
rect 42932 638361 42988 638370
rect 42644 635910 42700 635919
rect 42644 635845 42700 635854
rect 42164 633542 42220 633551
rect 42164 633477 42220 633486
rect 42178 632492 42206 633477
rect 42260 632506 42316 632515
rect 42178 632464 42260 632492
rect 42260 632441 42262 632450
rect 42314 632441 42316 632450
rect 42262 632409 42314 632415
rect 42946 628477 42974 638361
rect 43124 638130 43180 638139
rect 43124 638065 43180 638074
rect 42934 628471 42986 628477
rect 42934 628413 42986 628419
rect 42454 627953 42506 627959
rect 42454 627895 42506 627901
rect 41876 627409 41932 627418
rect 42070 627435 42122 627441
rect 41782 627377 41834 627383
rect 42070 627377 42122 627383
rect 41782 627213 41834 627219
rect 41782 627155 41834 627161
rect 41794 626632 41822 627155
rect 42164 625254 42220 625263
rect 42164 625189 42220 625198
rect 42178 624782 42206 625189
rect 42466 624703 42494 627895
rect 43138 627885 43166 638065
rect 43126 627879 43178 627885
rect 43126 627821 43178 627827
rect 43126 627731 43178 627737
rect 43126 627673 43178 627679
rect 43030 627435 43082 627441
rect 43030 627377 43082 627383
rect 42934 625215 42986 625221
rect 42934 625157 42986 625163
rect 42166 624697 42218 624703
rect 42166 624639 42218 624645
rect 42454 624697 42506 624703
rect 42454 624639 42506 624645
rect 42178 624161 42206 624639
rect 42452 624514 42508 624523
rect 42452 624449 42508 624458
rect 42166 623513 42218 623519
rect 42166 623455 42218 623461
rect 42178 622965 42206 623455
rect 42466 623371 42494 624449
rect 42946 623519 42974 625157
rect 42934 623513 42986 623519
rect 42934 623455 42986 623461
rect 42454 623365 42506 623371
rect 42454 623307 42506 623313
rect 42934 623365 42986 623371
rect 42934 623307 42986 623313
rect 42164 622146 42220 622155
rect 42164 622081 42220 622090
rect 42178 621748 42206 622081
rect 42166 621663 42218 621669
rect 42166 621605 42218 621611
rect 42178 621125 42206 621605
rect 42068 620962 42124 620971
rect 42068 620897 42124 620906
rect 42082 620490 42110 620897
rect 42452 620814 42508 620823
rect 42452 620749 42508 620758
rect 42166 620405 42218 620411
rect 42166 620347 42218 620353
rect 42178 619929 42206 620347
rect 41780 619186 41836 619195
rect 41780 619121 41836 619130
rect 41794 618640 41822 619121
rect 41876 618298 41932 618307
rect 41876 618233 41932 618242
rect 41890 617974 41918 618233
rect 42466 617895 42494 620749
rect 42836 618298 42892 618307
rect 42836 618233 42892 618242
rect 42740 618150 42796 618159
rect 42740 618085 42796 618094
rect 42070 617889 42122 617895
rect 42070 617831 42122 617837
rect 42454 617889 42506 617895
rect 42454 617831 42506 617837
rect 42082 617456 42110 617831
rect 42452 617706 42508 617715
rect 42452 617641 42508 617650
rect 42166 617223 42218 617229
rect 42166 617165 42218 617171
rect 42178 616790 42206 617165
rect 42166 616705 42218 616711
rect 42166 616647 42218 616653
rect 42178 616157 42206 616647
rect 42166 615891 42218 615897
rect 42166 615833 42218 615839
rect 42178 615606 42206 615833
rect 42166 614041 42218 614047
rect 42166 613983 42218 613989
rect 42178 613756 42206 613983
rect 42466 613677 42494 617641
rect 42166 613671 42218 613677
rect 42166 613613 42218 613619
rect 42454 613671 42506 613677
rect 42454 613613 42506 613619
rect 42178 613121 42206 613613
rect 42454 613523 42506 613529
rect 42454 613465 42506 613471
rect 42070 612857 42122 612863
rect 42070 612799 42122 612805
rect 42082 612498 42110 612799
rect 42466 606319 42494 613465
rect 42754 612863 42782 618085
rect 42850 614047 42878 618233
rect 42946 616711 42974 623307
rect 43042 621669 43070 627377
rect 43030 621663 43082 621669
rect 43030 621605 43082 621611
rect 43030 621515 43082 621521
rect 43030 621457 43082 621463
rect 42934 616705 42986 616711
rect 42934 616647 42986 616653
rect 43042 615897 43070 621457
rect 43138 620411 43166 627673
rect 43126 620405 43178 620411
rect 43126 620347 43178 620353
rect 43126 620257 43178 620263
rect 43126 620199 43178 620205
rect 43138 617229 43166 620199
rect 43126 617223 43178 617229
rect 43126 617165 43178 617171
rect 43030 615891 43082 615897
rect 43030 615833 43082 615839
rect 42838 614041 42890 614047
rect 42838 613983 42890 613989
rect 42742 612857 42794 612863
rect 42742 612799 42794 612805
rect 42742 607751 42794 607757
rect 42740 607716 42742 607725
rect 42794 607716 42796 607725
rect 42740 607651 42796 607660
rect 42740 606902 42796 606911
rect 42740 606837 42742 606846
rect 42794 606837 42796 606846
rect 42742 606805 42794 606811
rect 42452 606310 42508 606319
rect 42452 606245 42508 606254
rect 43234 604691 43262 648425
rect 43426 647611 43454 691641
rect 43604 679866 43660 679875
rect 43604 679801 43660 679810
rect 43510 670873 43562 670879
rect 43510 670815 43562 670821
rect 43522 664071 43550 670815
rect 43618 664737 43646 679801
rect 43606 664731 43658 664737
rect 43606 664673 43658 664679
rect 43510 664065 43562 664071
rect 43510 664007 43562 664013
rect 43412 647602 43468 647611
rect 43412 647537 43468 647546
rect 43316 646122 43372 646131
rect 43316 646057 43372 646066
rect 43220 604682 43276 604691
rect 43220 604617 43276 604626
rect 43330 602915 43358 646057
rect 43606 628471 43658 628477
rect 43606 628413 43658 628419
rect 43414 627879 43466 627885
rect 43414 627821 43466 627827
rect 43426 625221 43454 627821
rect 43510 627805 43562 627811
rect 43510 627747 43562 627753
rect 43414 625215 43466 625221
rect 43414 625157 43466 625163
rect 43522 621521 43550 627747
rect 43510 621515 43562 621521
rect 43510 621457 43562 621463
rect 43618 620263 43646 628413
rect 43606 620257 43658 620263
rect 43606 620199 43658 620205
rect 43508 605274 43564 605283
rect 43508 605209 43564 605218
rect 43316 602906 43372 602915
rect 43316 602841 43372 602850
rect 42932 602166 42988 602175
rect 42932 602101 42988 602110
rect 40052 600686 40108 600695
rect 40052 600621 40108 600630
rect 40066 586001 40094 600621
rect 41876 598466 41932 598475
rect 41876 598401 41932 598410
rect 41780 597578 41836 597587
rect 41780 597513 41836 597522
rect 40054 585995 40106 586001
rect 40054 585937 40106 585943
rect 41794 584225 41822 597513
rect 41890 584415 41918 598401
rect 41972 596246 42028 596255
rect 41972 596181 42028 596190
rect 41876 584406 41932 584415
rect 41876 584341 41932 584350
rect 41986 584267 42014 596181
rect 42068 595210 42124 595219
rect 42068 595145 42124 595154
rect 42082 584563 42110 595145
rect 42836 594914 42892 594923
rect 42836 594849 42892 594858
rect 42164 593730 42220 593739
rect 42164 593665 42220 593674
rect 42068 584554 42124 584563
rect 42068 584489 42124 584498
rect 41972 584258 42028 584267
rect 41782 584219 41834 584225
rect 42178 584225 42206 593665
rect 42452 592398 42508 592407
rect 42452 592333 42508 592342
rect 42466 586149 42494 592333
rect 42548 591954 42604 591963
rect 42604 591912 42686 591940
rect 42548 591889 42604 591898
rect 42548 590770 42604 590779
rect 42548 590705 42604 590714
rect 42562 589299 42590 590705
rect 42548 589290 42604 589299
rect 42548 589225 42550 589234
rect 42602 589225 42604 589234
rect 42550 589193 42602 589199
rect 42550 586587 42602 586593
rect 42550 586529 42602 586535
rect 42454 586143 42506 586149
rect 42454 586085 42506 586091
rect 42454 585995 42506 586001
rect 42454 585937 42506 585943
rect 42466 584563 42494 585937
rect 42562 585007 42590 586529
rect 42548 584998 42604 585007
rect 42548 584933 42604 584942
rect 42658 584836 42686 591912
rect 42850 585113 42878 594849
rect 42946 586635 42974 602101
rect 43028 599650 43084 599659
rect 43028 599585 43084 599594
rect 42932 586626 42988 586635
rect 43042 586593 43070 599585
rect 43124 593434 43180 593443
rect 43124 593369 43180 593378
rect 42932 586561 42988 586570
rect 43030 586587 43082 586593
rect 43030 586529 43082 586535
rect 43138 586464 43166 593369
rect 42946 586436 43166 586464
rect 42838 585107 42890 585113
rect 42838 585049 42890 585055
rect 42562 584817 42686 584836
rect 42550 584811 42686 584817
rect 42602 584808 42686 584811
rect 42550 584753 42602 584759
rect 42838 584737 42890 584743
rect 42838 584679 42890 584685
rect 42452 584554 42508 584563
rect 42452 584489 42508 584498
rect 42452 584258 42508 584267
rect 41972 584193 42028 584202
rect 42166 584219 42218 584225
rect 41782 584161 41834 584167
rect 42452 584193 42508 584202
rect 42166 584161 42218 584167
rect 41782 583997 41834 584003
rect 41782 583939 41834 583945
rect 41794 583445 41822 583939
rect 42466 582153 42494 584193
rect 42166 582147 42218 582153
rect 42166 582089 42218 582095
rect 42454 582147 42506 582153
rect 42454 582089 42506 582095
rect 42178 581605 42206 582089
rect 42850 581487 42878 584679
rect 42946 584415 42974 586436
rect 43030 586143 43082 586149
rect 43030 586085 43082 586091
rect 42932 584406 42988 584415
rect 42932 584341 42988 584350
rect 42934 584219 42986 584225
rect 42934 584161 42986 584167
rect 42070 581481 42122 581487
rect 42070 581423 42122 581429
rect 42838 581481 42890 581487
rect 42838 581423 42890 581429
rect 42082 580974 42110 581423
rect 42836 581298 42892 581307
rect 42836 581233 42892 581242
rect 42070 580297 42122 580303
rect 42070 580239 42122 580245
rect 42082 579790 42110 580239
rect 42166 579039 42218 579045
rect 42166 578981 42218 578987
rect 42178 578569 42206 578981
rect 42070 578447 42122 578453
rect 42070 578389 42122 578395
rect 42082 577940 42110 578389
rect 42166 577707 42218 577713
rect 42166 577649 42218 577655
rect 42178 577274 42206 577649
rect 41780 577154 41836 577163
rect 41780 577089 41836 577098
rect 41794 576756 41822 577089
rect 42452 577006 42508 577015
rect 42452 576941 42508 576950
rect 42262 576079 42314 576085
rect 42262 576021 42314 576027
rect 41794 574943 41822 575424
rect 41876 575082 41932 575091
rect 41876 575017 41932 575026
rect 41780 574934 41836 574943
rect 41780 574869 41836 574878
rect 41890 574797 41918 575017
rect 42274 574254 42302 576021
rect 42192 574226 42302 574254
rect 42260 574046 42316 574055
rect 42260 573981 42316 573990
rect 41780 573898 41836 573907
rect 41780 573833 41836 573842
rect 41794 573574 41822 573833
rect 42070 573489 42122 573495
rect 42070 573431 42122 573437
rect 42082 572982 42110 573431
rect 42166 572675 42218 572681
rect 42166 572617 42218 572623
rect 42178 572390 42206 572617
rect 42274 572533 42302 573981
rect 42466 572681 42494 576941
rect 42850 573495 42878 581233
rect 42946 578453 42974 584161
rect 42934 578447 42986 578453
rect 42934 578389 42986 578395
rect 42932 578338 42988 578347
rect 42932 578273 42988 578282
rect 42946 576085 42974 578273
rect 43042 577713 43070 586085
rect 43126 585107 43178 585113
rect 43126 585049 43178 585055
rect 43138 584984 43166 585049
rect 43138 584956 43262 584984
rect 43126 584811 43178 584817
rect 43126 584753 43178 584759
rect 43138 579045 43166 584753
rect 43234 580303 43262 584956
rect 43222 580297 43274 580303
rect 43222 580239 43274 580245
rect 43330 580081 43358 602841
rect 43318 580075 43370 580081
rect 43318 580017 43370 580023
rect 43126 579039 43178 579045
rect 43126 578981 43178 578987
rect 43030 577707 43082 577713
rect 43030 577649 43082 577655
rect 43028 577598 43084 577607
rect 43028 577533 43084 577542
rect 42934 576079 42986 576085
rect 42934 576021 42986 576027
rect 42838 573489 42890 573495
rect 42838 573431 42890 573437
rect 42836 573306 42892 573315
rect 42836 573241 42892 573250
rect 42454 572675 42506 572681
rect 42454 572617 42506 572623
rect 42262 572527 42314 572533
rect 42262 572469 42314 572475
rect 42454 572527 42506 572533
rect 42454 572469 42506 572475
rect 42166 571047 42218 571053
rect 42166 570989 42218 570995
rect 42178 570540 42206 570989
rect 42358 570307 42410 570313
rect 42358 570249 42410 570255
rect 42070 570233 42122 570239
rect 42070 570175 42122 570181
rect 42082 569948 42110 570175
rect 42070 569715 42122 569721
rect 42070 569657 42122 569663
rect 42082 569282 42110 569657
rect 34484 564722 34540 564731
rect 34484 564657 34540 564666
rect 34498 564541 34526 564657
rect 34486 564535 34538 564541
rect 34486 564477 34538 564483
rect 42370 563103 42398 570249
rect 42466 570239 42494 572469
rect 42454 570233 42506 570239
rect 42454 570175 42506 570181
rect 42850 569721 42878 573241
rect 43042 571053 43070 577533
rect 43030 571047 43082 571053
rect 43030 570989 43082 570995
rect 42838 569715 42890 569721
rect 42838 569657 42890 569663
rect 43316 564574 43372 564583
rect 43316 564509 43372 564518
rect 42452 563538 42508 563547
rect 42452 563473 42454 563482
rect 42506 563473 42508 563482
rect 42454 563441 42506 563447
rect 42356 563094 42412 563103
rect 42356 563029 42412 563038
rect 43220 562058 43276 562067
rect 43220 561993 43276 562002
rect 41972 558654 42028 558663
rect 41972 558589 42028 558598
rect 40148 557470 40204 557479
rect 40148 557405 40204 557414
rect 40162 542933 40190 557405
rect 41684 555990 41740 555999
rect 41684 555925 41740 555934
rect 40150 542927 40202 542933
rect 40150 542869 40202 542875
rect 41698 541305 41726 555925
rect 41876 555250 41932 555259
rect 41876 555185 41932 555194
rect 41780 554362 41836 554371
rect 41780 554297 41836 554306
rect 41686 541299 41738 541305
rect 41686 541241 41738 541247
rect 41794 541009 41822 554297
rect 41890 541347 41918 555185
rect 41986 544635 42014 558589
rect 42068 553030 42124 553039
rect 42068 552965 42124 552974
rect 41974 544629 42026 544635
rect 41974 544571 42026 544577
rect 41974 542927 42026 542933
rect 41974 542869 42026 542875
rect 41876 541338 41932 541347
rect 41876 541273 41932 541282
rect 41986 541199 42014 542869
rect 41972 541190 42028 541199
rect 41972 541125 42028 541134
rect 42082 541051 42110 552965
rect 42356 551994 42412 552003
rect 42356 551929 42412 551938
rect 42164 550070 42220 550079
rect 42164 550005 42220 550014
rect 42068 541042 42124 541051
rect 41782 541003 41834 541009
rect 42178 541009 42206 550005
rect 42370 545597 42398 551929
rect 42932 551698 42988 551707
rect 42932 551633 42988 551642
rect 42836 551106 42892 551115
rect 42836 551041 42892 551050
rect 42644 546296 42700 546305
rect 42644 546231 42646 546240
rect 42698 546231 42700 546240
rect 42646 546199 42698 546205
rect 42358 545591 42410 545597
rect 42358 545533 42410 545539
rect 42646 545591 42698 545597
rect 42646 545533 42698 545539
rect 42068 540977 42124 540986
rect 42166 541003 42218 541009
rect 41782 540945 41834 540951
rect 42166 540945 42218 540951
rect 41782 540781 41834 540787
rect 41782 540723 41834 540729
rect 41794 540245 41822 540723
rect 42068 538970 42124 538979
rect 42068 538905 42124 538914
rect 42082 538424 42110 538905
rect 42166 538191 42218 538197
rect 42166 538133 42218 538139
rect 42178 537758 42206 538133
rect 42070 537081 42122 537087
rect 42070 537023 42122 537029
rect 42082 536574 42110 537023
rect 42070 535823 42122 535829
rect 42070 535765 42122 535771
rect 42082 535390 42110 535765
rect 42166 535305 42218 535311
rect 42166 535247 42218 535253
rect 42178 534724 42206 535247
rect 42166 534491 42218 534497
rect 42166 534433 42218 534439
rect 42178 534058 42206 534433
rect 42070 533751 42122 533757
rect 42070 533693 42122 533699
rect 42082 533540 42110 533693
rect 42658 532869 42686 545533
rect 42850 544876 42878 551041
rect 42754 544848 42878 544876
rect 42754 535311 42782 544848
rect 42946 544728 42974 551633
rect 43028 549330 43084 549339
rect 43028 549265 43084 549274
rect 42850 544700 42974 544728
rect 42850 537087 42878 544700
rect 42934 544629 42986 544635
rect 42934 544571 42986 544577
rect 42946 538789 42974 544571
rect 42934 538783 42986 538789
rect 42934 538725 42986 538731
rect 42932 538674 42988 538683
rect 42932 538609 42988 538618
rect 42838 537081 42890 537087
rect 42838 537023 42890 537029
rect 42836 536898 42892 536907
rect 42836 536833 42892 536842
rect 42742 535305 42794 535311
rect 42742 535247 42794 535253
rect 42262 532863 42314 532869
rect 42262 532805 42314 532811
rect 42646 532863 42698 532869
rect 42646 532805 42698 532811
rect 41794 531727 41822 532241
rect 41780 531718 41836 531727
rect 41780 531653 41836 531662
rect 41890 531283 41918 531616
rect 42166 531383 42218 531389
rect 42166 531325 42218 531331
rect 41876 531274 41932 531283
rect 41876 531209 41932 531218
rect 42178 531024 42206 531325
rect 42274 530415 42302 532805
rect 42644 532606 42700 532615
rect 42644 532541 42700 532550
rect 42192 530387 42302 530415
rect 42262 530347 42314 530353
rect 42262 530289 42314 530295
rect 42274 529780 42302 530289
rect 42192 529752 42302 529780
rect 42262 529681 42314 529687
rect 42262 529623 42314 529629
rect 42274 529219 42302 529623
rect 42192 529191 42302 529219
rect 42166 527683 42218 527689
rect 42166 527625 42218 527631
rect 42178 527365 42206 527625
rect 42658 527245 42686 532541
rect 42740 532310 42796 532319
rect 42740 532245 42796 532254
rect 42070 527239 42122 527245
rect 42070 527181 42122 527187
rect 42646 527239 42698 527245
rect 42646 527181 42698 527187
rect 42082 526732 42110 527181
rect 42358 527091 42410 527097
rect 42358 527033 42410 527039
rect 42166 526499 42218 526505
rect 42166 526441 42218 526447
rect 42178 526066 42206 526441
rect 42370 435527 42398 527033
rect 42754 526505 42782 532245
rect 42850 530353 42878 536833
rect 42946 533757 42974 538609
rect 43042 534497 43070 549265
rect 43124 548590 43180 548599
rect 43124 548525 43180 548534
rect 43138 535829 43166 548525
rect 43234 535829 43262 561993
rect 43330 561304 43358 564509
rect 43522 561623 43550 605209
rect 43606 580075 43658 580081
rect 43606 580017 43658 580023
rect 43618 564583 43646 580017
rect 43604 564574 43660 564583
rect 43604 564509 43660 564518
rect 43508 561614 43564 561623
rect 43508 561549 43564 561558
rect 43330 561276 43646 561304
rect 43618 559847 43646 561276
rect 43796 560578 43852 560587
rect 43796 560513 43852 560522
rect 43604 559838 43660 559847
rect 43604 559773 43660 559782
rect 43414 541299 43466 541305
rect 43414 541241 43466 541247
rect 43318 541003 43370 541009
rect 43318 540945 43370 540951
rect 43126 535823 43178 535829
rect 43126 535765 43178 535771
rect 43222 535823 43274 535829
rect 43222 535765 43274 535771
rect 43330 535700 43358 540945
rect 43138 535672 43358 535700
rect 43030 534491 43082 534497
rect 43030 534433 43082 534439
rect 43030 534343 43082 534349
rect 43030 534285 43082 534291
rect 42934 533751 42986 533757
rect 42934 533693 42986 533699
rect 42934 533603 42986 533609
rect 42934 533545 42986 533551
rect 42838 530347 42890 530353
rect 42838 530289 42890 530295
rect 42946 527689 42974 533545
rect 43042 529687 43070 534285
rect 43138 531389 43166 535672
rect 43222 535601 43274 535607
rect 43222 535543 43274 535549
rect 43126 531383 43178 531389
rect 43126 531325 43178 531331
rect 43030 529681 43082 529687
rect 43030 529623 43082 529629
rect 42934 527683 42986 527689
rect 42934 527625 42986 527631
rect 42742 526499 42794 526505
rect 42742 526441 42794 526447
rect 42646 436959 42698 436965
rect 42644 436924 42646 436933
rect 42698 436924 42700 436933
rect 42644 436859 42700 436868
rect 42646 436145 42698 436151
rect 42644 436110 42646 436119
rect 42698 436110 42700 436119
rect 42644 436045 42700 436054
rect 42356 435518 42412 435527
rect 42356 435453 42412 435462
rect 43234 433603 43262 535543
rect 43426 534349 43454 541241
rect 43510 538783 43562 538789
rect 43510 538725 43562 538731
rect 43414 534343 43466 534349
rect 43414 534285 43466 534291
rect 43522 533609 43550 538725
rect 43510 533603 43562 533609
rect 43510 533545 43562 533551
rect 43412 434482 43468 434491
rect 43412 434417 43468 434426
rect 43220 433594 43276 433603
rect 43220 433529 43276 433538
rect 41876 429894 41932 429903
rect 41876 429829 41932 429838
rect 41780 426786 41836 426795
rect 41780 426721 41836 426730
rect 41794 413433 41822 426721
rect 41890 420019 41918 429829
rect 43426 429140 43454 434417
rect 43618 432123 43646 559773
rect 43702 541521 43754 541527
rect 43702 541463 43754 541469
rect 43714 538197 43742 541463
rect 43702 538191 43754 538197
rect 43702 538133 43754 538139
rect 43810 433011 43838 560513
rect 43796 433002 43852 433011
rect 43796 432937 43852 432946
rect 43604 432114 43660 432123
rect 43604 432049 43660 432058
rect 43234 429112 43454 429140
rect 43124 424418 43180 424427
rect 43124 424353 43180 424362
rect 42740 424122 42796 424131
rect 42740 424057 42796 424066
rect 42164 423234 42220 423243
rect 42164 423169 42220 423178
rect 41878 420013 41930 420019
rect 41878 419955 41930 419961
rect 42178 413581 42206 423169
rect 42644 420126 42700 420135
rect 42644 420061 42700 420070
rect 42358 420013 42410 420019
rect 42358 419955 42410 419961
rect 42166 413575 42218 413581
rect 42166 413517 42218 413523
rect 41782 413427 41834 413433
rect 41782 413369 41834 413375
rect 41782 413205 41834 413211
rect 41782 413147 41834 413153
rect 41794 412624 41822 413147
rect 42370 411361 42398 419955
rect 42658 418655 42686 420061
rect 42644 418646 42700 418655
rect 42644 418581 42646 418590
rect 42698 418581 42700 418590
rect 42646 418549 42698 418555
rect 42166 411355 42218 411361
rect 42166 411297 42218 411303
rect 42358 411355 42410 411361
rect 42358 411297 42410 411303
rect 42178 410805 42206 411297
rect 42358 411207 42410 411213
rect 42358 411149 42410 411155
rect 42070 410541 42122 410547
rect 42070 410483 42122 410489
rect 42082 410182 42110 410483
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42178 408965 42206 409447
rect 42166 408247 42218 408253
rect 42166 408189 42218 408195
rect 42178 407769 42206 408189
rect 42070 407507 42122 407513
rect 42070 407449 42122 407455
rect 42082 407148 42110 407449
rect 42166 406915 42218 406921
rect 42166 406857 42218 406863
rect 42178 406482 42206 406857
rect 41780 406066 41836 406075
rect 41780 406001 41836 406010
rect 41794 405929 41822 406001
rect 41794 404299 41822 404632
rect 41780 404290 41836 404299
rect 41780 404225 41836 404234
rect 42082 403855 42110 403997
rect 42166 403881 42218 403887
rect 42068 403846 42124 403855
rect 42166 403823 42218 403829
rect 42068 403781 42124 403790
rect 42178 403448 42206 403823
rect 42370 402999 42398 411149
rect 42754 409511 42782 424057
rect 42932 422642 42988 422651
rect 42932 422577 42988 422586
rect 42836 421014 42892 421023
rect 42836 420949 42892 420958
rect 42742 409505 42794 409511
rect 42742 409447 42794 409453
rect 42850 408253 42878 420949
rect 42838 408247 42890 408253
rect 42838 408189 42890 408195
rect 42946 403887 42974 422577
rect 43028 421310 43084 421319
rect 43028 421245 43084 421254
rect 43042 406921 43070 421245
rect 43138 411213 43166 424353
rect 43234 419076 43262 429112
rect 43234 419048 43358 419076
rect 43222 413575 43274 413581
rect 43222 413517 43274 413523
rect 43126 411207 43178 411213
rect 43126 411149 43178 411155
rect 43234 411084 43262 413517
rect 43138 411056 43262 411084
rect 43138 407513 43166 411056
rect 43126 407507 43178 407513
rect 43126 407449 43178 407455
rect 43030 406915 43082 406921
rect 43030 406857 43082 406863
rect 42934 403881 42986 403887
rect 42934 403823 42986 403829
rect 42070 402993 42122 402999
rect 42070 402935 42122 402941
rect 42358 402993 42410 402999
rect 42358 402935 42410 402941
rect 42082 402782 42110 402935
rect 41780 402514 41836 402523
rect 41780 402449 41836 402458
rect 41794 402157 41822 402449
rect 41780 402070 41836 402079
rect 41780 402005 41836 402014
rect 41794 401598 41822 402005
rect 41780 400146 41836 400155
rect 41780 400081 41836 400090
rect 41794 399748 41822 400081
rect 41780 399554 41836 399563
rect 41780 399489 41836 399498
rect 41794 399121 41822 399489
rect 41780 398814 41836 398823
rect 41780 398749 41836 398758
rect 41794 398490 41822 398749
rect 42358 393965 42410 393971
rect 42356 393930 42358 393939
rect 42410 393930 42412 393939
rect 42356 393865 42412 393874
rect 42358 393225 42410 393231
rect 42356 393190 42358 393199
rect 42410 393190 42412 393199
rect 42356 393125 42412 393134
rect 42358 392337 42410 392343
rect 42356 392302 42358 392311
rect 42410 392302 42412 392311
rect 42356 392237 42412 392246
rect 43220 391266 43276 391275
rect 43220 391201 43276 391210
rect 42068 386678 42124 386687
rect 42068 386613 42124 386622
rect 37364 380018 37420 380027
rect 37364 379953 37420 379962
rect 37378 372585 37406 379953
rect 37366 372579 37418 372585
rect 37366 372521 37418 372527
rect 42082 370217 42110 386613
rect 42356 383570 42412 383579
rect 42356 383505 42412 383514
rect 42260 378834 42316 378843
rect 42260 378769 42316 378778
rect 42164 376614 42220 376623
rect 42164 376549 42220 376558
rect 42178 375291 42206 376549
rect 42164 375282 42220 375291
rect 42164 375217 42166 375226
rect 42218 375217 42220 375226
rect 42166 375185 42218 375191
rect 42274 370217 42302 378769
rect 42070 370211 42122 370217
rect 42070 370153 42122 370159
rect 42262 370211 42314 370217
rect 42262 370153 42314 370159
rect 42370 369995 42398 383505
rect 42836 381794 42892 381803
rect 42836 381729 42892 381738
rect 42740 377798 42796 377807
rect 42740 377733 42796 377742
rect 42166 369989 42218 369995
rect 42166 369931 42218 369937
rect 42358 369989 42410 369995
rect 42358 369931 42410 369937
rect 42178 369445 42206 369931
rect 42358 369841 42410 369847
rect 42358 369783 42410 369789
rect 42370 368145 42398 369783
rect 42070 368139 42122 368145
rect 42070 368081 42122 368087
rect 42358 368139 42410 368145
rect 42358 368081 42410 368087
rect 42082 367632 42110 368081
rect 42070 367399 42122 367405
rect 42070 367341 42122 367347
rect 42082 366966 42110 367341
rect 42070 366289 42122 366295
rect 42070 366231 42122 366237
rect 42082 365782 42110 366231
rect 42754 365037 42782 377733
rect 42166 365031 42218 365037
rect 42166 364973 42218 364979
rect 42742 365031 42794 365037
rect 42742 364973 42794 364979
rect 42178 364569 42206 364973
rect 42070 364291 42122 364297
rect 42070 364233 42122 364239
rect 42082 363932 42110 364233
rect 42850 364149 42878 381729
rect 43028 380906 43084 380915
rect 43028 380841 43084 380850
rect 42934 372579 42986 372585
rect 42934 372521 42986 372527
rect 42946 364297 42974 372521
rect 43042 366295 43070 380841
rect 43124 378538 43180 378547
rect 43124 378473 43180 378482
rect 43030 366289 43082 366295
rect 43030 366231 43082 366237
rect 43030 366141 43082 366147
rect 43030 366083 43082 366089
rect 42934 364291 42986 364297
rect 42934 364233 42986 364239
rect 42358 364143 42410 364149
rect 42358 364085 42410 364091
rect 42838 364143 42890 364149
rect 42838 364085 42890 364091
rect 42166 363699 42218 363705
rect 42166 363641 42218 363647
rect 42178 363266 42206 363641
rect 41780 362850 41836 362859
rect 41780 362785 41836 362794
rect 41794 362748 41822 362785
rect 42262 362145 42314 362151
rect 42262 362087 42314 362093
rect 42082 360935 42110 361416
rect 42068 360926 42124 360935
rect 42068 360861 42124 360870
rect 41794 360639 41822 360824
rect 41780 360630 41836 360639
rect 41780 360565 41836 360574
rect 42274 360246 42302 362087
rect 42192 360218 42302 360246
rect 42370 359615 42398 364085
rect 43042 362151 43070 366083
rect 43138 363705 43166 378473
rect 43126 363699 43178 363705
rect 43126 363641 43178 363647
rect 43030 362145 43082 362151
rect 43030 362087 43082 362093
rect 42192 359587 42398 359615
rect 42068 359446 42124 359455
rect 42068 359381 42124 359390
rect 42082 358974 42110 359381
rect 41780 358706 41836 358715
rect 41780 358641 41836 358650
rect 41794 358382 41822 358641
rect 41876 356930 41932 356939
rect 41876 356865 41932 356874
rect 41890 356565 41918 356865
rect 41780 356486 41836 356495
rect 41780 356421 41836 356430
rect 41794 355940 41822 356421
rect 41780 355598 41836 355607
rect 41780 355533 41836 355542
rect 41794 355274 41822 355533
rect 42358 350749 42410 350755
rect 42356 350714 42358 350723
rect 42410 350714 42412 350723
rect 42356 350649 42412 350658
rect 42646 349713 42698 349719
rect 42644 349678 42646 349687
rect 42698 349678 42700 349687
rect 42644 349613 42700 349622
rect 42358 349121 42410 349127
rect 42356 349086 42358 349095
rect 42410 349086 42412 349095
rect 42356 349021 42412 349030
rect 43234 347763 43262 391201
rect 43330 390979 43358 419048
rect 43316 390970 43372 390979
rect 43316 390905 43372 390914
rect 43318 370211 43370 370217
rect 43318 370153 43370 370159
rect 43330 366147 43358 370153
rect 43318 366141 43370 366147
rect 43318 366083 43370 366089
rect 43316 348050 43372 348059
rect 43316 347985 43372 347994
rect 43220 347754 43276 347763
rect 43220 347689 43276 347698
rect 42740 344128 42796 344137
rect 42740 344063 42796 344072
rect 37268 340354 37324 340363
rect 37268 340289 37324 340298
rect 37172 337246 37228 337255
rect 37172 337181 37228 337190
rect 37186 328407 37214 337181
rect 37282 329369 37310 340289
rect 37364 337246 37420 337255
rect 37364 337181 37420 337190
rect 37270 329363 37322 329369
rect 37270 329305 37322 329311
rect 37378 329221 37406 337181
rect 42356 333398 42412 333407
rect 42356 333333 42412 333342
rect 42370 332075 42398 333333
rect 42356 332066 42412 332075
rect 42356 332001 42358 332010
rect 42410 332001 42412 332010
rect 42358 331969 42410 331975
rect 41782 329363 41834 329369
rect 41782 329305 41834 329311
rect 37366 329215 37418 329221
rect 37366 329157 37418 329163
rect 41686 329215 41738 329221
rect 41686 329157 41738 329163
rect 37174 328401 37226 328407
rect 37174 328343 37226 328349
rect 41698 327297 41726 329157
rect 41686 327291 41738 327297
rect 41686 327233 41738 327239
rect 41794 327075 41822 329305
rect 42358 327291 42410 327297
rect 42358 327233 42410 327239
rect 41782 327069 41834 327075
rect 41782 327011 41834 327017
rect 41782 326773 41834 326779
rect 41782 326715 41834 326721
rect 41794 326266 41822 326715
rect 42070 324923 42122 324929
rect 42070 324865 42122 324871
rect 42082 324416 42110 324865
rect 42166 324183 42218 324189
rect 42166 324125 42218 324131
rect 42178 323750 42206 324125
rect 42166 323147 42218 323153
rect 42166 323089 42218 323095
rect 42178 322566 42206 323089
rect 42070 321815 42122 321821
rect 42070 321757 42122 321763
rect 42082 321382 42110 321757
rect 42370 321303 42398 327233
rect 42754 324929 42782 344063
rect 43124 335470 43180 335479
rect 43124 335405 43180 335414
rect 43028 334582 43084 334591
rect 43028 334517 43084 334526
rect 43042 328204 43070 334517
rect 43138 328333 43166 335405
rect 43330 329388 43358 347985
rect 43412 338578 43468 338587
rect 43412 338513 43468 338522
rect 43234 329360 43358 329388
rect 43126 328327 43178 328333
rect 43126 328269 43178 328275
rect 43042 328176 43166 328204
rect 43030 328105 43082 328111
rect 43030 328047 43082 328053
rect 42742 324923 42794 324929
rect 42742 324865 42794 324871
rect 43042 323153 43070 328047
rect 43030 323147 43082 323153
rect 43030 323089 43082 323095
rect 43030 322999 43082 323005
rect 43030 322941 43082 322947
rect 42166 321297 42218 321303
rect 42166 321239 42218 321245
rect 42358 321297 42410 321303
rect 42358 321239 42410 321245
rect 42178 320716 42206 321239
rect 43042 320637 43070 322941
rect 43138 321821 43166 328176
rect 43126 321815 43178 321821
rect 43126 321757 43178 321763
rect 42166 320631 42218 320637
rect 42166 320573 42218 320579
rect 43030 320631 43082 320637
rect 43030 320573 43082 320579
rect 42178 320081 42206 320573
rect 41780 319782 41836 319791
rect 41780 319717 41836 319726
rect 41794 319532 41822 319717
rect 42164 318746 42220 318755
rect 42164 318681 42220 318690
rect 42178 318241 42206 318681
rect 41780 318006 41836 318015
rect 41780 317941 41836 317950
rect 41794 317608 41822 317941
rect 41876 317414 41932 317423
rect 41876 317349 41932 317358
rect 41890 317045 41918 317349
rect 42070 316931 42122 316937
rect 42070 316873 42122 316879
rect 42082 316424 42110 316873
rect 41780 316082 41836 316091
rect 41780 316017 41836 316026
rect 41794 315758 41822 316017
rect 41780 315638 41836 315647
rect 41780 315573 41836 315582
rect 41794 315205 41822 315573
rect 41780 313714 41836 313723
rect 41780 313649 41836 313658
rect 41794 313390 41822 313649
rect 41780 313270 41836 313279
rect 41780 313205 41836 313214
rect 41794 312724 41822 313205
rect 41780 312382 41836 312391
rect 41780 312317 41836 312326
rect 41794 312058 41822 312317
rect 42262 307533 42314 307539
rect 42260 307498 42262 307507
rect 42314 307498 42316 307507
rect 42260 307433 42316 307442
rect 42262 306793 42314 306799
rect 42260 306758 42262 306767
rect 42314 306758 42316 306767
rect 42260 306693 42316 306702
rect 42836 305722 42892 305731
rect 42836 305657 42892 305666
rect 42850 305541 42878 305657
rect 42838 305535 42890 305541
rect 42838 305477 42890 305483
rect 43234 304103 43262 329360
rect 43318 328327 43370 328333
rect 43318 328269 43370 328275
rect 43330 323005 43358 328269
rect 43318 322999 43370 323005
rect 43318 322941 43370 322947
rect 43426 316937 43454 338513
rect 43414 316931 43466 316937
rect 43414 316873 43466 316879
rect 43412 304834 43468 304843
rect 43412 304769 43468 304778
rect 43220 304094 43276 304103
rect 43220 304029 43276 304038
rect 39956 300394 40012 300403
rect 39956 300329 40012 300338
rect 37364 294030 37420 294039
rect 37364 293965 37420 293974
rect 37378 286893 37406 293965
rect 39970 288003 39998 300329
rect 41780 297286 41836 297295
rect 41780 297221 41836 297230
rect 39958 287997 40010 288003
rect 39958 287939 40010 287945
rect 37366 286887 37418 286893
rect 37366 286829 37418 286835
rect 41794 283859 41822 297221
rect 42164 294770 42220 294779
rect 42164 294705 42220 294714
rect 42178 283859 42206 294705
rect 43124 293882 43180 293891
rect 43124 293817 43180 293826
rect 42260 292402 42316 292411
rect 42260 292337 42316 292346
rect 41782 283853 41834 283859
rect 41782 283795 41834 283801
rect 42166 283853 42218 283859
rect 42166 283795 42218 283801
rect 42274 283679 42302 292337
rect 42836 292254 42892 292263
rect 42836 292189 42892 292198
rect 42548 290922 42604 290931
rect 42548 290857 42604 290866
rect 42260 283670 42316 283679
rect 42260 283605 42316 283614
rect 41782 283409 41834 283415
rect 41782 283351 41834 283357
rect 41794 283050 41822 283351
rect 42166 281781 42218 281787
rect 42166 281723 42218 281729
rect 42178 281200 42206 281723
rect 42166 281115 42218 281121
rect 42166 281057 42218 281063
rect 42178 280534 42206 281057
rect 42166 279931 42218 279937
rect 42166 279873 42218 279879
rect 42178 279350 42206 279873
rect 42562 278605 42590 290857
rect 42644 289146 42700 289155
rect 42644 289081 42646 289090
rect 42698 289081 42700 289090
rect 42646 289049 42698 289055
rect 42646 287997 42698 288003
rect 42646 287939 42698 287945
rect 42658 281787 42686 287939
rect 42742 286887 42794 286893
rect 42742 286829 42794 286835
rect 42646 281781 42698 281787
rect 42646 281723 42698 281729
rect 42644 281598 42700 281607
rect 42644 281533 42700 281542
rect 42658 279808 42686 281533
rect 42754 279937 42782 286829
rect 42742 279931 42794 279937
rect 42742 279873 42794 279879
rect 42658 279780 42782 279808
rect 42166 278599 42218 278605
rect 42166 278541 42218 278547
rect 42550 278599 42602 278605
rect 42550 278541 42602 278547
rect 42178 278166 42206 278541
rect 42166 277859 42218 277865
rect 42166 277801 42218 277807
rect 42178 277500 42206 277801
rect 42070 277415 42122 277421
rect 42070 277357 42122 277363
rect 42082 276908 42110 277357
rect 41780 276566 41836 276575
rect 41780 276501 41836 276510
rect 41794 276316 41822 276501
rect 41986 274799 42014 275058
rect 41972 274790 42028 274799
rect 41972 274725 42028 274734
rect 42754 274535 42782 279780
rect 42850 277421 42878 292189
rect 43138 277865 43166 293817
rect 43220 290626 43276 290635
rect 43220 290561 43276 290570
rect 43234 289113 43262 290561
rect 43222 289107 43274 289113
rect 43222 289049 43274 289055
rect 43426 288984 43454 304769
rect 43234 288956 43454 288984
rect 43234 277865 43262 288956
rect 43318 283853 43370 283859
rect 43318 283795 43370 283801
rect 43126 277859 43178 277865
rect 43126 277801 43178 277807
rect 43222 277859 43274 277865
rect 43222 277801 43274 277807
rect 43330 277736 43358 283795
rect 43138 277708 43358 277736
rect 42838 277415 42890 277421
rect 42838 277357 42890 277363
rect 42262 274529 42314 274535
rect 42262 274471 42314 274477
rect 42742 274529 42794 274535
rect 42742 274471 42794 274477
rect 41986 274059 42014 274392
rect 41972 274050 42028 274059
rect 41972 273985 42028 273994
rect 42274 273859 42302 274471
rect 42192 273831 42302 273859
rect 43138 273795 43166 277708
rect 43222 277637 43274 277643
rect 43222 277579 43274 277585
rect 42262 273789 42314 273795
rect 42262 273731 42314 273737
rect 43126 273789 43178 273795
rect 43126 273731 43178 273737
rect 42274 273222 42302 273731
rect 42192 273194 42302 273222
rect 41780 272866 41836 272875
rect 41780 272801 41836 272810
rect 41794 272542 41822 272801
rect 41780 272422 41836 272431
rect 41780 272357 41836 272366
rect 41794 272024 41822 272357
rect 41780 270646 41836 270655
rect 41780 270581 41836 270590
rect 41794 270174 41822 270581
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 41780 269166 41836 269175
rect 41780 269101 41836 269110
rect 41794 268877 41822 269101
rect 42262 264317 42314 264323
rect 42260 264282 42262 264291
rect 42314 264282 42316 264291
rect 42260 264217 42316 264226
rect 42262 263577 42314 263583
rect 42260 263542 42262 263551
rect 42314 263542 42316 263551
rect 42260 263477 42316 263486
rect 42836 262506 42892 262515
rect 42836 262441 42892 262450
rect 42850 262325 42878 262441
rect 42838 262319 42890 262325
rect 42838 262261 42890 262267
rect 43234 260887 43262 277579
rect 43316 264874 43372 264883
rect 43316 264809 43372 264818
rect 43220 260878 43276 260887
rect 43220 260813 43276 260822
rect 43330 260147 43358 264809
rect 43796 261618 43852 261627
rect 43796 261553 43852 261562
rect 43316 260138 43372 260147
rect 43316 260073 43372 260082
rect 42260 257178 42316 257187
rect 42260 257113 42316 257122
rect 37268 254070 37324 254079
rect 37268 254005 37324 254014
rect 37172 250814 37228 250823
rect 37172 250749 37228 250758
rect 34582 247667 34634 247673
rect 34582 247609 34634 247615
rect 34594 247123 34622 247609
rect 34580 247114 34636 247123
rect 34580 247049 34636 247058
rect 34594 246087 34622 247049
rect 34580 246078 34636 246087
rect 34580 246013 34636 246022
rect 37186 242049 37214 250749
rect 37282 244491 37310 254005
rect 41972 251554 42028 251563
rect 41972 251489 42028 251498
rect 37364 250814 37420 250823
rect 37364 250749 37420 250758
rect 37270 244485 37322 244491
rect 37270 244427 37322 244433
rect 37174 242043 37226 242049
rect 37174 241985 37226 241991
rect 37378 241975 37406 250749
rect 41782 244485 41834 244491
rect 41782 244427 41834 244433
rect 37366 241969 37418 241975
rect 37366 241911 37418 241917
rect 41794 240643 41822 244427
rect 41986 242345 42014 251489
rect 42166 250627 42218 250633
rect 42166 250569 42218 250575
rect 42068 248446 42124 248455
rect 42068 248381 42124 248390
rect 42082 244787 42110 248381
rect 42178 247673 42206 250569
rect 42166 247667 42218 247673
rect 42166 247609 42218 247615
rect 42070 244781 42122 244787
rect 42070 244723 42122 244729
rect 41974 242339 42026 242345
rect 41974 242281 42026 242287
rect 41782 240637 41834 240643
rect 41782 240579 41834 240585
rect 42274 240588 42302 257113
rect 43124 249778 43180 249787
rect 43124 249713 43180 249722
rect 43028 248150 43084 248159
rect 43028 248085 43084 248094
rect 42550 244781 42602 244787
rect 42550 244723 42602 244729
rect 42274 240560 42398 240588
rect 41782 240415 41834 240421
rect 41782 240357 41834 240363
rect 41794 239834 41822 240357
rect 42370 238571 42398 240560
rect 42166 238565 42218 238571
rect 42166 238507 42218 238513
rect 42358 238565 42410 238571
rect 42358 238507 42410 238513
rect 42178 237984 42206 238507
rect 42562 238497 42590 244723
rect 42742 242339 42794 242345
rect 42742 242281 42794 242287
rect 42646 242043 42698 242049
rect 42646 241985 42698 241991
rect 42658 240759 42686 241985
rect 42754 240791 42782 242281
rect 42742 240785 42794 240791
rect 42644 240750 42700 240759
rect 42742 240727 42794 240733
rect 42644 240685 42700 240694
rect 42550 238491 42602 238497
rect 42550 238433 42602 238439
rect 42358 238417 42410 238423
rect 42358 238359 42410 238365
rect 42166 237751 42218 237757
rect 42166 237693 42218 237699
rect 42178 237361 42206 237693
rect 42166 236715 42218 236721
rect 42166 236657 42218 236663
rect 42178 236165 42206 236657
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42164 234830 42220 234839
rect 42370 234816 42398 238359
rect 43042 235463 43070 248085
rect 43138 242123 43166 249713
rect 43126 242117 43178 242123
rect 43126 242059 43178 242065
rect 43126 241969 43178 241975
rect 43126 241911 43178 241917
rect 43138 236721 43166 241911
rect 43222 240785 43274 240791
rect 43222 240727 43274 240733
rect 43126 236715 43178 236721
rect 43126 236657 43178 236663
rect 43234 236592 43262 240727
rect 43138 236564 43262 236592
rect 43030 235457 43082 235463
rect 43030 235399 43082 235405
rect 42370 234788 42494 234816
rect 42164 234765 42220 234774
rect 42178 234325 42206 234765
rect 42358 234717 42410 234723
rect 42358 234659 42410 234665
rect 42070 234051 42122 234057
rect 42070 233993 42122 233999
rect 42082 233692 42110 233993
rect 41780 233350 41836 233359
rect 41780 233285 41836 233294
rect 41794 233129 41822 233285
rect 41780 231722 41836 231731
rect 41780 231657 41836 231666
rect 41794 231176 41822 231657
rect 41890 231583 41918 231842
rect 41876 231574 41932 231583
rect 41876 231509 41932 231518
rect 42370 230672 42398 234659
rect 42466 234205 42494 234788
rect 42454 234199 42506 234205
rect 42454 234141 42506 234147
rect 43138 234057 43166 236564
rect 42454 234051 42506 234057
rect 42454 233993 42506 233999
rect 43126 234051 43178 234057
rect 43126 233993 43178 233999
rect 42192 230644 42398 230672
rect 42466 230006 42494 233993
rect 42192 229978 42494 230006
rect 41780 229798 41836 229807
rect 41780 229733 41836 229742
rect 41794 229357 41822 229733
rect 41780 229058 41836 229067
rect 41780 228993 41836 229002
rect 41794 228808 41822 228993
rect 41780 227282 41836 227291
rect 41780 227217 41836 227226
rect 41794 226958 41822 227217
rect 41780 226838 41836 226847
rect 41780 226773 41836 226782
rect 41794 226321 41822 226773
rect 41780 225950 41836 225959
rect 41780 225885 41836 225894
rect 41794 225700 41822 225885
rect 42358 221101 42410 221107
rect 42356 221066 42358 221075
rect 42410 221066 42412 221075
rect 42356 221001 42412 221010
rect 42358 220361 42410 220367
rect 42356 220326 42358 220335
rect 42410 220326 42412 220335
rect 42356 220261 42412 220270
rect 42358 219473 42410 219479
rect 42356 219438 42358 219447
rect 42410 219438 42412 219447
rect 42356 219373 42412 219382
rect 43330 216931 43358 260073
rect 43604 259398 43660 259407
rect 43604 259333 43660 259342
rect 43618 255517 43646 259333
rect 43606 255511 43658 255517
rect 43606 255453 43658 255459
rect 43510 242117 43562 242123
rect 43510 242059 43562 242065
rect 43522 234723 43550 242059
rect 43510 234717 43562 234723
rect 43510 234659 43562 234665
rect 43618 227712 43646 255453
rect 43522 227684 43646 227712
rect 43522 227564 43550 227684
rect 43810 227564 43838 261553
rect 44578 252113 44606 889633
rect 44758 805183 44810 805189
rect 44758 805125 44810 805131
rect 44662 418607 44714 418613
rect 44662 418549 44714 418555
rect 44566 252107 44618 252113
rect 44566 252049 44618 252055
rect 44674 252039 44702 418549
rect 44770 252187 44798 805125
rect 44866 800897 44894 985019
rect 44854 800891 44906 800897
rect 44854 800833 44906 800839
rect 44852 762302 44908 762311
rect 44852 762237 44908 762246
rect 44866 252483 44894 762237
rect 44962 757977 44990 985093
rect 44950 757971 45002 757977
rect 44950 757913 45002 757919
rect 44950 718751 45002 718757
rect 44950 718693 45002 718699
rect 44854 252477 44906 252483
rect 44854 252419 44906 252425
rect 44962 252261 44990 718693
rect 45058 717129 45086 985167
rect 45046 717123 45098 717129
rect 45046 717065 45098 717071
rect 45046 675683 45098 675689
rect 45046 675625 45098 675631
rect 45058 252631 45086 675625
rect 45154 671397 45182 985463
rect 50518 985447 50570 985453
rect 50518 985389 50570 985395
rect 47734 985373 47786 985379
rect 47734 985315 47786 985321
rect 47446 913001 47498 913007
rect 47446 912943 47498 912949
rect 45142 671391 45194 671397
rect 45142 671333 45194 671339
rect 45142 632467 45194 632473
rect 45142 632409 45194 632415
rect 45046 252625 45098 252631
rect 45046 252567 45098 252573
rect 45154 252335 45182 632409
rect 45238 589251 45290 589257
rect 45238 589193 45290 589199
rect 45250 252409 45278 589193
rect 45334 546257 45386 546263
rect 45334 546199 45386 546205
rect 45346 252705 45374 546199
rect 45430 455089 45482 455095
rect 45430 455031 45482 455037
rect 45442 393231 45470 455031
rect 45526 440733 45578 440739
rect 45526 440675 45578 440681
rect 45430 393225 45482 393231
rect 45430 393167 45482 393173
rect 45430 375243 45482 375249
rect 45430 375185 45482 375191
rect 45334 252699 45386 252705
rect 45334 252641 45386 252647
rect 45442 252557 45470 375185
rect 45538 349127 45566 440675
rect 47458 410547 47486 912943
rect 47542 812213 47594 812219
rect 47542 812155 47594 812161
rect 47554 779955 47582 812155
rect 47542 779949 47594 779955
rect 47542 779891 47594 779897
rect 47542 743097 47594 743103
rect 47542 743039 47594 743045
rect 47446 410541 47498 410547
rect 47446 410483 47498 410489
rect 45718 383087 45770 383093
rect 45718 383029 45770 383035
rect 45526 349121 45578 349127
rect 45526 349063 45578 349069
rect 45622 332027 45674 332033
rect 45622 331969 45674 331975
rect 45526 311085 45578 311091
rect 45526 311027 45578 311033
rect 45430 252551 45482 252557
rect 45430 252493 45482 252499
rect 45238 252403 45290 252409
rect 45238 252345 45290 252351
rect 45142 252329 45194 252335
rect 45142 252271 45194 252277
rect 44950 252255 45002 252261
rect 44950 252197 45002 252203
rect 44758 252181 44810 252187
rect 44758 252123 44810 252129
rect 44662 252033 44714 252039
rect 44662 251975 44714 251981
rect 44566 250035 44618 250041
rect 44566 249977 44618 249983
rect 43426 227536 43550 227564
rect 43618 227536 43838 227564
rect 43316 216922 43372 216931
rect 43316 216857 43372 216866
rect 43426 216191 43454 227536
rect 43618 217671 43646 227536
rect 43604 217662 43660 217671
rect 43604 217597 43660 217606
rect 43412 216182 43468 216191
rect 43412 216117 43468 216126
rect 41876 213962 41932 213971
rect 41876 213897 41932 213906
rect 37364 210854 37420 210863
rect 37364 210789 37420 210798
rect 37378 200831 37406 210789
rect 41684 206118 41740 206127
rect 41684 206053 41740 206062
rect 37366 200825 37418 200831
rect 37366 200767 37418 200773
rect 41698 197691 41726 206053
rect 41782 200825 41834 200831
rect 41782 200767 41834 200773
rect 41684 197682 41740 197691
rect 41684 197617 41740 197626
rect 41794 197427 41822 200767
rect 41890 198241 41918 213897
rect 41972 209226 42028 209235
rect 41972 209161 42028 209170
rect 41878 198235 41930 198241
rect 41878 198177 41930 198183
rect 41986 197501 42014 209161
rect 42068 208338 42124 208347
rect 42068 208273 42124 208282
rect 42082 201349 42110 208273
rect 42740 208116 42796 208125
rect 42740 208051 42796 208060
rect 42358 204377 42410 204383
rect 42356 204342 42358 204351
rect 42410 204342 42412 204351
rect 42356 204277 42412 204286
rect 42370 202871 42398 204277
rect 42356 202862 42412 202871
rect 42356 202797 42412 202806
rect 42070 201343 42122 201349
rect 42070 201285 42122 201291
rect 42754 198907 42782 208051
rect 43028 207450 43084 207459
rect 43028 207385 43084 207394
rect 43042 204772 43070 207385
rect 43124 205822 43180 205831
rect 43124 205757 43180 205766
rect 42850 204744 43070 204772
rect 42742 198901 42794 198907
rect 42742 198843 42794 198849
rect 42850 198833 42878 204744
rect 43028 204638 43084 204647
rect 43028 204573 43084 204582
rect 42934 201343 42986 201349
rect 42934 201285 42986 201291
rect 42838 198827 42890 198833
rect 42838 198769 42890 198775
rect 42358 198235 42410 198241
rect 42358 198177 42410 198183
rect 41974 197495 42026 197501
rect 41974 197437 42026 197443
rect 41782 197421 41834 197427
rect 41782 197363 41834 197369
rect 41782 197199 41834 197205
rect 41782 197141 41834 197147
rect 41794 196618 41822 197141
rect 42370 195355 42398 198177
rect 42454 197495 42506 197501
rect 42454 197437 42506 197443
rect 42166 195349 42218 195355
rect 42166 195291 42218 195297
rect 42358 195349 42410 195355
rect 42358 195291 42410 195297
rect 42178 194805 42206 195291
rect 42358 195201 42410 195207
rect 42358 195143 42410 195149
rect 42070 194535 42122 194541
rect 42070 194477 42122 194483
rect 42082 194176 42110 194477
rect 42070 193499 42122 193505
rect 42070 193441 42122 193447
rect 42082 192992 42110 193441
rect 42166 192241 42218 192247
rect 42166 192183 42218 192189
rect 42178 191769 42206 192183
rect 42370 191507 42398 195143
rect 42070 191501 42122 191507
rect 42070 191443 42122 191449
rect 42358 191501 42410 191507
rect 42358 191443 42410 191449
rect 42082 191142 42110 191443
rect 42166 191057 42218 191063
rect 42166 190999 42218 191005
rect 42178 190476 42206 190999
rect 41780 190134 41836 190143
rect 41780 190069 41836 190078
rect 41794 189929 41822 190069
rect 42262 189281 42314 189287
rect 42262 189223 42314 189229
rect 41972 189098 42028 189107
rect 41972 189033 42028 189042
rect 41986 188626 42014 189033
rect 41780 188358 41836 188367
rect 41780 188293 41836 188302
rect 41794 188011 41822 188293
rect 41794 187997 42192 188011
rect 41808 187983 42206 187997
rect 42178 187881 42206 187983
rect 42166 187875 42218 187881
rect 42166 187817 42218 187823
rect 42274 187456 42302 189223
rect 42192 187428 42302 187456
rect 42166 187135 42218 187141
rect 42166 187077 42218 187083
rect 42178 186776 42206 187077
rect 42466 186697 42494 197437
rect 42644 195758 42700 195767
rect 42644 195693 42700 195702
rect 42658 189287 42686 195693
rect 42646 189281 42698 189287
rect 42646 189223 42698 189229
rect 42946 188196 42974 201285
rect 43042 192247 43070 204573
rect 43030 192241 43082 192247
rect 43030 192183 43082 192189
rect 43138 191063 43166 205757
rect 44578 204383 44606 249977
rect 45538 219479 45566 311027
rect 45634 252007 45662 331969
rect 45730 307539 45758 383029
rect 45718 307533 45770 307539
rect 45718 307475 45770 307481
rect 45718 296729 45770 296735
rect 45718 296671 45770 296677
rect 45620 251998 45676 252007
rect 45620 251933 45676 251942
rect 45730 221107 45758 296671
rect 45910 289107 45962 289113
rect 45910 289049 45962 289055
rect 45814 282299 45866 282305
rect 45814 282241 45866 282247
rect 45718 221101 45770 221107
rect 45718 221043 45770 221049
rect 45826 220367 45854 282241
rect 45922 252155 45950 289049
rect 47554 281121 47582 743039
rect 47746 627959 47774 985315
rect 50326 927431 50378 927437
rect 50326 927373 50378 927379
rect 50338 907531 50366 927373
rect 50326 907525 50378 907531
rect 50326 907467 50378 907473
rect 50422 884215 50474 884221
rect 50422 884157 50474 884163
rect 50326 855429 50378 855435
rect 50326 855371 50378 855377
rect 47734 627953 47786 627959
rect 47734 627895 47786 627901
rect 47638 627879 47690 627885
rect 47638 627821 47690 627827
rect 47542 281115 47594 281121
rect 47542 281057 47594 281063
rect 46484 274790 46540 274799
rect 46484 274725 46540 274734
rect 46498 274059 46526 274725
rect 46292 274050 46348 274059
rect 46292 273985 46348 273994
rect 46484 274050 46540 274059
rect 46484 273985 46540 273994
rect 46306 273319 46334 273985
rect 46292 273310 46348 273319
rect 46292 273245 46348 273254
rect 45908 252146 45964 252155
rect 45908 252081 45964 252090
rect 45814 220361 45866 220367
rect 45814 220303 45866 220309
rect 45526 219473 45578 219479
rect 45526 219415 45578 219421
rect 44566 204377 44618 204383
rect 44566 204319 44618 204325
rect 43318 198901 43370 198907
rect 43318 198843 43370 198849
rect 43222 198827 43274 198833
rect 43222 198769 43274 198775
rect 43234 195207 43262 198769
rect 43222 195201 43274 195207
rect 43222 195143 43274 195149
rect 43330 193505 43358 198843
rect 47650 194541 47678 627821
rect 50338 367405 50366 855371
rect 50434 823911 50462 884157
rect 50422 823905 50474 823911
rect 50422 823847 50474 823853
rect 50422 757527 50474 757533
rect 50422 757469 50474 757475
rect 50434 736739 50462 757469
rect 50422 736733 50474 736739
rect 50422 736675 50474 736681
rect 50422 728667 50474 728673
rect 50422 728609 50474 728615
rect 50434 692487 50462 728609
rect 50422 692481 50474 692487
rect 50422 692423 50474 692429
rect 50422 685525 50474 685531
rect 50422 685467 50474 685473
rect 50326 367399 50378 367405
rect 50326 367341 50378 367347
rect 50434 237757 50462 685467
rect 50530 584743 50558 985389
rect 59540 973054 59596 973063
rect 59540 972989 59596 972998
rect 59554 970653 59582 972989
rect 53302 970647 53354 970653
rect 53302 970589 53354 970595
rect 59542 970647 59594 970653
rect 59542 970589 59594 970595
rect 53206 941787 53258 941793
rect 53206 941729 53258 941735
rect 53218 908123 53246 941729
rect 53206 908117 53258 908123
rect 53206 908059 53258 908065
rect 53206 898645 53258 898651
rect 53206 898587 53258 898593
rect 50614 829529 50666 829535
rect 50614 829471 50666 829477
rect 50626 780473 50654 829471
rect 53218 822283 53246 898587
rect 53206 822277 53258 822283
rect 53206 822219 53258 822225
rect 53206 797857 53258 797863
rect 53206 797799 53258 797805
rect 50614 780467 50666 780473
rect 50614 780409 50666 780415
rect 51862 649783 51914 649789
rect 51862 649725 51914 649731
rect 51874 644535 51902 649725
rect 51862 644529 51914 644535
rect 51862 644471 51914 644477
rect 51862 607751 51914 607757
rect 51862 607693 51914 607699
rect 51874 601911 51902 607693
rect 51862 601905 51914 601911
rect 51862 601847 51914 601853
rect 50518 584737 50570 584743
rect 50518 584679 50570 584685
rect 50518 563499 50570 563505
rect 50518 563441 50570 563447
rect 50530 543747 50558 563441
rect 50518 543741 50570 543747
rect 50518 543683 50570 543689
rect 50614 512735 50666 512741
rect 50614 512677 50666 512683
rect 50518 469519 50570 469525
rect 50518 469461 50570 469467
rect 50530 393971 50558 469461
rect 50626 436965 50654 512677
rect 50614 436959 50666 436965
rect 50614 436901 50666 436907
rect 50518 393965 50570 393971
rect 50518 393907 50570 393913
rect 50518 368731 50570 368737
rect 50518 368673 50570 368679
rect 50530 306799 50558 368673
rect 53218 324189 53246 797799
rect 53314 541527 53342 970589
rect 61858 962259 61886 999375
rect 74722 997335 74750 999375
rect 74708 997326 74764 997335
rect 74708 997261 74764 997270
rect 74900 997326 74956 997335
rect 74900 997261 74956 997270
rect 74914 995739 74942 997261
rect 92386 995961 92414 1005221
rect 92578 996151 92606 1005295
rect 92950 999433 93002 999439
rect 92950 999375 93002 999381
rect 92564 996142 92620 996151
rect 92564 996077 92620 996086
rect 92374 995955 92426 995961
rect 92374 995897 92426 995903
rect 92470 995955 92522 995961
rect 92470 995897 92522 995903
rect 78644 995846 78700 995855
rect 78384 995804 78644 995832
rect 80784 995813 81086 995832
rect 84528 995813 84830 995832
rect 91248 995813 91550 995832
rect 80784 995807 81098 995813
rect 80784 995804 81046 995807
rect 78644 995781 78700 995790
rect 84528 995807 84842 995813
rect 84528 995804 84790 995807
rect 81046 995749 81098 995755
rect 91248 995807 91562 995813
rect 91248 995804 91510 995807
rect 84790 995749 84842 995755
rect 91510 995749 91562 995755
rect 74902 995733 74954 995739
rect 74902 995675 74954 995681
rect 82486 995733 82538 995739
rect 85366 995733 85418 995739
rect 82486 995675 82538 995681
rect 85104 995681 85366 995684
rect 89684 995698 89740 995707
rect 85104 995675 85418 995681
rect 82498 995536 82526 995675
rect 85104 995656 85406 995675
rect 89424 995656 89684 995684
rect 89684 995633 89740 995642
rect 77088 995508 77342 995536
rect 77314 993741 77342 995508
rect 77698 993815 77726 995522
rect 77686 993809 77738 993815
rect 80194 993783 80222 995522
rect 81408 995508 81662 995536
rect 82032 995517 82334 995536
rect 82498 995522 82608 995536
rect 82032 995511 82346 995517
rect 82032 995508 82294 995511
rect 81634 995443 81662 995508
rect 82498 995508 82622 995522
rect 83232 995508 83486 995536
rect 82294 995453 82346 995459
rect 81622 995437 81674 995443
rect 81622 995379 81674 995385
rect 82594 994111 82622 995508
rect 82582 994105 82634 994111
rect 82582 994047 82634 994053
rect 77686 993751 77738 993757
rect 80180 993774 80236 993783
rect 77302 993735 77354 993741
rect 80180 993709 80236 993718
rect 77302 993677 77354 993683
rect 83458 993635 83486 995508
rect 85714 995369 85742 995522
rect 86352 995508 86558 995536
rect 87552 995508 87902 995536
rect 86530 995411 86558 995508
rect 86516 995402 86572 995411
rect 85702 995363 85754 995369
rect 86516 995337 86572 995346
rect 85702 995305 85754 995311
rect 87874 995263 87902 995508
rect 87860 995254 87916 995263
rect 87860 995189 87916 995198
rect 88738 993931 88766 995522
rect 92482 995369 92510 995897
rect 92470 995363 92522 995369
rect 92470 995305 92522 995311
rect 88724 993922 88780 993931
rect 88724 993857 88780 993866
rect 92962 993635 92990 999375
rect 62036 993626 62092 993635
rect 62036 993561 62092 993570
rect 83444 993626 83500 993635
rect 83444 993561 83500 993570
rect 92948 993626 93004 993635
rect 92948 993561 93004 993570
rect 61844 962250 61900 962259
rect 61844 962185 61900 962194
rect 62050 962111 62078 993561
rect 93634 986415 93662 1005443
rect 93718 1005427 93770 1005433
rect 93718 1005369 93770 1005375
rect 73366 986409 73418 986415
rect 73366 986351 73418 986357
rect 93622 986409 93674 986415
rect 93622 986351 93674 986357
rect 63286 985521 63338 985527
rect 63286 985463 63338 985469
rect 63298 985305 63326 985463
rect 63286 985299 63338 985305
rect 63286 985241 63338 985247
rect 65206 983893 65258 983899
rect 65206 983835 65258 983841
rect 65110 983597 65162 983603
rect 65110 983539 65162 983545
rect 65014 983523 65066 983529
rect 65014 983465 65066 983471
rect 64918 980859 64970 980865
rect 64918 980801 64970 980807
rect 64822 980785 64874 980791
rect 64822 980727 64874 980733
rect 64630 980711 64682 980717
rect 64630 980653 64682 980659
rect 62036 962102 62092 962111
rect 62036 962037 62092 962046
rect 59348 958698 59404 958707
rect 59348 958633 59404 958642
rect 59362 956223 59390 958633
rect 59350 956217 59402 956223
rect 59350 956159 59402 956165
rect 59540 944342 59596 944351
rect 59540 944277 59596 944286
rect 59554 941793 59582 944277
rect 59542 941787 59594 941793
rect 59542 941729 59594 941735
rect 59540 929986 59596 929995
rect 59540 929921 59596 929930
rect 59554 927437 59582 929921
rect 59542 927431 59594 927437
rect 59542 927373 59594 927379
rect 59540 915482 59596 915491
rect 59540 915417 59596 915426
rect 59554 913007 59582 915417
rect 59542 913001 59594 913007
rect 59542 912943 59594 912949
rect 59540 901274 59596 901283
rect 59540 901209 59596 901218
rect 59554 898651 59582 901209
rect 59542 898645 59594 898651
rect 59542 898587 59594 898593
rect 59540 886770 59596 886779
rect 59540 886705 59596 886714
rect 59554 884221 59582 886705
rect 59542 884215 59594 884221
rect 59542 884157 59594 884163
rect 58964 872414 59020 872423
rect 58964 872349 59020 872358
rect 53398 840999 53450 841005
rect 53398 840941 53450 840947
rect 53410 778919 53438 840941
rect 58198 829529 58250 829535
rect 58196 829494 58198 829503
rect 58250 829494 58252 829503
rect 58196 829429 58252 829438
rect 58978 821913 59006 872349
rect 59540 858058 59596 858067
rect 59540 857993 59596 858002
rect 59554 855435 59582 857993
rect 59542 855429 59594 855435
rect 59542 855371 59594 855377
rect 59540 843702 59596 843711
rect 59540 843637 59596 843646
rect 59554 841005 59582 843637
rect 59542 840999 59594 841005
rect 59542 840941 59594 840947
rect 58966 821907 59018 821913
rect 58966 821849 59018 821855
rect 59540 814990 59596 814999
rect 59540 814925 59596 814934
rect 59554 812219 59582 814925
rect 59542 812213 59594 812219
rect 59542 812155 59594 812161
rect 59540 800634 59596 800643
rect 59540 800569 59596 800578
rect 59554 797863 59582 800569
rect 59542 797857 59594 797863
rect 59542 797799 59594 797805
rect 58964 786278 59020 786287
rect 58964 786213 59020 786222
rect 53398 778913 53450 778919
rect 53398 778855 53450 778861
rect 53398 771883 53450 771889
rect 53398 771825 53450 771831
rect 53410 737257 53438 771825
rect 58196 757566 58252 757575
rect 58196 757501 58198 757510
rect 58250 757501 58252 757510
rect 58198 757469 58250 757475
rect 58580 743210 58636 743219
rect 58580 743145 58636 743154
rect 58594 743103 58622 743145
rect 58582 743097 58634 743103
rect 58582 743039 58634 743045
rect 53398 737251 53450 737257
rect 53398 737193 53450 737199
rect 58978 735481 59006 786213
rect 59540 771922 59596 771931
rect 59540 771857 59542 771866
rect 59594 771857 59596 771866
rect 59542 771825 59594 771831
rect 58966 735475 59018 735481
rect 58966 735417 59018 735423
rect 59540 728854 59596 728863
rect 59540 728789 59596 728798
rect 59554 728673 59582 728789
rect 59542 728667 59594 728673
rect 59542 728609 59594 728615
rect 59540 714350 59596 714359
rect 53398 714311 53450 714317
rect 59540 714285 59542 714294
rect 53398 714253 53450 714259
rect 59594 714285 59596 714294
rect 59542 714253 59594 714259
rect 53410 694041 53438 714253
rect 59540 700142 59596 700151
rect 59540 700077 59596 700086
rect 59554 699887 59582 700077
rect 59542 699881 59594 699887
rect 59542 699823 59594 699829
rect 53398 694035 53450 694041
rect 53398 693977 53450 693983
rect 58676 685638 58732 685647
rect 58676 685573 58732 685582
rect 58690 685531 58718 685573
rect 58678 685525 58730 685531
rect 58678 685467 58730 685473
rect 58388 671430 58444 671439
rect 58388 671365 58444 671374
rect 58402 671101 58430 671365
rect 53398 671095 53450 671101
rect 53398 671037 53450 671043
rect 58390 671095 58442 671101
rect 58390 671037 58442 671043
rect 53410 649567 53438 671037
rect 59540 656926 59596 656935
rect 59540 656861 59596 656870
rect 59554 656745 59582 656861
rect 59542 656739 59594 656745
rect 59542 656681 59594 656687
rect 53398 649561 53450 649567
rect 53398 649503 53450 649509
rect 59542 644529 59594 644535
rect 59542 644471 59594 644477
rect 59554 642727 59582 644471
rect 59540 642718 59596 642727
rect 59540 642653 59596 642662
rect 58388 628214 58444 628223
rect 58388 628149 58444 628158
rect 58402 627885 58430 628149
rect 58390 627879 58442 627885
rect 58390 627821 58442 627827
rect 58388 613858 58444 613867
rect 58388 613793 58444 613802
rect 58402 613529 58430 613793
rect 58390 613523 58442 613529
rect 58390 613465 58442 613471
rect 53398 606863 53450 606869
rect 53398 606805 53450 606811
rect 53410 587481 53438 606805
rect 59542 601905 59594 601911
rect 59542 601847 59594 601853
rect 59554 599511 59582 601847
rect 59540 599502 59596 599511
rect 59540 599437 59596 599446
rect 53398 587475 53450 587481
rect 53398 587417 53450 587423
rect 59542 587475 59594 587481
rect 59542 587417 59594 587423
rect 59554 585303 59582 587417
rect 59540 585294 59596 585303
rect 59540 585229 59596 585238
rect 59540 570790 59596 570799
rect 59540 570725 59596 570734
rect 59554 570313 59582 570725
rect 59542 570307 59594 570313
rect 59542 570249 59594 570255
rect 53398 564535 53450 564541
rect 53398 564477 53450 564483
rect 53410 558695 53438 564477
rect 53398 558689 53450 558695
rect 53398 558631 53450 558637
rect 59542 558689 59594 558695
rect 59542 558631 59594 558637
rect 59554 556591 59582 558631
rect 59540 556582 59596 556591
rect 59540 556517 59596 556526
rect 59542 543741 59594 543747
rect 59542 543683 59594 543689
rect 59554 542235 59582 543683
rect 59540 542226 59596 542235
rect 59540 542161 59596 542170
rect 53302 541521 53354 541527
rect 53302 541463 53354 541469
rect 59444 527574 59500 527583
rect 59444 527509 59500 527518
rect 59458 527097 59486 527509
rect 59446 527091 59498 527097
rect 59446 527033 59498 527039
rect 59540 513366 59596 513375
rect 59540 513301 59596 513310
rect 59554 512741 59582 513301
rect 59542 512735 59594 512741
rect 59542 512677 59594 512683
rect 58100 499010 58156 499019
rect 58100 498945 58156 498954
rect 58114 498311 58142 498945
rect 53398 498305 53450 498311
rect 53398 498247 53450 498253
rect 58102 498305 58154 498311
rect 58102 498247 58154 498253
rect 53302 483875 53354 483881
rect 53302 483817 53354 483823
rect 53314 392343 53342 483817
rect 53410 436151 53438 498247
rect 59540 484506 59596 484515
rect 59540 484441 59596 484450
rect 59554 483881 59582 484441
rect 59542 483875 59594 483881
rect 59542 483817 59594 483823
rect 59540 470298 59596 470307
rect 59540 470233 59596 470242
rect 59554 469525 59582 470233
rect 59542 469519 59594 469525
rect 59542 469461 59594 469467
rect 59540 455794 59596 455803
rect 59540 455729 59596 455738
rect 59554 455095 59582 455729
rect 59542 455089 59594 455095
rect 59542 455031 59594 455037
rect 59540 441438 59596 441447
rect 59540 441373 59596 441382
rect 59554 440739 59582 441373
rect 59542 440733 59594 440739
rect 59542 440675 59594 440681
rect 53398 436145 53450 436151
rect 53398 436087 53450 436093
rect 59348 427082 59404 427091
rect 59348 427017 59404 427026
rect 59362 426309 59390 427017
rect 53398 426303 53450 426309
rect 53398 426245 53450 426251
rect 59350 426303 59402 426309
rect 59350 426245 59402 426251
rect 53302 392337 53354 392343
rect 53302 392279 53354 392285
rect 53410 350755 53438 426245
rect 57812 412726 57868 412735
rect 57812 412661 57868 412670
rect 57826 411879 57854 412661
rect 53494 411873 53546 411879
rect 53494 411815 53546 411821
rect 57814 411873 57866 411879
rect 57814 411815 57866 411821
rect 53398 350749 53450 350755
rect 53398 350691 53450 350697
rect 53506 349719 53534 411815
rect 59060 398370 59116 398379
rect 59060 398305 59116 398314
rect 58964 355302 59020 355311
rect 58964 355237 59020 355246
rect 53494 349713 53546 349719
rect 53494 349655 53546 349661
rect 53302 339871 53354 339877
rect 53302 339813 53354 339819
rect 53206 324183 53258 324189
rect 53206 324125 53258 324131
rect 50518 306793 50570 306799
rect 50518 306735 50570 306741
rect 53314 264323 53342 339813
rect 53398 325515 53450 325521
rect 53398 325457 53450 325463
rect 53302 264317 53354 264323
rect 53302 264259 53354 264265
rect 53410 263583 53438 325457
rect 57620 283522 57676 283531
rect 57620 283457 57676 283466
rect 57634 282305 57662 283457
rect 57622 282299 57674 282305
rect 57622 282241 57674 282247
rect 53398 263577 53450 263583
rect 53398 263519 53450 263525
rect 58978 262325 59006 355237
rect 59074 305541 59102 398305
rect 59540 384014 59596 384023
rect 59540 383949 59596 383958
rect 59554 383093 59582 383949
rect 59542 383087 59594 383093
rect 59542 383029 59594 383035
rect 59540 369658 59596 369667
rect 59540 369593 59596 369602
rect 59554 368737 59582 369593
rect 59542 368731 59594 368737
rect 59542 368673 59594 368679
rect 59540 340946 59596 340955
rect 59540 340881 59596 340890
rect 59554 339877 59582 340881
rect 59542 339871 59594 339877
rect 59542 339813 59594 339819
rect 59540 326442 59596 326451
rect 59540 326377 59596 326386
rect 59554 325521 59582 326377
rect 59542 325515 59594 325521
rect 59542 325457 59594 325463
rect 59540 312234 59596 312243
rect 59540 312169 59596 312178
rect 59554 311091 59582 312169
rect 59542 311085 59594 311091
rect 59542 311027 59594 311033
rect 59062 305535 59114 305541
rect 59062 305477 59114 305483
rect 59540 297730 59596 297739
rect 59540 297665 59596 297674
rect 59554 296735 59582 297665
rect 59542 296729 59594 296735
rect 59542 296671 59594 296677
rect 64642 275201 64670 980653
rect 64726 980637 64778 980643
rect 64726 980579 64778 980585
rect 64630 275195 64682 275201
rect 64630 275137 64682 275143
rect 64738 275127 64766 980579
rect 64726 275121 64778 275127
rect 64726 275063 64778 275069
rect 64834 273499 64862 980727
rect 64822 273493 64874 273499
rect 64822 273435 64874 273441
rect 64930 270983 64958 980801
rect 64918 270977 64970 270983
rect 64918 270919 64970 270925
rect 58966 262319 59018 262325
rect 58966 262261 59018 262267
rect 60598 255585 60650 255591
rect 60598 255527 60650 255533
rect 60502 255511 60554 255517
rect 60502 255453 60554 255459
rect 60514 255388 60542 255453
rect 60610 255388 60638 255527
rect 60514 255360 60638 255388
rect 65026 254967 65054 983465
rect 65012 254958 65068 254967
rect 65012 254893 65068 254902
rect 65122 254819 65150 983539
rect 65218 254925 65246 983835
rect 73378 981314 73406 986351
rect 93730 985897 93758 1005369
rect 95074 995855 95102 1005517
rect 100726 1005501 100778 1005507
rect 108694 1005501 108746 1005507
rect 100726 1005443 100778 1005449
rect 108692 1005466 108694 1005475
rect 433270 1005501 433322 1005507
rect 108746 1005466 108748 1005475
rect 100738 1004989 100766 1005443
rect 108692 1005401 108748 1005410
rect 115220 1005466 115276 1005475
rect 115220 1005401 115222 1005410
rect 115274 1005401 115276 1005410
rect 321044 1005466 321100 1005475
rect 321428 1005466 321484 1005475
rect 321100 1005424 321428 1005452
rect 321044 1005401 321100 1005410
rect 321428 1005401 321484 1005410
rect 325460 1005466 325516 1005475
rect 325460 1005401 325516 1005410
rect 358676 1005466 358732 1005475
rect 431636 1005466 431692 1005475
rect 358676 1005401 358678 1005410
rect 115222 1005369 115274 1005375
rect 109462 1005353 109514 1005359
rect 106580 1005318 106636 1005327
rect 106580 1005253 106582 1005262
rect 106634 1005253 106636 1005262
rect 109460 1005318 109462 1005327
rect 298294 1005353 298346 1005359
rect 109514 1005318 109516 1005327
rect 109460 1005253 109516 1005262
rect 217268 1005318 217324 1005327
rect 217268 1005253 217270 1005262
rect 106582 1005221 106634 1005227
rect 217322 1005253 217324 1005262
rect 218900 1005318 218956 1005327
rect 218900 1005253 218902 1005262
rect 217270 1005221 217322 1005227
rect 218954 1005253 218956 1005262
rect 223124 1005318 223180 1005327
rect 308758 1005353 308810 1005359
rect 298294 1005295 298346 1005301
rect 308756 1005318 308758 1005327
rect 308810 1005318 308812 1005327
rect 223124 1005253 223180 1005262
rect 218902 1005221 218954 1005227
rect 198742 1005205 198794 1005211
rect 114164 1005170 114220 1005179
rect 207286 1005205 207338 1005211
rect 198742 1005147 198794 1005153
rect 207284 1005170 207286 1005179
rect 207338 1005170 207340 1005179
rect 114164 1005105 114220 1005114
rect 114178 1004989 114206 1005105
rect 100726 1004983 100778 1004989
rect 100726 1004925 100778 1004931
rect 114166 1004983 114218 1004989
rect 114166 1004925 114218 1004931
rect 195286 1003725 195338 1003731
rect 195286 1003667 195338 1003673
rect 151508 1002654 151564 1002663
rect 144214 1002615 144266 1002621
rect 151508 1002589 151510 1002598
rect 144214 1002557 144266 1002563
rect 151562 1002589 151564 1002598
rect 151510 1002557 151562 1002563
rect 143734 1002541 143786 1002547
rect 143734 1002483 143786 1002489
rect 143746 999532 143774 1002483
rect 143926 1002467 143978 1002473
rect 143926 1002409 143978 1002415
rect 143830 1000839 143882 1000845
rect 143830 1000781 143882 1000787
rect 143650 999504 143774 999532
rect 123862 999433 123914 999439
rect 123862 999375 123914 999381
rect 103894 996029 103946 996035
rect 101492 995994 101548 996003
rect 101492 995929 101494 995938
rect 101546 995929 101548 995938
rect 103892 995994 103894 996003
rect 115222 996029 115274 996035
rect 103946 995994 103948 996003
rect 106964 995994 107020 996003
rect 103892 995929 103948 995938
rect 106486 995955 106538 995961
rect 101494 995897 101546 995903
rect 106964 995929 107020 995938
rect 113396 995994 113452 996003
rect 115222 995971 115274 995977
rect 113396 995929 113398 995938
rect 106486 995897 106538 995903
rect 95060 995846 95116 995855
rect 95060 995781 95116 995790
rect 99764 995846 99820 995855
rect 99764 995781 99820 995790
rect 105428 995846 105484 995855
rect 105428 995781 105430 995790
rect 99778 995739 99806 995781
rect 105482 995781 105484 995790
rect 105430 995749 105482 995755
rect 99766 995733 99818 995739
rect 94964 995698 95020 995707
rect 94964 995633 95020 995642
rect 98900 995698 98956 995707
rect 98900 995633 98956 995642
rect 99668 995698 99724 995707
rect 99766 995675 99818 995681
rect 103124 995698 103180 995707
rect 99668 995633 99724 995642
rect 103124 995633 103180 995642
rect 89590 985891 89642 985897
rect 89590 985833 89642 985839
rect 93718 985891 93770 985897
rect 93718 985833 93770 985839
rect 89602 981314 89630 985833
rect 90646 985817 90698 985823
rect 90646 985759 90698 985765
rect 90658 985305 90686 985759
rect 90646 985299 90698 985305
rect 90646 985241 90698 985247
rect 94978 983899 95006 995633
rect 98914 995411 98942 995633
rect 99682 995517 99710 995633
rect 99670 995511 99722 995517
rect 99670 995453 99722 995459
rect 103138 995443 103166 995633
rect 103126 995437 103178 995443
rect 98900 995402 98956 995411
rect 103126 995379 103178 995385
rect 98900 995337 98956 995346
rect 100724 995106 100780 995115
rect 100724 995041 100780 995050
rect 100738 993815 100766 995041
rect 100726 993809 100778 993815
rect 100726 993751 100778 993757
rect 94966 983893 95018 983899
rect 94966 983835 95018 983841
rect 106498 981476 106526 995897
rect 106978 993783 107006 995929
rect 113450 995929 113452 995938
rect 113398 995897 113450 995903
rect 113396 995846 113452 995855
rect 113396 995781 113398 995790
rect 113450 995781 113452 995790
rect 113398 995749 113450 995755
rect 115234 995707 115262 995971
rect 123874 995855 123902 999375
rect 123860 995846 123916 995855
rect 118102 995807 118154 995813
rect 134516 995846 134572 995855
rect 132144 995813 132446 995832
rect 132144 995807 132458 995813
rect 132144 995804 132406 995807
rect 123860 995781 123916 995790
rect 118102 995749 118154 995755
rect 136724 995846 136780 995855
rect 134572 995818 134640 995832
rect 134572 995804 134654 995818
rect 136464 995804 136724 995832
rect 134516 995781 134572 995790
rect 132406 995749 132458 995755
rect 115220 995698 115276 995707
rect 115220 995633 115276 995642
rect 108212 995550 108268 995559
rect 108212 995485 108268 995494
rect 115316 995550 115372 995559
rect 115316 995485 115372 995494
rect 106964 993774 107020 993783
rect 108226 993741 108254 995485
rect 115220 995402 115276 995411
rect 115220 995337 115276 995346
rect 106964 993709 107020 993718
rect 108214 993735 108266 993741
rect 108214 993677 108266 993683
rect 115234 993445 115262 995337
rect 115330 993519 115358 995485
rect 115318 993513 115370 993519
rect 115318 993455 115370 993461
rect 115222 993439 115274 993445
rect 115222 993381 115274 993387
rect 115234 983751 115262 993381
rect 115330 983825 115358 993455
rect 115318 983819 115370 983825
rect 115318 983761 115370 983767
rect 115222 983745 115274 983751
rect 115222 983687 115274 983693
rect 118114 983677 118142 995749
rect 132816 995665 133118 995684
rect 132816 995659 133130 995665
rect 132816 995656 133078 995659
rect 133078 995601 133130 995607
rect 128482 993741 128510 995522
rect 129120 995508 129374 995536
rect 129346 995443 129374 995508
rect 129334 995437 129386 995443
rect 129334 995379 129386 995385
rect 129730 994227 129758 995522
rect 131616 995508 131870 995536
rect 129716 994218 129772 994227
rect 129716 994153 129772 994162
rect 131842 993815 131870 995508
rect 133426 995295 133454 995522
rect 134002 995369 134030 995522
rect 133990 995363 134042 995369
rect 133990 995305 134042 995311
rect 133414 995289 133466 995295
rect 134002 995240 134030 995305
rect 133414 995231 133466 995237
rect 133954 995212 134030 995240
rect 133954 994111 133982 995212
rect 133942 994105 133994 994111
rect 134626 994079 134654 995804
rect 137972 995846 138028 995855
rect 137760 995804 137972 995832
rect 136724 995781 136780 995790
rect 142656 995813 143006 995832
rect 142656 995807 143018 995813
rect 142656 995804 142966 995807
rect 137972 995781 138028 995790
rect 142966 995749 143018 995755
rect 141046 995733 141098 995739
rect 137396 995698 137452 995707
rect 137136 995656 137396 995684
rect 140784 995681 141046 995684
rect 143650 995707 143678 999504
rect 143734 999433 143786 999439
rect 143734 999375 143786 999381
rect 143746 995813 143774 999375
rect 143734 995807 143786 995813
rect 143734 995749 143786 995755
rect 143842 995739 143870 1000781
rect 143830 995733 143882 995739
rect 140784 995675 141098 995681
rect 143636 995698 143692 995707
rect 140784 995656 141086 995675
rect 137396 995633 137452 995642
rect 143830 995675 143882 995681
rect 143636 995633 143692 995642
rect 143938 995591 143966 1002409
rect 144022 1002393 144074 1002399
rect 144022 1002335 144074 1002341
rect 144034 995855 144062 1002335
rect 144118 999507 144170 999513
rect 144118 999449 144170 999455
rect 144130 995961 144158 999449
rect 144226 996003 144254 1002557
rect 152854 1002541 152906 1002547
rect 152852 1002506 152854 1002515
rect 152906 1002506 152908 1002515
rect 152852 1002441 152908 1002450
rect 153620 1002506 153676 1002515
rect 153620 1002441 153622 1002450
rect 153674 1002441 153676 1002450
rect 153622 1002409 153674 1002415
rect 150358 1002393 150410 1002399
rect 150356 1002358 150358 1002367
rect 150410 1002358 150412 1002367
rect 144310 1002319 144362 1002325
rect 150356 1002293 150412 1002302
rect 178486 1002319 178538 1002325
rect 144310 1002261 144362 1002267
rect 178486 1002261 178538 1002267
rect 144212 995994 144268 996003
rect 144118 995955 144170 995961
rect 144212 995929 144268 995938
rect 144118 995897 144170 995903
rect 144020 995846 144076 995855
rect 144020 995781 144076 995790
rect 139318 995585 139370 995591
rect 135936 995508 136190 995536
rect 138960 995533 139318 995536
rect 143926 995585 143978 995591
rect 138960 995527 139370 995533
rect 138960 995508 139358 995527
rect 140160 995508 140414 995536
rect 143926 995527 143978 995533
rect 136162 994375 136190 995508
rect 136148 994366 136204 994375
rect 136148 994301 136204 994310
rect 133942 994047 133994 994053
rect 134612 994070 134668 994079
rect 134612 994005 134668 994014
rect 131830 993809 131882 993815
rect 140386 993783 140414 995508
rect 144322 995369 144350 1002261
rect 160244 1000878 160300 1000887
rect 160244 1000813 160246 1000822
rect 160298 1000813 160300 1000822
rect 160246 1000781 160298 1000787
rect 155156 999546 155212 999555
rect 155156 999481 155158 999490
rect 155210 999481 155212 999490
rect 155158 999449 155210 999455
rect 156886 999433 156938 999439
rect 156884 999398 156886 999407
rect 156938 999398 156940 999407
rect 156884 999333 156940 999342
rect 162646 996177 162698 996183
rect 162646 996119 162698 996125
rect 164084 996142 164140 996151
rect 145268 995994 145324 996003
rect 144406 995955 144458 995961
rect 145268 995929 145324 995938
rect 149108 995994 149164 996003
rect 149492 995994 149548 996003
rect 149164 995952 149492 995980
rect 149108 995929 149164 995938
rect 149492 995929 149548 995938
rect 151988 995994 152044 996003
rect 151988 995929 151990 995938
rect 144406 995897 144458 995903
rect 144310 995363 144362 995369
rect 144310 995305 144362 995311
rect 144418 995295 144446 995897
rect 144406 995289 144458 995295
rect 144406 995231 144458 995237
rect 131830 993751 131882 993757
rect 140372 993774 140428 993783
rect 128470 993735 128522 993741
rect 140372 993709 140428 993718
rect 128470 993677 128522 993683
rect 126742 993513 126794 993519
rect 126742 993455 126794 993461
rect 126754 993371 126782 993455
rect 126742 993365 126794 993371
rect 126742 993307 126794 993313
rect 138262 986409 138314 986415
rect 138262 986351 138314 986357
rect 122038 985447 122090 985453
rect 122038 985389 122090 985395
rect 118102 983671 118154 983677
rect 118102 983613 118154 983619
rect 106114 981448 106526 981476
rect 106114 981328 106142 981448
rect 105840 981300 106142 981328
rect 122050 981314 122078 985389
rect 138274 981314 138302 986351
rect 145282 983603 145310 995929
rect 152042 995929 152044 995938
rect 159476 995994 159532 996003
rect 159476 995929 159532 995938
rect 151990 995897 152042 995903
rect 158612 995846 158668 995855
rect 158612 995781 158668 995790
rect 146804 995698 146860 995707
rect 146804 995633 146806 995642
rect 146858 995633 146860 995642
rect 158324 995698 158380 995707
rect 158324 995633 158380 995642
rect 146806 995601 146858 995607
rect 146804 995550 146860 995559
rect 146804 995485 146860 995494
rect 146818 995443 146846 995485
rect 146806 995437 146858 995443
rect 146806 995379 146858 995385
rect 158338 994227 158366 995633
rect 158324 994218 158380 994227
rect 158324 994153 158380 994162
rect 158626 993815 158654 995781
rect 158614 993809 158666 993815
rect 158614 993751 158666 993757
rect 159490 993741 159518 995929
rect 162658 995559 162686 996119
rect 164084 996077 164086 996086
rect 164138 996077 164140 996086
rect 164086 996045 164138 996051
rect 164182 996029 164234 996035
rect 164180 995994 164182 996003
rect 164234 995994 164236 996003
rect 164180 995929 164236 995938
rect 178498 995855 178526 1002261
rect 195094 1000913 195146 1000919
rect 195094 1000855 195146 1000861
rect 165620 995846 165676 995855
rect 164086 995807 164138 995813
rect 165620 995781 165622 995790
rect 164086 995749 164138 995755
rect 165674 995781 165676 995790
rect 166196 995846 166252 995855
rect 166196 995781 166252 995790
rect 178484 995846 178540 995855
rect 178484 995781 178540 995790
rect 185204 995846 185260 995855
rect 187604 995846 187660 995855
rect 185260 995818 185424 995832
rect 185260 995804 185438 995818
rect 187344 995804 187604 995832
rect 185204 995781 185260 995790
rect 165622 995749 165674 995755
rect 163990 995733 164042 995739
rect 162932 995698 162988 995707
rect 163990 995675 164042 995681
rect 162932 995633 162988 995642
rect 162644 995550 162700 995559
rect 162644 995485 162700 995494
rect 159478 993735 159530 993741
rect 159478 993677 159530 993683
rect 162658 993445 162686 995485
rect 162946 993519 162974 995633
rect 162934 993513 162986 993519
rect 162934 993455 162986 993461
rect 162646 993439 162698 993445
rect 162646 993381 162698 993387
rect 164002 986785 164030 995675
rect 154486 986779 154538 986785
rect 154486 986721 154538 986727
rect 163990 986779 164042 986785
rect 163990 986721 164042 986727
rect 145270 983597 145322 983603
rect 145270 983539 145322 983545
rect 154498 981314 154526 986721
rect 164098 986415 164126 995749
rect 166210 995739 166238 995781
rect 166198 995733 166250 995739
rect 166198 995675 166250 995681
rect 170228 995698 170284 995707
rect 170228 995633 170284 995642
rect 164086 986409 164138 986415
rect 164086 986351 164138 986357
rect 170242 983992 170270 995633
rect 185108 995550 185164 995559
rect 179842 993667 179870 995522
rect 180514 993889 180542 995522
rect 181152 995508 181406 995536
rect 180502 993883 180554 993889
rect 180502 993825 180554 993831
rect 181378 993741 181406 995508
rect 183010 993815 183038 995522
rect 183552 995508 183806 995536
rect 184176 995517 184382 995536
rect 184176 995511 184394 995517
rect 184176 995508 184342 995511
rect 183778 995443 183806 995508
rect 184848 995508 185108 995536
rect 185108 995485 185164 995494
rect 184342 995453 184394 995459
rect 183766 995437 183818 995443
rect 183766 995379 183818 995385
rect 185410 994227 185438 995804
rect 192500 995846 192556 995855
rect 187872 995813 188126 995832
rect 187872 995807 188138 995813
rect 187872 995804 188086 995807
rect 187604 995781 187660 995790
rect 192192 995804 192500 995832
rect 192500 995781 192556 995790
rect 188086 995749 188138 995755
rect 188854 995733 188906 995739
rect 188544 995681 188854 995684
rect 189428 995698 189484 995707
rect 188544 995675 188906 995681
rect 188544 995656 188894 995675
rect 189168 995656 189428 995684
rect 194064 995665 194462 995684
rect 195106 995665 195134 1000855
rect 195190 999433 195242 999439
rect 195190 999375 195242 999381
rect 194064 995659 194474 995665
rect 194064 995656 194422 995659
rect 189428 995633 189484 995642
rect 194422 995601 194474 995607
rect 195094 995659 195146 995665
rect 195094 995601 195146 995607
rect 195202 995591 195230 999375
rect 195298 995855 195326 1003667
rect 195382 997953 195434 997959
rect 195382 997895 195434 997901
rect 195394 996003 195422 997895
rect 195380 995994 195436 996003
rect 195380 995929 195436 995938
rect 195670 995955 195722 995961
rect 195670 995897 195722 995903
rect 195284 995846 195340 995855
rect 195284 995781 195340 995790
rect 191926 995585 191978 995591
rect 190580 995550 190636 995559
rect 185986 995508 186048 995536
rect 190368 995508 190580 995536
rect 185396 994218 185452 994227
rect 185396 994153 185452 994162
rect 185986 994079 186014 995508
rect 191568 995533 191926 995536
rect 191568 995527 191978 995533
rect 195190 995585 195242 995591
rect 195190 995527 195242 995533
rect 191568 995508 191966 995527
rect 190580 995485 190636 995494
rect 185972 994070 186028 994079
rect 185972 994005 186028 994014
rect 182998 993809 183050 993815
rect 182998 993751 183050 993757
rect 181366 993735 181418 993741
rect 181366 993677 181418 993683
rect 179830 993661 179882 993667
rect 179830 993603 179882 993609
rect 181462 985521 181514 985527
rect 181460 985486 181462 985495
rect 181514 985486 181516 985495
rect 181460 985421 181516 985430
rect 187316 985486 187372 985495
rect 187316 985421 187372 985430
rect 187330 985379 187358 985421
rect 186934 985373 186986 985379
rect 186934 985315 186986 985321
rect 187318 985373 187370 985379
rect 187318 985315 187370 985321
rect 170242 983964 170462 983992
rect 170434 981328 170462 983964
rect 170434 981300 170736 981328
rect 186946 981314 186974 985315
rect 195682 983529 195710 995897
rect 198754 993889 198782 1005147
rect 207284 1005105 207340 1005114
rect 221876 1005170 221932 1005179
rect 221876 1005105 221932 1005114
rect 211702 1003725 211754 1003731
rect 211700 1003690 211702 1003699
rect 211754 1003690 211756 1003699
rect 211700 1003625 211756 1003634
rect 208150 1000913 208202 1000919
rect 208148 1000878 208150 1000887
rect 208202 1000878 208204 1000887
rect 208148 1000813 208204 1000822
rect 209398 997953 209450 997959
rect 209396 997918 209398 997927
rect 209450 997918 209452 997927
rect 209396 997853 209452 997862
rect 213334 996177 213386 996183
rect 213332 996142 213334 996151
rect 213386 996142 213388 996151
rect 213332 996077 213388 996086
rect 215636 996142 215692 996151
rect 215636 996077 215638 996086
rect 215690 996077 215692 996086
rect 218902 996103 218954 996109
rect 215638 996045 215690 996051
rect 218902 996045 218954 996051
rect 200276 995994 200332 996003
rect 200276 995929 200278 995938
rect 200330 995929 200332 995938
rect 200948 995994 201004 996003
rect 200948 995929 200950 995938
rect 200278 995897 200330 995903
rect 201002 995929 201004 995938
rect 204212 995994 204268 996003
rect 204212 995929 204268 995938
rect 206612 995994 206668 996003
rect 216788 995994 216844 996003
rect 206612 995929 206668 995938
rect 213046 995955 213098 995961
rect 200950 995897 201002 995903
rect 202868 995846 202924 995855
rect 202868 995781 202870 995790
rect 202922 995781 202924 995790
rect 203348 995846 203404 995855
rect 203348 995781 203404 995790
rect 202870 995749 202922 995755
rect 201526 995511 201578 995517
rect 201526 995453 201578 995459
rect 201538 995263 201566 995453
rect 203362 995411 203390 995781
rect 204226 995739 204254 995929
rect 204214 995733 204266 995739
rect 204214 995675 204266 995681
rect 206626 995443 206654 995929
rect 216788 995929 216790 995938
rect 213046 995897 213098 995903
rect 216842 995929 216844 995938
rect 216790 995897 216842 995903
rect 206614 995437 206666 995443
rect 203348 995402 203404 995411
rect 206614 995379 206666 995385
rect 212660 995402 212716 995411
rect 203348 995337 203404 995346
rect 212660 995337 212716 995346
rect 201524 995254 201580 995263
rect 201524 995189 201580 995198
rect 210164 995254 210220 995263
rect 210164 995189 210220 995198
rect 211028 995254 211084 995263
rect 211028 995189 211084 995198
rect 198742 993883 198794 993889
rect 198742 993825 198794 993831
rect 210178 993815 210206 995189
rect 210166 993809 210218 993815
rect 210166 993751 210218 993757
rect 211042 993667 211070 995189
rect 212674 993741 212702 995337
rect 212662 993735 212714 993741
rect 212662 993677 212714 993683
rect 211030 993661 211082 993667
rect 211030 993603 211082 993609
rect 213058 986341 213086 995897
rect 218914 995707 218942 996045
rect 218900 995698 218956 995707
rect 218900 995633 218956 995642
rect 214388 995402 214444 995411
rect 214388 995337 214444 995346
rect 214402 993593 214430 995337
rect 214390 993587 214442 993593
rect 214390 993529 214442 993535
rect 221890 987155 221918 1005105
rect 223138 987821 223166 1005253
rect 298198 1000395 298250 1000401
rect 298198 1000337 298250 1000343
rect 246646 999581 246698 999587
rect 260758 999581 260810 999587
rect 246646 999523 246698 999529
rect 258836 999546 258892 999555
rect 226006 999433 226058 999439
rect 226006 999375 226058 999381
rect 246550 999433 246602 999439
rect 246550 999375 246602 999381
rect 226018 995073 226046 999375
rect 246454 995955 246506 995961
rect 246454 995897 246506 995903
rect 238868 995846 238924 995855
rect 236256 995813 236510 995832
rect 236256 995807 236522 995813
rect 236256 995804 236470 995807
rect 238704 995804 238868 995832
rect 239540 995846 239596 995855
rect 239280 995804 239540 995832
rect 238868 995781 238924 995790
rect 245424 995813 245726 995832
rect 245424 995807 245738 995813
rect 245424 995804 245686 995807
rect 239540 995781 239596 995790
rect 236470 995749 236522 995755
rect 245686 995749 245738 995755
rect 240212 995698 240268 995707
rect 239952 995656 240212 995684
rect 240212 995633 240268 995642
rect 240788 995550 240844 995559
rect 231264 995508 231518 995536
rect 231936 995508 232190 995536
rect 226006 995067 226058 995073
rect 226006 995009 226058 995015
rect 227542 994475 227594 994481
rect 227542 994417 227594 994423
rect 227554 994227 227582 994417
rect 231490 994375 231518 995508
rect 231476 994366 231532 994375
rect 231476 994301 231532 994310
rect 227540 994218 227596 994227
rect 227540 994153 227596 994162
rect 232162 993815 232190 995508
rect 232150 993809 232202 993815
rect 232150 993751 232202 993757
rect 232546 993741 232574 995522
rect 234370 994523 234398 995522
rect 234356 994514 234412 994523
rect 234356 994449 234412 994458
rect 234946 993889 234974 995522
rect 235584 995508 235838 995536
rect 235810 993963 235838 995508
rect 236770 994481 236798 995522
rect 236758 994475 236810 994481
rect 236758 994417 236810 994423
rect 237442 994079 237470 995522
rect 240576 995508 240788 995536
rect 241776 995508 241886 995536
rect 242976 995508 243230 995536
rect 240788 995485 240844 995494
rect 241858 995411 241886 995508
rect 241844 995402 241900 995411
rect 241844 995337 241900 995346
rect 238966 994475 239018 994481
rect 238966 994417 239018 994423
rect 237428 994070 237484 994079
rect 237428 994005 237484 994014
rect 235798 993957 235850 993963
rect 235798 993899 235850 993905
rect 234934 993883 234986 993889
rect 234934 993825 234986 993831
rect 232534 993735 232586 993741
rect 232534 993677 232586 993683
rect 238978 993667 239006 994417
rect 243202 994079 243230 995508
rect 243586 994671 243614 995522
rect 243572 994662 243628 994671
rect 243572 994597 243628 994606
rect 243188 994070 243244 994079
rect 243094 994031 243146 994037
rect 243188 994005 243244 994014
rect 243094 993973 243146 993979
rect 243106 993815 243134 993973
rect 246466 993963 246494 995897
rect 246562 995813 246590 999375
rect 246658 996003 246686 999523
rect 247702 999507 247754 999513
rect 258836 999481 258838 999490
rect 247702 999449 247754 999455
rect 258890 999481 258892 999490
rect 260756 999546 260758 999555
rect 260810 999546 260812 999555
rect 260756 999481 260812 999490
rect 258838 999449 258890 999455
rect 246644 995994 246700 996003
rect 246644 995929 246700 995938
rect 247604 995994 247660 996003
rect 247604 995929 247660 995938
rect 246550 995807 246602 995813
rect 246550 995749 246602 995755
rect 246454 993957 246506 993963
rect 246454 993899 246506 993905
rect 243094 993809 243146 993815
rect 243094 993751 243146 993757
rect 247618 993741 247646 995929
rect 247714 994037 247742 999449
rect 259606 999433 259658 999439
rect 259604 999398 259606 999407
rect 298102 999433 298154 999439
rect 259658 999398 259660 999407
rect 298102 999375 298154 999381
rect 259604 999333 259660 999342
rect 263924 996586 263980 996595
rect 259126 996547 259178 996553
rect 263924 996521 263926 996530
rect 259126 996489 259178 996495
rect 263978 996521 263980 996530
rect 263926 996489 263978 996495
rect 254902 995881 254954 995887
rect 250484 995846 250540 995855
rect 250484 995781 250486 995790
rect 250538 995781 250540 995790
rect 254036 995846 254092 995855
rect 254036 995781 254038 995790
rect 250486 995749 250538 995755
rect 254090 995781 254092 995790
rect 254900 995846 254902 995855
rect 257302 995881 257354 995887
rect 254954 995846 254956 995855
rect 254900 995781 254956 995790
rect 255668 995846 255724 995855
rect 255668 995781 255724 995790
rect 257300 995846 257302 995855
rect 257354 995846 257356 995855
rect 257300 995781 257356 995790
rect 254038 995749 254090 995755
rect 255682 995739 255710 995781
rect 250390 995733 250442 995739
rect 250388 995698 250390 995707
rect 255670 995733 255722 995739
rect 250442 995698 250444 995707
rect 255670 995675 255722 995681
rect 250388 995633 250444 995642
rect 250484 995106 250540 995115
rect 250484 995041 250540 995050
rect 250498 994185 250526 995041
rect 247798 994179 247850 994185
rect 247798 994121 247850 994127
rect 250486 994179 250538 994185
rect 250486 994121 250538 994127
rect 247702 994031 247754 994037
rect 247702 993973 247754 993979
rect 247810 993908 247838 994121
rect 259138 994111 259166 996489
rect 265078 996177 265130 996183
rect 265076 996142 265078 996151
rect 276502 996177 276554 996183
rect 265130 996142 265132 996151
rect 266996 996142 267052 996151
rect 265076 996077 265132 996086
rect 266902 996103 266954 996109
rect 276502 996119 276554 996125
rect 266996 996077 266998 996086
rect 266902 996045 266954 996051
rect 267050 996077 267052 996086
rect 266998 996045 267050 996051
rect 266914 996003 266942 996045
rect 276514 996035 276542 996119
rect 276502 996029 276554 996035
rect 266900 995994 266956 996003
rect 276502 995971 276554 995977
rect 266900 995929 266956 995938
rect 262676 995846 262732 995855
rect 262676 995781 262732 995790
rect 268532 995846 268588 995855
rect 268532 995781 268534 995790
rect 262690 994671 262718 995781
rect 268586 995781 268588 995790
rect 273620 995846 273676 995855
rect 292532 995846 292588 995855
rect 290880 995813 291230 995832
rect 273620 995781 273676 995790
rect 273718 995807 273770 995813
rect 268534 995749 268586 995755
rect 265748 995698 265804 995707
rect 265748 995633 265804 995642
rect 268052 995698 268108 995707
rect 268052 995633 268108 995642
rect 262676 994662 262732 994671
rect 262676 994597 262732 994606
rect 259126 994105 259178 994111
rect 259126 994047 259178 994053
rect 247714 993889 247838 993908
rect 247702 993883 247838 993889
rect 247754 993880 247838 993883
rect 247702 993825 247754 993831
rect 243286 993735 243338 993741
rect 243286 993677 243338 993683
rect 247606 993735 247658 993741
rect 247606 993677 247658 993683
rect 238966 993661 239018 993667
rect 238966 993603 239018 993609
rect 223126 987815 223178 987821
rect 223126 987757 223178 987763
rect 235606 987815 235658 987821
rect 235606 987757 235658 987763
rect 219382 987149 219434 987155
rect 219382 987091 219434 987097
rect 221878 987149 221930 987155
rect 221878 987091 221930 987097
rect 203158 986335 203210 986341
rect 203158 986277 203210 986283
rect 213046 986335 213098 986341
rect 213046 986277 213098 986283
rect 195670 983523 195722 983529
rect 195670 983465 195722 983471
rect 203170 981314 203198 986277
rect 219394 981314 219422 987091
rect 235618 981314 235646 987757
rect 243298 980865 243326 993677
rect 265762 993593 265790 995633
rect 265750 993587 265802 993593
rect 265750 993529 265802 993535
rect 251734 985299 251786 985305
rect 251734 985241 251786 985247
rect 251746 981314 251774 985241
rect 268066 981314 268094 995633
rect 273634 986489 273662 995781
rect 290880 995807 291242 995813
rect 290880 995804 291190 995807
rect 273718 995749 273770 995755
rect 292176 995804 292532 995832
rect 292532 995781 292588 995790
rect 291190 995749 291242 995755
rect 273622 986483 273674 986489
rect 273622 986425 273674 986431
rect 273730 986415 273758 995749
rect 298114 995739 298142 999375
rect 297334 995733 297386 995739
rect 295412 995698 295468 995707
rect 287184 995665 287486 995684
rect 291504 995665 291806 995684
rect 287184 995659 287498 995665
rect 287184 995656 287446 995659
rect 291504 995659 291818 995665
rect 291504 995656 291766 995659
rect 287446 995601 287498 995607
rect 295200 995656 295412 995684
rect 297072 995681 297334 995684
rect 297072 995675 297386 995681
rect 298102 995733 298154 995739
rect 298210 995707 298238 1000337
rect 298306 995887 298334 1005295
rect 299542 1005279 299594 1005285
rect 308756 1005253 308812 1005262
rect 309620 1005318 309676 1005327
rect 309620 1005253 309622 1005262
rect 299542 1005221 299594 1005227
rect 309674 1005253 309676 1005262
rect 309622 1005221 309674 1005227
rect 298294 995881 298346 995887
rect 299446 995881 299498 995887
rect 298294 995823 298346 995829
rect 299444 995846 299446 995855
rect 299498 995846 299500 995855
rect 299444 995781 299500 995790
rect 298102 995675 298154 995681
rect 298196 995698 298252 995707
rect 297072 995656 297374 995675
rect 295412 995633 295468 995642
rect 298196 995633 298252 995642
rect 298484 995698 298540 995707
rect 298484 995633 298540 995642
rect 291766 995601 291818 995607
rect 287926 995585 287978 995591
rect 286772 995550 286828 995559
rect 282850 993667 282878 995522
rect 283522 993741 283550 995522
rect 284160 995508 284414 995536
rect 286032 995508 286334 995536
rect 286560 995508 286772 995536
rect 284386 994523 284414 995508
rect 286306 994671 286334 995508
rect 287856 995533 287926 995536
rect 287856 995527 287978 995533
rect 287856 995508 287966 995527
rect 288384 995508 288446 995536
rect 286772 995485 286828 995494
rect 286292 994662 286348 994671
rect 286292 994597 286348 994606
rect 284372 994514 284428 994523
rect 284372 994449 284428 994458
rect 283510 993735 283562 993741
rect 283510 993677 283562 993683
rect 279286 993661 279338 993667
rect 279284 993626 279286 993635
rect 282838 993661 282890 993667
rect 279338 993626 279340 993635
rect 288418 993635 288446 995508
rect 288994 995508 289056 995536
rect 288994 994227 289022 995508
rect 290338 994819 290366 995522
rect 293376 995508 293630 995536
rect 293602 995411 293630 995508
rect 293588 995402 293644 995411
rect 293588 995337 293644 995346
rect 290324 994810 290380 994819
rect 290324 994745 290380 994754
rect 294562 994227 294590 995522
rect 288980 994218 289036 994227
rect 288980 994153 289036 994162
rect 294548 994218 294604 994227
rect 294548 994153 294604 994162
rect 282838 993603 282890 993609
rect 288404 993626 288460 993635
rect 279284 993561 279340 993570
rect 288404 993561 288460 993570
rect 284278 986483 284330 986489
rect 284278 986425 284330 986431
rect 273718 986409 273770 986415
rect 273718 986351 273770 986357
rect 284290 981314 284318 986425
rect 243286 980859 243338 980865
rect 243286 980801 243338 980807
rect 298498 980791 298526 995633
rect 299554 995559 299582 1005221
rect 325474 1005211 325502 1005401
rect 358730 1005401 358732 1005410
rect 379126 1005427 379178 1005433
rect 358678 1005369 358730 1005375
rect 431636 1005401 431638 1005410
rect 379126 1005369 379178 1005375
rect 431690 1005401 431692 1005410
rect 433268 1005466 433270 1005475
rect 433322 1005466 433324 1005475
rect 433268 1005401 433324 1005410
rect 431638 1005369 431690 1005375
rect 365014 1005353 365066 1005359
rect 365012 1005318 365014 1005327
rect 365066 1005318 365068 1005327
rect 365012 1005253 365068 1005262
rect 305302 1005205 305354 1005211
rect 314230 1005205 314282 1005211
rect 305302 1005147 305354 1005153
rect 314228 1005170 314230 1005179
rect 325462 1005205 325514 1005211
rect 314282 1005170 314284 1005179
rect 305314 1000401 305342 1005147
rect 325462 1005147 325514 1005153
rect 331222 1005205 331274 1005211
rect 358006 1005205 358058 1005211
rect 331222 1005147 331274 1005153
rect 358004 1005170 358006 1005179
rect 358058 1005170 358060 1005179
rect 314228 1005105 314284 1005114
rect 305302 1000395 305354 1000401
rect 305302 1000337 305354 1000343
rect 311254 999433 311306 999439
rect 311252 999398 311254 999407
rect 311306 999398 311308 999407
rect 311252 999333 311308 999342
rect 328342 997953 328394 997959
rect 328342 997895 328394 997901
rect 325462 997879 325514 997885
rect 325462 997821 325514 997827
rect 318454 997805 318506 997811
rect 318452 997770 318454 997779
rect 318506 997770 318508 997779
rect 318452 997705 318508 997714
rect 316342 996473 316394 996479
rect 316342 996415 316394 996421
rect 316354 996183 316382 996415
rect 302326 996177 302378 996183
rect 316342 996177 316394 996183
rect 302326 996119 302378 996125
rect 316340 996142 316342 996151
rect 316394 996142 316396 996151
rect 302338 995647 302366 996119
rect 316340 996077 316396 996086
rect 318644 996142 318700 996151
rect 318644 996077 318646 996086
rect 318698 996077 318700 996086
rect 318646 996045 318698 996051
rect 305684 995994 305740 996003
rect 305684 995929 305740 995938
rect 313844 995994 313900 996003
rect 313844 995929 313900 995938
rect 304726 995881 304778 995887
rect 304724 995846 304726 995855
rect 304778 995846 304780 995855
rect 305698 995813 305726 995929
rect 307316 995846 307372 995855
rect 304724 995781 304780 995790
rect 305686 995807 305738 995813
rect 307316 995781 307372 995790
rect 310292 995846 310348 995855
rect 310292 995781 310294 995790
rect 305686 995749 305738 995755
rect 302422 995733 302474 995739
rect 302422 995675 302474 995681
rect 302242 995619 302366 995647
rect 299540 995550 299596 995559
rect 302242 995517 302270 995619
rect 302326 995585 302378 995591
rect 302324 995550 302326 995559
rect 302378 995550 302380 995559
rect 299540 995485 299596 995494
rect 302230 995511 302282 995517
rect 302324 995485 302380 995494
rect 302230 995453 302282 995459
rect 302434 993741 302462 995675
rect 307330 995665 307358 995781
rect 310346 995781 310348 995790
rect 310294 995749 310346 995755
rect 309236 995698 309292 995707
rect 307318 995659 307370 995665
rect 309236 995633 309292 995642
rect 313364 995698 313420 995707
rect 313364 995633 313420 995642
rect 307318 995601 307370 995607
rect 309250 994819 309278 995633
rect 309236 994810 309292 994819
rect 309236 994745 309292 994754
rect 313378 994523 313406 995633
rect 313364 994514 313420 994523
rect 313364 994449 313420 994458
rect 302422 993735 302474 993741
rect 302422 993677 302474 993683
rect 313858 993667 313886 995929
rect 317492 995846 317548 995855
rect 317492 995781 317548 995790
rect 313846 993661 313898 993667
rect 313846 993603 313898 993609
rect 317506 993593 317534 995781
rect 323924 995698 323980 995707
rect 323924 995633 323980 995642
rect 320758 994771 320810 994777
rect 320758 994713 320810 994719
rect 317494 993587 317546 993593
rect 317494 993529 317546 993535
rect 320770 986489 320798 994713
rect 316918 986483 316970 986489
rect 316918 986425 316970 986431
rect 320758 986483 320810 986489
rect 320758 986425 320810 986431
rect 300406 986409 300458 986415
rect 300406 986351 300458 986357
rect 300418 981314 300446 986351
rect 316726 985225 316778 985231
rect 316726 985167 316778 985173
rect 316738 981314 316766 985167
rect 298486 980785 298538 980791
rect 298486 980727 298538 980733
rect 316930 980717 316958 986425
rect 323938 986415 323966 995633
rect 325474 994777 325502 997821
rect 326804 995994 326860 996003
rect 326804 995929 326860 995938
rect 325462 994771 325514 994777
rect 325462 994713 325514 994719
rect 326818 986489 326846 995929
rect 328354 993593 328382 997895
rect 328342 993587 328394 993593
rect 328342 993529 328394 993535
rect 331234 992187 331262 1005147
rect 358004 1005105 358060 1005114
rect 356756 1003986 356812 1003995
rect 356756 1003921 356758 1003930
rect 356810 1003921 356812 1003930
rect 377206 1003947 377258 1003953
rect 356758 1003889 356810 1003895
rect 377206 1003889 377258 1003895
rect 359062 1003873 359114 1003879
rect 355988 1003838 356044 1003847
rect 355988 1003773 355990 1003782
rect 356042 1003773 356044 1003782
rect 359060 1003838 359062 1003847
rect 359114 1003838 359116 1003847
rect 359060 1003773 359116 1003782
rect 377110 1003799 377162 1003805
rect 355990 1003741 356042 1003747
rect 377110 1003741 377162 1003747
rect 359926 1003725 359978 1003731
rect 359924 1003690 359926 1003699
rect 359978 1003690 359980 1003699
rect 359924 1003625 359980 1003634
rect 361556 1000878 361612 1000887
rect 361556 1000813 361558 1000822
rect 361610 1000813 361612 1000822
rect 361558 1000781 361610 1000787
rect 377122 999439 377150 1003741
rect 377110 999433 377162 999439
rect 377110 999375 377162 999381
rect 367894 997953 367946 997959
rect 367892 997918 367894 997927
rect 371446 997953 371498 997959
rect 367946 997918 367948 997927
rect 350134 997879 350186 997885
rect 371446 997895 371498 997901
rect 367892 997853 367948 997862
rect 350134 997821 350186 997827
rect 350146 995855 350174 997821
rect 369046 997805 369098 997811
rect 369044 997770 369046 997779
rect 369098 997770 369100 997779
rect 369044 997705 369100 997714
rect 367124 996142 367180 996151
rect 367124 996077 367126 996086
rect 367178 996077 367180 996086
rect 367126 996045 367178 996051
rect 362324 995994 362380 996003
rect 362324 995929 362380 995938
rect 370196 995994 370252 996003
rect 370196 995929 370198 995938
rect 350132 995846 350188 995855
rect 350132 995781 350188 995790
rect 360980 995846 361036 995855
rect 360980 995781 360982 995790
rect 361034 995781 361036 995790
rect 360982 995749 361034 995755
rect 362338 993667 362366 995929
rect 370250 995929 370252 995938
rect 370198 995897 370250 995903
rect 368854 995881 368906 995887
rect 365876 995846 365932 995855
rect 365782 995807 365834 995813
rect 368854 995823 368906 995829
rect 365876 995781 365932 995790
rect 365782 995749 365834 995755
rect 365794 994523 365822 995749
rect 365890 995739 365918 995781
rect 365878 995733 365930 995739
rect 368866 995707 368894 995823
rect 371458 995813 371486 997895
rect 377218 997145 377246 1003889
rect 379138 999661 379166 1005369
rect 383638 1005353 383690 1005359
rect 425302 1005353 425354 1005359
rect 383638 1005295 383690 1005301
rect 424532 1005318 424588 1005327
rect 383542 1005205 383594 1005211
rect 383542 1005147 383594 1005153
rect 379990 1003873 380042 1003879
rect 379990 1003815 380042 1003821
rect 379126 999655 379178 999661
rect 379126 999597 379178 999603
rect 379030 999433 379082 999439
rect 379030 999375 379082 999381
rect 377206 997139 377258 997145
rect 377206 997081 377258 997087
rect 377492 995994 377548 996003
rect 374518 995955 374570 995961
rect 377492 995929 377548 995938
rect 374518 995897 374570 995903
rect 371446 995807 371498 995813
rect 371446 995749 371498 995755
rect 365878 995675 365930 995681
rect 368852 995698 368908 995707
rect 368852 995633 368908 995642
rect 374420 995698 374476 995707
rect 374420 995633 374476 995642
rect 365780 994514 365836 994523
rect 365780 994449 365836 994458
rect 362326 993661 362378 993667
rect 362326 993603 362378 993609
rect 331222 992181 331274 992187
rect 331222 992123 331274 992129
rect 332566 992181 332618 992187
rect 332566 992123 332618 992129
rect 326806 986483 326858 986489
rect 326806 986425 326858 986431
rect 323926 986409 323978 986415
rect 323926 986351 323978 986357
rect 332578 981328 332606 992123
rect 374434 986563 374462 995633
rect 374422 986557 374474 986563
rect 374422 986499 374474 986505
rect 349078 986483 349130 986489
rect 349078 986425 349130 986431
rect 332578 981300 332976 981328
rect 349090 981314 349118 986425
rect 374530 986415 374558 995897
rect 377300 995846 377356 995855
rect 377300 995781 377356 995790
rect 377314 995739 377342 995781
rect 377302 995733 377354 995739
rect 377302 995675 377354 995681
rect 377506 986489 377534 995929
rect 379042 994967 379070 999375
rect 380002 996553 380030 1003815
rect 380086 1003725 380138 1003731
rect 380086 1003667 380138 1003673
rect 380098 996572 380126 1003667
rect 381430 999655 381482 999661
rect 381430 999597 381482 999603
rect 379990 996547 380042 996553
rect 380098 996544 380222 996572
rect 379990 996489 380042 996495
rect 380194 995855 380222 996544
rect 380278 996547 380330 996553
rect 380278 996489 380330 996495
rect 380290 996151 380318 996489
rect 380276 996142 380332 996151
rect 380276 996077 380332 996086
rect 380180 995846 380236 995855
rect 380180 995781 380236 995790
rect 381442 995707 381470 999597
rect 382006 997139 382058 997145
rect 382006 997081 382058 997087
rect 381428 995698 381484 995707
rect 381428 995633 381484 995642
rect 382018 995115 382046 997081
rect 383554 995887 383582 1005147
rect 383650 1001012 383678 1005295
rect 424532 1005253 424534 1005262
rect 424586 1005253 424588 1005262
rect 425300 1005318 425302 1005327
rect 434710 1005353 434762 1005359
rect 425354 1005318 425356 1005327
rect 434806 1005353 434858 1005359
rect 434710 1005295 434762 1005301
rect 434804 1005318 434806 1005327
rect 434858 1005318 434860 1005327
rect 425300 1005253 425356 1005262
rect 424534 1005221 424586 1005227
rect 426070 1005205 426122 1005211
rect 426068 1005170 426070 1005179
rect 426122 1005170 426124 1005179
rect 426068 1005105 426124 1005114
rect 434722 1005063 434750 1005295
rect 434804 1005253 434860 1005262
rect 435572 1005170 435628 1005179
rect 435572 1005105 435574 1005114
rect 435626 1005105 435628 1005114
rect 435574 1005073 435626 1005079
rect 437218 1005063 437246 1005517
rect 440566 1005501 440618 1005507
rect 440566 1005443 440618 1005449
rect 441622 1005501 441674 1005507
rect 443446 1005501 443498 1005507
rect 441674 1005449 441854 1005452
rect 441622 1005443 441854 1005449
rect 443446 1005443 443498 1005449
rect 440578 1005359 440606 1005443
rect 441634 1005433 441854 1005443
rect 441634 1005427 441866 1005433
rect 441634 1005424 441814 1005427
rect 441814 1005369 441866 1005375
rect 437782 1005353 437834 1005359
rect 440566 1005353 440618 1005359
rect 437782 1005295 437834 1005301
rect 438740 1005318 438796 1005327
rect 434710 1005057 434762 1005063
rect 434710 1004999 434762 1005005
rect 437206 1005057 437258 1005063
rect 437206 1004999 437258 1005005
rect 428086 1003873 428138 1003879
rect 423380 1003838 423436 1003847
rect 423380 1003773 423382 1003782
rect 423434 1003773 423436 1003782
rect 428084 1003838 428086 1003847
rect 428138 1003838 428140 1003847
rect 428084 1003773 428140 1003782
rect 423382 1003741 423434 1003747
rect 426454 1003725 426506 1003731
rect 426452 1003690 426454 1003699
rect 426506 1003690 426508 1003699
rect 426452 1003625 426508 1003634
rect 434036 1001174 434092 1001183
rect 434036 1001109 434038 1001118
rect 434090 1001109 434092 1001118
rect 434038 1001077 434090 1001083
rect 432502 1001061 432554 1001067
rect 430868 1001026 430924 1001035
rect 383650 1000984 383774 1001012
rect 383638 1000839 383690 1000845
rect 383638 1000781 383690 1000787
rect 383542 995881 383594 995887
rect 383542 995823 383594 995829
rect 383650 995813 383678 1000781
rect 383638 995807 383690 995813
rect 383638 995749 383690 995755
rect 383746 995739 383774 1000984
rect 430868 1000961 430870 1000970
rect 430922 1000961 430924 1000970
rect 432500 1001026 432502 1001035
rect 432554 1001026 432556 1001035
rect 432500 1000961 432556 1000970
rect 430870 1000929 430922 1000935
rect 428950 1000913 429002 1000919
rect 427316 1000878 427372 1000887
rect 427316 1000813 427318 1000822
rect 427370 1000813 427372 1000822
rect 428948 1000878 428950 1000887
rect 429002 1000878 429004 1000887
rect 428948 1000813 429004 1000822
rect 427318 1000781 427370 1000787
rect 423286 996399 423338 996405
rect 423286 996341 423338 996347
rect 423298 996183 423326 996341
rect 399862 996177 399914 996183
rect 399862 996119 399914 996125
rect 408886 996177 408938 996183
rect 408982 996177 409034 996183
rect 408938 996125 408982 996128
rect 408886 996119 409034 996125
rect 423286 996177 423338 996183
rect 436438 996177 436490 996183
rect 423286 996119 423338 996125
rect 436436 996142 436438 996151
rect 436490 996142 436492 996151
rect 399874 995961 399902 996119
rect 408898 996100 409022 996119
rect 437794 996109 437822 1005295
rect 439700 1005318 439756 1005327
rect 438796 1005276 439700 1005304
rect 438740 1005253 438796 1005262
rect 440566 1005295 440618 1005301
rect 440866 1005285 441086 1005304
rect 439700 1005253 439756 1005262
rect 440854 1005279 441098 1005285
rect 440906 1005276 441046 1005279
rect 440854 1005221 440906 1005227
rect 441046 1005221 441098 1005227
rect 443458 1005211 443486 1005443
rect 444884 1005318 444940 1005327
rect 444884 1005253 444940 1005262
rect 443446 1005205 443498 1005211
rect 443446 1005147 443498 1005153
rect 440758 1005131 440810 1005137
rect 440758 1005073 440810 1005079
rect 440770 996405 440798 1005073
rect 440758 996399 440810 996405
rect 440758 996341 440810 996347
rect 436436 996077 436492 996086
rect 437782 996103 437834 996109
rect 437782 996045 437834 996051
rect 436438 996029 436490 996035
rect 429716 995994 429772 996003
rect 399862 995955 399914 995961
rect 429716 995929 429772 995938
rect 436436 995994 436438 996003
rect 436490 995994 436492 996003
rect 436436 995929 436492 995938
rect 399862 995897 399914 995903
rect 388820 995846 388876 995855
rect 384994 995813 385296 995832
rect 384982 995807 385296 995813
rect 385034 995804 385296 995807
rect 396692 995846 396748 995855
rect 389410 995813 389664 995832
rect 388820 995781 388876 995790
rect 389398 995807 389664 995813
rect 384982 995749 385034 995755
rect 383734 995733 383786 995739
rect 383734 995675 383786 995681
rect 384406 995733 384458 995739
rect 388834 995684 388862 995781
rect 389450 995804 389664 995807
rect 396748 995804 397008 995832
rect 396692 995781 396748 995790
rect 389398 995749 389450 995755
rect 393044 995698 393100 995707
rect 384458 995681 384672 995684
rect 384406 995675 384672 995681
rect 384418 995656 384672 995675
rect 388834 995656 388992 995684
rect 410324 995698 410380 995707
rect 393100 995656 393312 995684
rect 393044 995633 393100 995642
rect 410324 995633 410380 995642
rect 385844 995550 385900 995559
rect 394868 995550 394924 995559
rect 385900 995508 385968 995536
rect 387490 995508 387792 995536
rect 385844 995485 385900 995494
rect 387490 995411 387518 995508
rect 387476 995402 387532 995411
rect 387476 995337 387532 995346
rect 382004 995106 382060 995115
rect 382004 995041 382060 995050
rect 379028 994958 379084 994967
rect 379028 994893 379084 994902
rect 388354 994523 388382 995522
rect 388340 994514 388396 994523
rect 388340 994449 388396 994458
rect 390178 993635 390206 995522
rect 390864 995508 391166 995536
rect 391138 994523 391166 995508
rect 392098 995263 392126 995522
rect 392084 995254 392140 995263
rect 392084 995189 392140 995198
rect 392674 995115 392702 995522
rect 393730 995508 393984 995536
rect 392660 995106 392716 995115
rect 392660 995041 392716 995050
rect 393730 994967 393758 995508
rect 394924 995508 395184 995536
rect 394868 995485 394924 995494
rect 393716 994958 393772 994967
rect 393716 994893 393772 994902
rect 391124 994514 391180 994523
rect 391124 994449 391180 994458
rect 396322 994375 396350 995522
rect 396308 994366 396364 994375
rect 396308 994301 396364 994310
rect 398818 993667 398846 995522
rect 398806 993661 398858 993667
rect 390164 993626 390220 993635
rect 398806 993603 398858 993609
rect 390164 993561 390220 993570
rect 390178 992155 390206 993561
rect 390164 992146 390220 992155
rect 390164 992081 390220 992090
rect 397750 986557 397802 986563
rect 397750 986499 397802 986505
rect 377494 986483 377546 986489
rect 377494 986425 377546 986431
rect 365398 986409 365450 986415
rect 365398 986351 365450 986357
rect 374518 986409 374570 986415
rect 374518 986351 374570 986357
rect 365410 981314 365438 986351
rect 381622 985151 381674 985157
rect 381622 985093 381674 985099
rect 381634 981314 381662 985093
rect 397762 981314 397790 986499
rect 316918 980711 316970 980717
rect 316918 980653 316970 980659
rect 410338 980643 410366 995633
rect 429730 993667 429758 995929
rect 440660 995698 440716 995707
rect 440660 995633 440716 995642
rect 429718 993661 429770 993667
rect 429718 993603 429770 993609
rect 414070 986483 414122 986489
rect 414070 986425 414122 986431
rect 414082 981314 414110 986425
rect 440674 986415 440702 995633
rect 430294 986409 430346 986415
rect 430294 986351 430346 986357
rect 440662 986409 440714 986415
rect 440662 986351 440714 986357
rect 430306 981314 430334 986351
rect 444898 985157 444926 1005253
rect 447778 1005211 447806 1005665
rect 469174 1005649 469226 1005655
rect 469174 1005591 469226 1005597
rect 466486 1005575 466538 1005581
rect 466486 1005517 466538 1005523
rect 452950 1005353 453002 1005359
rect 452950 1005295 453002 1005301
rect 447766 1005205 447818 1005211
rect 445076 1005170 445132 1005179
rect 447766 1005147 447818 1005153
rect 445076 1005105 445132 1005114
rect 445090 986489 445118 1005105
rect 452962 1002103 452990 1005295
rect 466498 1005008 466526 1005517
rect 466498 1004980 466622 1005008
rect 466486 1003873 466538 1003879
rect 466486 1003815 466538 1003821
rect 452950 1002097 453002 1002103
rect 452950 1002039 453002 1002045
rect 461590 1002097 461642 1002103
rect 461590 1002039 461642 1002045
rect 461602 998773 461630 1002039
rect 461590 998767 461642 998773
rect 461590 998709 461642 998715
rect 466498 995855 466526 1003815
rect 466594 999439 466622 1004980
rect 469186 1000771 469214 1005591
rect 470998 1005501 471050 1005507
rect 504598 1005501 504650 1005507
rect 470998 1005443 471050 1005449
rect 504596 1005466 504598 1005475
rect 504650 1005466 504652 1005475
rect 469366 1005205 469418 1005211
rect 469366 1005147 469418 1005153
rect 469270 1003799 469322 1003805
rect 469270 1003741 469322 1003747
rect 469174 1000765 469226 1000771
rect 469174 1000707 469226 1000713
rect 466582 999433 466634 999439
rect 466582 999375 466634 999381
rect 469282 998792 469310 1003741
rect 469378 1002103 469406 1005147
rect 470134 1003725 470186 1003731
rect 470134 1003667 470186 1003673
rect 469366 1002097 469418 1002103
rect 469366 1002039 469418 1002045
rect 469558 1000765 469610 1000771
rect 469558 1000707 469610 1000713
rect 466582 998767 466634 998773
rect 469282 998764 469502 998792
rect 466582 998709 466634 998715
rect 466484 995846 466540 995855
rect 466484 995781 466540 995790
rect 466594 995517 466622 998709
rect 466582 995511 466634 995517
rect 466582 995453 466634 995459
rect 469474 995295 469502 998764
rect 469462 995289 469514 995295
rect 469462 995231 469514 995237
rect 469570 994671 469598 1000707
rect 469556 994662 469612 994671
rect 469556 994597 469612 994606
rect 470146 993815 470174 1003667
rect 471010 996035 471038 1005443
rect 471862 1005427 471914 1005433
rect 471862 1005369 471914 1005375
rect 498742 1005427 498794 1005433
rect 504596 1005401 504652 1005410
rect 512662 1005427 512714 1005433
rect 498742 1005369 498794 1005375
rect 512662 1005369 512714 1005375
rect 572854 1005427 572906 1005433
rect 572854 1005369 572906 1005375
rect 471874 996109 471902 1005369
rect 472054 1005279 472106 1005285
rect 472054 1005221 472106 1005227
rect 471862 996103 471914 996109
rect 471862 996045 471914 996051
rect 470998 996029 471050 996035
rect 472066 996003 472094 1005221
rect 498754 1005179 498782 1005369
rect 502292 1005318 502348 1005327
rect 502292 1005253 502294 1005262
rect 502346 1005253 502348 1005262
rect 502294 1005221 502346 1005227
rect 508630 1005205 508682 1005211
rect 498356 1005170 498412 1005179
rect 498740 1005170 498796 1005179
rect 498412 1005128 498740 1005156
rect 498356 1005105 498412 1005114
rect 498740 1005105 498796 1005114
rect 508628 1005170 508630 1005179
rect 508682 1005170 508684 1005179
rect 508628 1005105 508684 1005114
rect 512674 1004915 512702 1005369
rect 554516 1005318 554572 1005327
rect 516790 1005279 516842 1005285
rect 516790 1005221 516842 1005227
rect 521398 1005279 521450 1005285
rect 554516 1005253 554518 1005262
rect 521398 1005221 521450 1005227
rect 554570 1005253 554572 1005262
rect 571894 1005279 571946 1005285
rect 554518 1005221 554570 1005227
rect 571894 1005221 571946 1005227
rect 512662 1004909 512714 1004915
rect 512662 1004851 512714 1004857
rect 501142 1003873 501194 1003879
rect 501140 1003838 501142 1003847
rect 501194 1003838 501196 1003847
rect 501140 1003773 501196 1003782
rect 500374 1003725 500426 1003731
rect 500372 1003690 500374 1003699
rect 500426 1003690 500428 1003699
rect 500372 1003625 500428 1003634
rect 502774 1002541 502826 1002547
rect 502772 1002506 502774 1002515
rect 515446 1002541 515498 1002547
rect 502826 1002506 502828 1002515
rect 489526 1002467 489578 1002473
rect 502772 1002441 502828 1002450
rect 503444 1002506 503500 1002515
rect 515446 1002483 515498 1002489
rect 503444 1002441 503446 1002450
rect 489526 1002409 489578 1002415
rect 503498 1002441 503500 1002450
rect 513526 1002467 513578 1002473
rect 503446 1002409 503498 1002415
rect 513526 1002409 513578 1002415
rect 472150 1002097 472202 1002103
rect 472150 1002039 472202 1002045
rect 470998 995971 471050 995977
rect 472052 995994 472108 996003
rect 472052 995929 472108 995938
rect 472162 995443 472190 1002039
rect 472630 1001135 472682 1001141
rect 472630 1001077 472682 1001083
rect 472534 1001061 472586 1001067
rect 472534 1001003 472586 1001009
rect 472642 1001012 472670 1001077
rect 472342 1000987 472394 1000993
rect 472342 1000929 472394 1000935
rect 472246 999433 472298 999439
rect 472246 999375 472298 999381
rect 472258 995591 472286 999375
rect 472354 995961 472382 1000929
rect 472438 1000839 472490 1000845
rect 472438 1000781 472490 1000787
rect 472342 995955 472394 995961
rect 472342 995897 472394 995903
rect 472450 995887 472478 1000781
rect 472438 995881 472490 995887
rect 472438 995823 472490 995829
rect 472546 995739 472574 1001003
rect 472642 1000984 472766 1001012
rect 472630 1000913 472682 1000919
rect 472630 1000855 472682 1000861
rect 472642 995813 472670 1000855
rect 472630 995807 472682 995813
rect 472630 995749 472682 995755
rect 472534 995733 472586 995739
rect 472534 995675 472586 995681
rect 472738 995665 472766 1000984
rect 488852 999398 488908 999407
rect 488852 999333 488908 999342
rect 477044 995846 477100 995855
rect 474082 995813 474336 995832
rect 474070 995807 474336 995813
rect 474122 995804 474336 995807
rect 481460 995846 481516 995855
rect 477100 995804 477360 995832
rect 477730 995813 477984 995832
rect 480994 995813 481104 995832
rect 477718 995807 477984 995813
rect 477044 995781 477100 995790
rect 474070 995749 474122 995755
rect 477770 995804 477984 995807
rect 480982 995807 481104 995813
rect 477718 995749 477770 995755
rect 481034 995804 481104 995807
rect 481516 995804 481680 995832
rect 481460 995781 481516 995790
rect 480982 995749 481034 995755
rect 473302 995733 473354 995739
rect 488866 995707 488894 999333
rect 480116 995698 480172 995707
rect 473354 995681 473664 995684
rect 473302 995675 473664 995681
rect 472726 995659 472778 995665
rect 473314 995656 473664 995675
rect 474658 995665 474960 995684
rect 479856 995670 480116 995684
rect 474646 995659 474960 995665
rect 472726 995601 472778 995607
rect 474698 995656 474960 995659
rect 479842 995656 480116 995670
rect 474646 995601 474698 995607
rect 472246 995585 472298 995591
rect 472246 995527 472298 995533
rect 476374 995585 476426 995591
rect 476426 995533 476784 995536
rect 476374 995527 476784 995533
rect 476386 995508 476784 995527
rect 478306 995517 478656 995536
rect 478294 995511 478656 995517
rect 478346 995508 478656 995511
rect 478294 995453 478346 995459
rect 472150 995437 472202 995443
rect 472150 995379 472202 995385
rect 470134 993809 470186 993815
rect 470134 993751 470186 993757
rect 469460 993626 469516 993635
rect 479170 993593 479198 995522
rect 479842 994523 479870 995656
rect 480116 995633 480172 995642
rect 488852 995698 488908 995707
rect 488852 995633 488908 995642
rect 482038 995585 482090 995591
rect 482090 995533 482352 995536
rect 482038 995527 482352 995533
rect 482050 995508 482352 995527
rect 482722 995508 482976 995536
rect 482722 995443 482750 995508
rect 482710 995437 482762 995443
rect 482710 995379 482762 995385
rect 479828 994514 479884 994523
rect 479828 994449 479884 994458
rect 484162 993815 484190 995522
rect 485376 995508 485630 995536
rect 485602 995147 485630 995508
rect 485590 995141 485642 995147
rect 485590 995083 485642 995089
rect 485986 994671 486014 995522
rect 485972 994662 486028 994671
rect 485972 994597 486028 994606
rect 484150 993809 484202 993815
rect 484150 993751 484202 993757
rect 487810 993667 487838 995522
rect 487798 993661 487850 993667
rect 487798 993603 487850 993609
rect 489538 993593 489566 1002409
rect 505076 1002358 505132 1002367
rect 505076 1002293 505078 1002302
rect 505130 1002293 505132 1002302
rect 505078 1002261 505130 1002267
rect 513538 1001511 513566 1002409
rect 513526 1001505 513578 1001511
rect 513526 1001447 513578 1001453
rect 510932 1001026 510988 1001035
rect 510932 1000961 510934 1000970
rect 510986 1000961 510988 1000970
rect 510934 1000929 510986 1000935
rect 509300 1000878 509356 1000887
rect 509300 1000813 509302 1000822
rect 509354 1000813 509356 1000822
rect 509302 1000781 509354 1000787
rect 497590 999507 497642 999513
rect 497590 999449 497642 999455
rect 497602 999407 497630 999449
rect 497588 999398 497644 999407
rect 497588 999333 497644 999342
rect 506324 999398 506380 999407
rect 515458 999384 515486 1002483
rect 515734 1001505 515786 1001511
rect 515734 1001447 515786 1001453
rect 515458 999356 515582 999384
rect 506324 999333 506326 999342
rect 506378 999333 506380 999342
rect 506326 999301 506378 999307
rect 510262 996621 510314 996627
rect 507860 996586 507916 996595
rect 507860 996521 507862 996530
rect 507914 996521 507916 996530
rect 510260 996586 510262 996595
rect 510314 996586 510316 996595
rect 510260 996521 510316 996530
rect 507862 996489 507914 996495
rect 511894 996251 511946 996257
rect 511894 996193 511946 996199
rect 511124 996142 511180 996151
rect 511124 996077 511126 996086
rect 511178 996077 511180 996086
rect 511126 996045 511178 996051
rect 511906 996035 511934 996193
rect 513430 996177 513482 996183
rect 513428 996142 513430 996151
rect 513482 996142 513484 996151
rect 513428 996077 513484 996086
rect 511894 996029 511946 996035
rect 511892 995994 511894 996003
rect 513430 996029 513482 996035
rect 511946 995994 511948 996003
rect 511892 995929 511948 995938
rect 513428 995994 513430 996003
rect 513482 995994 513484 996003
rect 513428 995929 513484 995938
rect 506612 995402 506668 995411
rect 506612 995337 506668 995346
rect 506626 993741 506654 995337
rect 515554 994671 515582 999356
rect 515540 994662 515596 994671
rect 515540 994597 515596 994606
rect 515746 993815 515774 1001447
rect 516692 1001026 516748 1001035
rect 516692 1000961 516694 1000970
rect 516746 1000961 516748 1000970
rect 516694 1000929 516746 1000935
rect 516692 1000878 516748 1000887
rect 516692 1000813 516694 1000822
rect 516746 1000813 516748 1000822
rect 516694 1000781 516746 1000787
rect 516802 1000739 516830 1005221
rect 521206 1004909 521258 1004915
rect 521206 1004851 521258 1004857
rect 519478 1003873 519530 1003879
rect 519478 1003815 519530 1003821
rect 518614 1002393 518666 1002399
rect 518614 1002335 518666 1002341
rect 516788 1000730 516844 1000739
rect 516788 1000665 516844 1000674
rect 516692 999546 516748 999555
rect 516692 999481 516694 999490
rect 516746 999481 516748 999490
rect 516694 999449 516746 999455
rect 516692 999398 516748 999407
rect 516692 999333 516694 999342
rect 516746 999333 516748 999342
rect 516694 999301 516746 999307
rect 518420 995698 518476 995707
rect 518420 995633 518476 995642
rect 515734 993809 515786 993815
rect 515734 993751 515786 993757
rect 506614 993735 506666 993741
rect 506614 993677 506666 993683
rect 469460 993561 469462 993570
rect 469514 993561 469516 993570
rect 479158 993587 479210 993593
rect 469462 993529 469514 993535
rect 479158 993529 479210 993535
rect 489526 993587 489578 993593
rect 489526 993529 489578 993535
rect 518434 987821 518462 995633
rect 518516 995550 518572 995559
rect 518516 995485 518572 995494
rect 518422 987815 518474 987821
rect 518422 987757 518474 987763
rect 445078 986483 445130 986489
rect 445078 986425 445130 986431
rect 478966 986483 479018 986489
rect 478966 986425 479018 986431
rect 444886 985151 444938 985157
rect 444886 985093 444938 985099
rect 462742 985151 462794 985157
rect 462742 985093 462794 985099
rect 446422 985077 446474 985083
rect 446422 985019 446474 985025
rect 446434 981314 446462 985019
rect 462754 981314 462782 985093
rect 478978 981314 479006 986425
rect 518530 986415 518558 995485
rect 518626 995369 518654 1002335
rect 519490 995855 519518 1003815
rect 521014 1003725 521066 1003731
rect 521014 1003667 521066 1003673
rect 519476 995846 519532 995855
rect 519476 995781 519532 995790
rect 521026 995559 521054 1003667
rect 521218 998792 521246 1004851
rect 521410 999703 521438 1005221
rect 523990 1005205 524042 1005211
rect 553750 1005205 553802 1005211
rect 523990 1005147 524042 1005153
rect 547124 1005170 547180 1005179
rect 521494 1002319 521546 1002325
rect 521494 1002261 521546 1002267
rect 521396 999694 521452 999703
rect 521396 999629 521452 999638
rect 521506 999555 521534 1002261
rect 523604 1001026 523660 1001035
rect 523604 1000961 523660 1000970
rect 523508 1000730 523564 1000739
rect 523508 1000665 523564 1000674
rect 523412 999990 523468 999999
rect 523412 999925 523468 999934
rect 521492 999546 521548 999555
rect 521492 999481 521548 999490
rect 521218 998764 521342 998792
rect 521110 996621 521162 996627
rect 521110 996563 521162 996569
rect 521012 995550 521068 995559
rect 521012 995485 521068 995494
rect 521122 995443 521150 996563
rect 521206 996547 521258 996553
rect 521206 996489 521258 996495
rect 521218 995707 521246 996489
rect 521204 995698 521260 995707
rect 521204 995633 521260 995642
rect 521110 995437 521162 995443
rect 521110 995379 521162 995385
rect 518614 995363 518666 995369
rect 518614 995305 518666 995311
rect 521314 995221 521342 998764
rect 521396 995994 521452 996003
rect 521396 995929 521452 995938
rect 521302 995215 521354 995221
rect 521302 995157 521354 995163
rect 521410 986489 521438 995929
rect 523426 995411 523454 999925
rect 523522 995961 523550 1000665
rect 523510 995955 523562 995961
rect 523510 995897 523562 995903
rect 523618 995517 523646 1000961
rect 523700 1000878 523756 1000887
rect 523700 1000813 523756 1000822
rect 523714 995591 523742 1000813
rect 523892 999694 523948 999703
rect 523892 999629 523948 999638
rect 523796 999398 523852 999407
rect 523796 999333 523852 999342
rect 523810 995665 523838 999333
rect 523906 995887 523934 999629
rect 523894 995881 523946 995887
rect 523894 995823 523946 995829
rect 524002 995813 524030 1005147
rect 547124 1005105 547180 1005114
rect 553748 1005170 553750 1005179
rect 562486 1005205 562538 1005211
rect 553802 1005170 553804 1005179
rect 553748 1005105 553804 1005114
rect 562484 1005170 562486 1005179
rect 562538 1005170 562540 1005179
rect 562484 1005105 562540 1005114
rect 524084 999546 524140 999555
rect 524084 999481 524140 999490
rect 523990 995807 524042 995813
rect 523990 995749 524042 995755
rect 524098 995739 524126 999481
rect 540310 999433 540362 999439
rect 540310 999375 540362 999381
rect 532820 995846 532876 995855
rect 527842 995813 528192 995832
rect 528994 995813 529392 995832
rect 529858 995813 530064 995832
rect 527830 995807 528192 995813
rect 527882 995804 528192 995807
rect 528982 995807 529392 995813
rect 527830 995749 527882 995755
rect 529034 995804 529392 995807
rect 529846 995807 530064 995813
rect 528982 995749 529034 995755
rect 529898 995804 530064 995807
rect 532876 995804 533088 995832
rect 536784 995813 537182 995832
rect 540322 995813 540350 999375
rect 536784 995807 537194 995813
rect 536784 995804 537142 995807
rect 532820 995781 532876 995790
rect 529846 995749 529898 995755
rect 537142 995749 537194 995755
rect 540310 995807 540362 995813
rect 540310 995749 540362 995755
rect 524086 995733 524138 995739
rect 528406 995733 528458 995739
rect 524086 995675 524138 995681
rect 525346 995665 525744 995684
rect 532244 995698 532300 995707
rect 528458 995681 528768 995684
rect 528406 995675 528768 995681
rect 523798 995659 523850 995665
rect 523798 995601 523850 995607
rect 525334 995659 525744 995665
rect 525386 995656 525744 995659
rect 528418 995656 528768 995675
rect 532300 995656 532512 995684
rect 532244 995633 532300 995642
rect 525334 995601 525386 995607
rect 523702 995585 523754 995591
rect 523702 995527 523754 995533
rect 524758 995585 524810 995591
rect 534068 995550 534124 995559
rect 524810 995533 525072 995536
rect 524758 995527 525072 995533
rect 523606 995511 523658 995517
rect 524770 995508 525072 995527
rect 526114 995517 526368 995536
rect 530914 995522 531216 995536
rect 526102 995511 526368 995517
rect 523606 995453 523658 995459
rect 526154 995508 526368 995511
rect 526102 995453 526154 995459
rect 523412 995402 523468 995411
rect 530578 995369 530606 995522
rect 530914 995508 531230 995522
rect 530914 995411 530942 995508
rect 530900 995402 530956 995411
rect 523412 995337 523468 995346
rect 530566 995363 530618 995369
rect 530900 995337 530956 995346
rect 530566 995305 530618 995311
rect 530578 995240 530606 995305
rect 530578 995212 530654 995240
rect 530626 993667 530654 995212
rect 531202 994523 531230 995508
rect 533698 994671 533726 995522
rect 534124 995508 534384 995536
rect 535330 995508 535584 995536
rect 537154 995508 537408 995536
rect 538978 995508 539232 995536
rect 534068 995485 534124 995494
rect 533684 994662 533740 994671
rect 533684 994597 533740 994606
rect 531188 994514 531244 994523
rect 531188 994449 531244 994458
rect 535330 993815 535358 995508
rect 537154 995443 537182 995508
rect 537142 995437 537194 995443
rect 537142 995379 537194 995385
rect 535318 993809 535370 993815
rect 535318 993751 535370 993757
rect 538978 993741 539006 995508
rect 538966 993735 539018 993741
rect 538966 993677 539018 993683
rect 530614 993661 530666 993667
rect 530614 993603 530666 993609
rect 547138 992187 547166 1005105
rect 551734 1003873 551786 1003879
rect 551732 1003838 551734 1003847
rect 570646 1003873 570698 1003879
rect 551786 1003838 551788 1003847
rect 551732 1003773 551788 1003782
rect 556532 1003838 556588 1003847
rect 570646 1003815 570698 1003821
rect 556532 1003773 556534 1003782
rect 556586 1003773 556588 1003782
rect 556534 1003741 556586 1003747
rect 552598 1003725 552650 1003731
rect 552596 1003690 552598 1003699
rect 552650 1003690 552652 1003699
rect 552596 1003625 552652 1003634
rect 559126 1002541 559178 1002547
rect 559124 1002506 559126 1002515
rect 566134 1002541 566186 1002547
rect 559178 1002506 559180 1002515
rect 559124 1002441 559180 1002450
rect 559892 1002506 559948 1002515
rect 566134 1002483 566186 1002489
rect 559892 1002441 559894 1002450
rect 559946 1002441 559948 1002450
rect 564502 1002467 564554 1002473
rect 559894 1002409 559946 1002415
rect 564502 1002409 564554 1002415
rect 560566 1002393 560618 1002399
rect 560564 1002358 560566 1002367
rect 560618 1002358 560620 1002367
rect 560564 1002293 560620 1002302
rect 561524 1002358 561580 1002367
rect 561524 1002293 561526 1002302
rect 561578 1002293 561580 1002302
rect 561526 1002261 561578 1002267
rect 564514 1001067 564542 1002409
rect 564694 1002393 564746 1002399
rect 564790 1002393 564842 1002399
rect 564694 1002335 564746 1002341
rect 564788 1002358 564790 1002367
rect 564842 1002358 564844 1002367
rect 564502 1001061 564554 1001067
rect 564502 1001003 564554 1001009
rect 555190 997953 555242 997959
rect 555188 997918 555190 997927
rect 559894 997953 559946 997959
rect 555242 997918 555244 997927
rect 555188 997853 555244 997862
rect 557300 997918 557356 997927
rect 559894 997895 559946 997901
rect 557300 997853 557302 997862
rect 557354 997853 557356 997862
rect 557302 997821 557354 997827
rect 556150 997805 556202 997811
rect 556148 997770 556150 997779
rect 556202 997770 556204 997779
rect 556148 997705 556204 997714
rect 559906 997515 559934 997895
rect 564706 997737 564734 1002335
rect 564788 1002293 564844 1002302
rect 565366 1002319 565418 1002325
rect 565366 1002261 565418 1002267
rect 565378 999513 565406 1002261
rect 566146 1001659 566174 1002483
rect 568726 1002393 568778 1002399
rect 568726 1002335 568778 1002341
rect 566134 1001653 566186 1001659
rect 566134 1001595 566186 1001601
rect 567766 1001061 567818 1001067
rect 567766 1001003 567818 1001009
rect 565366 999507 565418 999513
rect 565366 999449 565418 999455
rect 567778 998625 567806 1001003
rect 567766 998619 567818 998625
rect 567766 998561 567818 998567
rect 564694 997731 564746 997737
rect 564694 997673 564746 997679
rect 559894 997509 559946 997515
rect 559894 997451 559946 997457
rect 563734 996177 563786 996183
rect 563734 996119 563786 996125
rect 562774 996103 562826 996109
rect 562774 996045 562826 996051
rect 562786 995707 562814 996045
rect 563746 995855 563774 996119
rect 564790 996029 564842 996035
rect 564788 995994 564790 996003
rect 564842 995994 564844 996003
rect 564788 995929 564844 995938
rect 563732 995846 563788 995855
rect 563732 995781 563734 995790
rect 563786 995781 563788 995790
rect 567478 995807 567530 995813
rect 563734 995749 563786 995755
rect 567478 995749 567530 995755
rect 562772 995698 562828 995707
rect 562772 995633 562774 995642
rect 562826 995633 562828 995642
rect 567382 995659 567434 995665
rect 562774 995601 562826 995607
rect 567382 995601 567434 995607
rect 557972 995402 558028 995411
rect 557972 995337 558028 995346
rect 557986 993741 558014 995337
rect 557974 993735 558026 993741
rect 557974 993677 558026 993683
rect 547126 992181 547178 992187
rect 547126 992123 547178 992129
rect 527542 987815 527594 987821
rect 527542 987757 527594 987763
rect 521398 986483 521450 986489
rect 521398 986425 521450 986431
rect 495094 986409 495146 986415
rect 495094 986351 495146 986357
rect 518518 986409 518570 986415
rect 518518 986351 518570 986357
rect 495106 981314 495134 986351
rect 511414 985003 511466 985009
rect 511414 984945 511466 984951
rect 511426 981314 511454 984945
rect 527554 981314 527582 987757
rect 543766 986483 543818 986489
rect 543766 986425 543818 986431
rect 543778 981314 543806 986425
rect 560086 986409 560138 986415
rect 560086 986351 560138 986357
rect 560098 981314 560126 986351
rect 567394 983677 567422 995601
rect 567382 983671 567434 983677
rect 567382 983613 567434 983619
rect 567490 983603 567518 995749
rect 567478 983597 567530 983603
rect 567478 983539 567530 983545
rect 568738 983529 568766 1002335
rect 570166 1001653 570218 1001659
rect 570166 1001595 570218 1001601
rect 570178 997756 570206 1001595
rect 570262 999433 570314 999439
rect 570262 999375 570314 999381
rect 570274 997959 570302 999375
rect 570262 997953 570314 997959
rect 570262 997895 570314 997901
rect 570178 997728 570398 997756
rect 570260 995698 570316 995707
rect 570260 995633 570316 995642
rect 570274 986563 570302 995633
rect 570370 994819 570398 997728
rect 570550 997509 570602 997515
rect 570550 997451 570602 997457
rect 570452 995550 570508 995559
rect 570452 995485 570508 995494
rect 570356 994810 570412 994819
rect 570356 994745 570412 994754
rect 570262 986557 570314 986563
rect 570262 986499 570314 986505
rect 570466 986415 570494 995485
rect 570562 993815 570590 997451
rect 570658 993889 570686 1003815
rect 571906 1001067 571934 1005221
rect 572866 1001511 572894 1005369
rect 572950 1005205 573002 1005211
rect 572950 1005147 573002 1005153
rect 572854 1001505 572906 1001511
rect 572854 1001447 572906 1001453
rect 571894 1001061 571946 1001067
rect 571894 1001003 571946 1001009
rect 571030 999359 571082 999365
rect 571030 999301 571082 999307
rect 570838 998619 570890 998625
rect 570838 998561 570890 998567
rect 570850 994967 570878 998561
rect 570836 994958 570892 994967
rect 570836 994893 570892 994902
rect 571042 994671 571070 999301
rect 572962 997515 572990 1005147
rect 574486 1003799 574538 1003805
rect 574486 1003741 574538 1003747
rect 573046 1003725 573098 1003731
rect 573046 1003667 573098 1003673
rect 573058 1002251 573086 1003667
rect 573046 1002245 573098 1002251
rect 573046 1002187 573098 1002193
rect 573334 1002245 573386 1002251
rect 573334 1002187 573386 1002193
rect 573238 1001061 573290 1001067
rect 573238 1001003 573290 1001009
rect 573250 997589 573278 1001003
rect 573346 997663 573374 1002187
rect 574102 1001505 574154 1001511
rect 574102 1001447 574154 1001453
rect 573334 997657 573386 997663
rect 573334 997599 573386 997605
rect 573238 997583 573290 997589
rect 573238 997525 573290 997531
rect 572950 997509 573002 997515
rect 572950 997451 573002 997457
rect 573140 995846 573196 995855
rect 573140 995781 573196 995790
rect 571028 994662 571084 994671
rect 571028 994597 571084 994606
rect 570646 993883 570698 993889
rect 570646 993825 570698 993831
rect 570550 993809 570602 993815
rect 570550 993751 570602 993757
rect 573154 986489 573182 995781
rect 574114 994037 574142 1001447
rect 574498 997441 574526 1003741
rect 613462 999877 613514 999883
rect 613462 999819 613514 999825
rect 625558 999877 625610 999883
rect 625558 999819 625610 999825
rect 610582 999803 610634 999809
rect 610582 999745 610634 999751
rect 601846 999729 601898 999735
rect 601846 999671 601898 999677
rect 596182 999655 596234 999661
rect 596182 999597 596234 999603
rect 590710 999581 590762 999587
rect 590710 999523 590762 999529
rect 590614 999507 590666 999513
rect 590614 999449 590666 999455
rect 590518 999433 590570 999439
rect 590518 999375 590570 999381
rect 590530 997811 590558 999375
rect 590518 997805 590570 997811
rect 590518 997747 590570 997753
rect 590626 997737 590654 999449
rect 590614 997731 590666 997737
rect 590614 997673 590666 997679
rect 590722 997663 590750 999523
rect 596194 997885 596222 999597
rect 596182 997879 596234 997885
rect 596182 997821 596234 997827
rect 590710 997657 590762 997663
rect 590710 997599 590762 997605
rect 601858 997515 601886 999671
rect 610594 997589 610622 999745
rect 610678 997953 610730 997959
rect 610678 997895 610730 997901
rect 610582 997583 610634 997589
rect 610582 997525 610634 997531
rect 601846 997509 601898 997515
rect 601846 997451 601898 997457
rect 574486 997435 574538 997441
rect 574486 997377 574538 997383
rect 610690 995887 610718 997895
rect 613474 997441 613502 999819
rect 625462 999803 625514 999809
rect 625462 999745 625514 999751
rect 625366 999581 625418 999587
rect 625366 999523 625418 999529
rect 613462 997435 613514 997441
rect 613462 997377 613514 997383
rect 625378 996035 625406 999523
rect 625366 996029 625418 996035
rect 625366 995971 625418 995977
rect 625474 995961 625502 999745
rect 625462 995955 625514 995961
rect 625462 995897 625514 995903
rect 610678 995881 610730 995887
rect 610678 995823 610730 995829
rect 616342 995881 616394 995887
rect 616342 995823 616394 995829
rect 574102 994031 574154 994037
rect 574102 993973 574154 993979
rect 576020 993922 576076 993931
rect 576020 993857 576076 993866
rect 573142 986483 573194 986489
rect 573142 986425 573194 986431
rect 570454 986409 570506 986415
rect 570454 986351 570506 986357
rect 568726 983523 568778 983529
rect 568726 983465 568778 983471
rect 576034 981328 576062 993857
rect 616354 989301 616382 995823
rect 625570 995591 625598 999819
rect 625846 999729 625898 999735
rect 625898 999677 625982 999680
rect 625846 999671 625982 999677
rect 625750 999655 625802 999661
rect 625858 999652 625982 999671
rect 625750 999597 625802 999603
rect 625654 999433 625706 999439
rect 625654 999375 625706 999381
rect 625666 995887 625694 999375
rect 625654 995881 625706 995887
rect 625654 995823 625706 995829
rect 625762 995739 625790 999597
rect 625846 999507 625898 999513
rect 625846 999449 625898 999455
rect 625858 995813 625886 999449
rect 625846 995807 625898 995813
rect 625846 995749 625898 995755
rect 625750 995733 625802 995739
rect 625750 995675 625802 995681
rect 625954 995665 625982 999652
rect 626530 995813 626880 995832
rect 630946 995813 631200 995832
rect 631522 995813 631824 995832
rect 634594 995813 634896 995832
rect 626518 995807 626880 995813
rect 626570 995804 626880 995807
rect 630934 995807 631200 995813
rect 626518 995749 626570 995755
rect 630986 995804 631200 995807
rect 631510 995807 631824 995813
rect 630934 995749 630986 995755
rect 631562 995804 631824 995807
rect 634582 995807 634896 995813
rect 631510 995749 631562 995755
rect 634634 995804 634896 995807
rect 634582 995749 634634 995755
rect 627094 995733 627146 995739
rect 627146 995681 627504 995684
rect 627094 995675 627504 995681
rect 625942 995659 625994 995665
rect 627106 995656 627504 995675
rect 627874 995665 628176 995684
rect 627862 995659 628176 995665
rect 625942 995601 625994 995607
rect 627914 995656 628176 995659
rect 627862 995601 627914 995607
rect 625558 995585 625610 995591
rect 625558 995527 625610 995533
rect 630166 995585 630218 995591
rect 630218 995533 630576 995536
rect 630166 995527 630576 995533
rect 629986 994967 630014 995522
rect 630178 995508 630576 995527
rect 629972 994958 630028 994967
rect 629972 994893 630028 994902
rect 630740 994514 630796 994523
rect 630740 994449 630796 994458
rect 616342 989295 616394 989301
rect 616342 989237 616394 989243
rect 592438 986557 592490 986563
rect 592438 986499 592490 986505
rect 576034 981300 576240 981328
rect 592450 981314 592478 986499
rect 608758 986483 608810 986489
rect 608758 986425 608810 986431
rect 608770 981314 608798 986425
rect 624886 986409 624938 986415
rect 624886 986351 624938 986357
rect 624898 981314 624926 986351
rect 630754 980643 630782 994449
rect 632386 994407 632414 995522
rect 632770 995508 633024 995536
rect 632770 994523 632798 995508
rect 633718 995215 633770 995221
rect 633718 995157 633770 995163
rect 632756 994514 632812 994523
rect 632756 994449 632812 994458
rect 630838 994401 630890 994407
rect 630838 994343 630890 994349
rect 632374 994401 632426 994407
rect 632374 994343 632426 994349
rect 630850 993667 630878 994343
rect 633620 993774 633676 993783
rect 633620 993709 633676 993718
rect 630838 993661 630890 993667
rect 630838 993603 630890 993609
rect 630850 980717 630878 993603
rect 633634 985009 633662 993709
rect 633730 990707 633758 995157
rect 634306 994819 634334 995522
rect 635266 995508 635520 995536
rect 634292 994810 634348 994819
rect 634292 994745 634348 994754
rect 635266 994037 635294 995508
rect 635254 994031 635306 994037
rect 635254 993973 635306 993979
rect 636130 993889 636158 995522
rect 636118 993883 636170 993889
rect 636118 993825 636170 993831
rect 637378 993815 637406 995522
rect 638544 995508 638942 995536
rect 638516 994366 638572 994375
rect 638516 994301 638572 994310
rect 637366 993809 637418 993815
rect 637366 993751 637418 993757
rect 633718 990701 633770 990707
rect 633718 990643 633770 990649
rect 638530 989375 638558 994301
rect 638914 993667 638942 995508
rect 639202 994671 639230 995522
rect 639188 994662 639244 994671
rect 639188 994597 639244 994606
rect 640724 994218 640780 994227
rect 640724 994153 640780 994162
rect 638902 993661 638954 993667
rect 638902 993603 638954 993609
rect 640438 990701 640490 990707
rect 640438 990643 640490 990649
rect 638518 989369 638570 989375
rect 638518 989311 638570 989317
rect 640450 986341 640478 990643
rect 640738 989819 640766 994153
rect 641026 993741 641054 995522
rect 643990 995141 644042 995147
rect 643990 995083 644042 995089
rect 642454 995067 642506 995073
rect 642454 995009 642506 995015
rect 641014 993735 641066 993741
rect 641014 993677 641066 993683
rect 640726 989813 640778 989819
rect 640726 989755 640778 989761
rect 642466 987821 642494 995009
rect 643606 993661 643658 993667
rect 643606 993603 643658 993609
rect 643222 989295 643274 989301
rect 643222 989237 643274 989243
rect 642454 987815 642506 987821
rect 642454 987757 642506 987763
rect 640438 986335 640490 986341
rect 640438 986277 640490 986283
rect 633622 985003 633674 985009
rect 633622 984945 633674 984951
rect 641110 985003 641162 985009
rect 641110 984945 641162 984951
rect 641122 981314 641150 984945
rect 643234 984935 643262 989237
rect 643222 984929 643274 984935
rect 643222 984871 643274 984877
rect 643618 980865 643646 993603
rect 644002 990707 644030 995083
rect 650036 994070 650092 994079
rect 650036 994005 650092 994014
rect 643990 990701 644042 990707
rect 643990 990643 644042 990649
rect 649846 990701 649898 990707
rect 649846 990643 649898 990649
rect 649558 989813 649610 989819
rect 649558 989755 649610 989761
rect 647350 987815 647402 987821
rect 647350 987757 647402 987763
rect 646102 986335 646154 986341
rect 646102 986277 646154 986283
rect 643606 980859 643658 980865
rect 643606 980801 643658 980807
rect 630838 980711 630890 980717
rect 630838 980653 630890 980659
rect 410326 980637 410378 980643
rect 410326 980579 410378 980585
rect 630742 980637 630794 980643
rect 630742 980579 630794 980585
rect 646114 980569 646142 986277
rect 647362 980791 647390 987757
rect 647350 980785 647402 980791
rect 647350 980727 647402 980733
rect 649462 980785 649514 980791
rect 649462 980727 649514 980733
rect 646102 980563 646154 980569
rect 646102 980505 646154 980511
rect 649366 980563 649418 980569
rect 649366 980505 649418 980511
rect 630658 275636 630864 275664
rect 65890 259111 65918 275502
rect 66838 275121 66890 275127
rect 66838 275063 66890 275069
rect 66164 273310 66220 273319
rect 66164 273245 66166 273254
rect 66218 273245 66220 273254
rect 66166 273213 66218 273219
rect 66850 266691 66878 275063
rect 66946 269323 66974 275502
rect 67222 275195 67274 275201
rect 67222 275137 67274 275143
rect 67234 270687 67262 275137
rect 67606 270977 67658 270983
rect 67606 270919 67658 270925
rect 67222 270681 67274 270687
rect 67222 270623 67274 270629
rect 66932 269314 66988 269323
rect 66932 269249 66988 269258
rect 66838 266685 66890 266691
rect 66838 266627 66890 266633
rect 65876 259102 65932 259111
rect 65876 259037 65932 259046
rect 65206 254919 65258 254925
rect 65206 254861 65258 254867
rect 65108 254810 65164 254819
rect 65108 254745 65164 254754
rect 67618 252779 67646 270919
rect 68194 269873 68222 275502
rect 68182 269867 68234 269873
rect 68182 269809 68234 269815
rect 69346 269767 69374 275502
rect 69332 269758 69388 269767
rect 69332 269693 69388 269702
rect 70594 258963 70622 275502
rect 71746 269471 71774 275502
rect 72598 273493 72650 273499
rect 72598 273435 72650 273441
rect 72118 270681 72170 270687
rect 72118 270623 72170 270629
rect 71732 269462 71788 269471
rect 71732 269397 71788 269406
rect 72130 266839 72158 270623
rect 72610 270613 72638 273435
rect 72598 270607 72650 270613
rect 72598 270549 72650 270555
rect 72118 266833 72170 266839
rect 72118 266775 72170 266781
rect 72994 263551 73022 275502
rect 72980 263542 73036 263551
rect 72980 263477 73036 263486
rect 70580 258954 70636 258963
rect 70580 258889 70636 258898
rect 74146 258815 74174 275502
rect 75298 270021 75326 275502
rect 75286 270015 75338 270021
rect 75286 269957 75338 269963
rect 74132 258806 74188 258815
rect 74132 258741 74188 258750
rect 76546 258667 76574 275502
rect 77698 269915 77726 275502
rect 77684 269906 77740 269915
rect 77684 269841 77740 269850
rect 76532 258658 76588 258667
rect 76532 258593 76588 258602
rect 78946 258519 78974 275502
rect 80098 270095 80126 275502
rect 80564 273310 80620 273319
rect 80564 273245 80566 273254
rect 80618 273245 80620 273254
rect 80566 273213 80618 273219
rect 80662 270607 80714 270613
rect 80662 270549 80714 270555
rect 80086 270089 80138 270095
rect 80086 270031 80138 270037
rect 80566 266685 80618 266691
rect 80566 266627 80618 266633
rect 80578 259088 80606 266627
rect 80674 261437 80702 270549
rect 81346 269619 81374 275502
rect 81332 269610 81388 269619
rect 81332 269545 81388 269554
rect 82498 266395 82526 275502
rect 83650 270063 83678 275502
rect 84802 270169 84830 275502
rect 84790 270163 84842 270169
rect 84790 270105 84842 270111
rect 83636 270054 83692 270063
rect 83636 269989 83692 269998
rect 83638 266833 83690 266839
rect 83638 266775 83690 266781
rect 82486 266389 82538 266395
rect 82486 266331 82538 266337
rect 80662 261431 80714 261437
rect 80662 261373 80714 261379
rect 83542 261431 83594 261437
rect 83542 261373 83594 261379
rect 80578 259060 80894 259088
rect 78932 258510 78988 258519
rect 78932 258445 78988 258454
rect 80662 255733 80714 255739
rect 80660 255698 80662 255707
rect 80714 255698 80716 255707
rect 80660 255633 80716 255642
rect 80866 252853 80894 259060
rect 83554 254999 83582 261373
rect 83650 258107 83678 266775
rect 86050 258371 86078 275502
rect 86228 273310 86284 273319
rect 86420 273310 86476 273319
rect 86284 273268 86420 273296
rect 86228 273245 86284 273254
rect 86420 273245 86476 273254
rect 86036 258362 86092 258371
rect 86036 258297 86092 258306
rect 83638 258101 83690 258107
rect 87202 258075 87230 275502
rect 83638 258043 83690 258049
rect 87188 258066 87244 258075
rect 87188 258001 87244 258010
rect 88450 257779 88478 275502
rect 89602 270243 89630 275502
rect 89590 270237 89642 270243
rect 90754 270211 90782 275502
rect 89590 270179 89642 270185
rect 90740 270202 90796 270211
rect 90740 270137 90796 270146
rect 92002 258223 92030 275502
rect 93154 270359 93182 275502
rect 93140 270350 93196 270359
rect 94402 270317 94430 275502
rect 95554 270507 95582 275502
rect 95540 270498 95596 270507
rect 95540 270433 95596 270442
rect 93140 270285 93196 270294
rect 94390 270311 94442 270317
rect 94390 270253 94442 270259
rect 91988 258214 92044 258223
rect 91988 258149 92044 258158
rect 96310 258101 96362 258107
rect 96310 258043 96362 258049
rect 88436 257770 88492 257779
rect 88436 257705 88492 257714
rect 86708 255698 86764 255707
rect 86708 255633 86710 255642
rect 86762 255633 86764 255642
rect 86710 255601 86762 255607
rect 83542 254993 83594 254999
rect 83542 254935 83594 254941
rect 96322 252927 96350 258043
rect 96802 257927 96830 275502
rect 97954 270391 97982 275502
rect 97942 270385 97994 270391
rect 97942 270327 97994 270333
rect 99202 257959 99230 275502
rect 100258 270655 100286 275502
rect 100916 273458 100972 273467
rect 100916 273393 100918 273402
rect 100970 273393 100972 273402
rect 100918 273361 100970 273367
rect 100244 270646 100300 270655
rect 100244 270581 100300 270590
rect 101506 270465 101534 275502
rect 101494 270459 101546 270465
rect 101494 270401 101546 270407
rect 102658 269281 102686 275502
rect 102646 269275 102698 269281
rect 102646 269217 102698 269223
rect 99190 257953 99242 257959
rect 96788 257918 96844 257927
rect 99190 257895 99242 257901
rect 96788 257853 96844 257862
rect 103906 257811 103934 275502
rect 105058 270539 105086 275502
rect 105046 270533 105098 270539
rect 105046 270475 105098 270481
rect 106210 258033 106238 275502
rect 107458 269175 107486 275502
rect 108610 270613 108638 275502
rect 108598 270607 108650 270613
rect 108598 270549 108650 270555
rect 109858 269355 109886 275502
rect 109846 269349 109898 269355
rect 109846 269291 109898 269297
rect 107444 269166 107500 269175
rect 107444 269101 107500 269110
rect 106198 258027 106250 258033
rect 106198 257969 106250 257975
rect 111010 257885 111038 275502
rect 112258 270687 112286 275502
rect 112246 270681 112298 270687
rect 112246 270623 112298 270629
rect 113410 263699 113438 275502
rect 114658 269429 114686 275502
rect 114646 269423 114698 269429
rect 114646 269365 114698 269371
rect 115810 269207 115838 275502
rect 115798 269201 115850 269207
rect 115798 269143 115850 269149
rect 116962 263847 116990 275502
rect 116948 263838 117004 263847
rect 116948 263773 117004 263782
rect 113396 263690 113452 263699
rect 113396 263625 113452 263634
rect 118114 258107 118142 275502
rect 119362 269133 119390 275502
rect 119350 269127 119402 269133
rect 119350 269069 119402 269075
rect 120514 263995 120542 275502
rect 120788 273458 120844 273467
rect 120788 273393 120790 273402
rect 120842 273393 120844 273402
rect 120790 273361 120842 273367
rect 121666 269577 121694 275502
rect 121654 269571 121706 269577
rect 121654 269513 121706 269519
rect 122914 268763 122942 275502
rect 122902 268757 122954 268763
rect 122902 268699 122954 268705
rect 120500 263986 120556 263995
rect 120500 263921 120556 263930
rect 124066 263065 124094 275502
rect 125314 266617 125342 275502
rect 126466 268985 126494 275502
rect 127714 269651 127742 275502
rect 127702 269645 127754 269651
rect 127702 269587 127754 269593
rect 128866 269503 128894 275502
rect 130114 270613 130142 275502
rect 130006 270607 130058 270613
rect 130006 270549 130058 270555
rect 130102 270607 130154 270613
rect 130102 270549 130154 270555
rect 128854 269497 128906 269503
rect 128854 269439 128906 269445
rect 126454 268979 126506 268985
rect 126454 268921 126506 268927
rect 130018 268911 130046 270549
rect 130006 268905 130058 268911
rect 130006 268847 130058 268853
rect 125302 266611 125354 266617
rect 125302 266553 125354 266559
rect 124054 263059 124106 263065
rect 124054 263001 124106 263007
rect 131266 260697 131294 275502
rect 132514 269799 132542 275502
rect 132982 270681 133034 270687
rect 132982 270623 133034 270629
rect 132994 270391 133022 270623
rect 132886 270385 132938 270391
rect 132886 270327 132938 270333
rect 132982 270385 133034 270391
rect 132982 270327 133034 270333
rect 132502 269793 132554 269799
rect 132502 269735 132554 269741
rect 132898 268837 132926 270327
rect 133570 270021 133598 275502
rect 133558 270015 133610 270021
rect 133558 269957 133610 269963
rect 133270 269867 133322 269873
rect 133270 269809 133322 269815
rect 133282 269059 133310 269809
rect 134818 269725 134846 275502
rect 134806 269719 134858 269725
rect 134806 269661 134858 269667
rect 133270 269053 133322 269059
rect 133270 268995 133322 269001
rect 132886 268831 132938 268837
rect 132886 268773 132938 268779
rect 135970 266691 135998 275502
rect 137122 270687 137150 275502
rect 137110 270681 137162 270687
rect 137110 270623 137162 270629
rect 135958 266685 136010 266691
rect 135958 266627 136010 266633
rect 138370 260771 138398 275502
rect 139318 270533 139370 270539
rect 139318 270475 139370 270481
rect 139126 270385 139178 270391
rect 139126 270327 139178 270333
rect 139138 269448 139166 270327
rect 139330 269596 139358 270475
rect 139414 270089 139466 270095
rect 139414 270031 139466 270037
rect 139426 269744 139454 270031
rect 139522 269947 139550 275502
rect 140784 275488 141086 275516
rect 140470 270681 140522 270687
rect 140470 270623 140522 270629
rect 139894 270607 139946 270613
rect 139894 270549 139946 270555
rect 139702 270459 139754 270465
rect 139702 270401 139754 270407
rect 139510 269941 139562 269947
rect 139510 269883 139562 269889
rect 139426 269716 139550 269744
rect 139330 269568 139454 269596
rect 139138 269420 139358 269448
rect 139222 267795 139274 267801
rect 139222 267737 139274 267743
rect 138358 260765 138410 260771
rect 138358 260707 138410 260713
rect 131254 260691 131306 260697
rect 131254 260633 131306 260639
rect 118102 258101 118154 258107
rect 118102 258043 118154 258049
rect 110998 257879 111050 257885
rect 110998 257821 111050 257827
rect 103894 257805 103946 257811
rect 103894 257747 103946 257753
rect 138164 255846 138220 255855
rect 138164 255781 138220 255790
rect 138178 255739 138206 255781
rect 106678 255733 106730 255739
rect 106498 255681 106678 255684
rect 118102 255733 118154 255739
rect 106498 255675 106730 255681
rect 118100 255698 118102 255707
rect 138166 255733 138218 255739
rect 118154 255698 118156 255707
rect 106498 255665 106718 255675
rect 106486 255659 106718 255665
rect 106538 255656 106718 255659
rect 138166 255675 138218 255681
rect 118100 255633 118156 255642
rect 106486 255601 106538 255607
rect 112150 254993 112202 254999
rect 112150 254935 112202 254941
rect 112162 253001 112190 254935
rect 112150 252995 112202 253001
rect 112150 252937 112202 252943
rect 96310 252921 96362 252927
rect 96310 252863 96362 252869
rect 80854 252847 80906 252853
rect 80854 252789 80906 252795
rect 67606 252773 67658 252779
rect 67606 252715 67658 252721
rect 139234 250781 139262 267737
rect 139222 250775 139274 250781
rect 139222 250717 139274 250723
rect 139330 250263 139358 269420
rect 139318 250257 139370 250263
rect 139318 250199 139370 250205
rect 50422 237751 50474 237757
rect 50422 237693 50474 237699
rect 139426 233484 139454 269568
rect 139522 239996 139550 269716
rect 139606 268905 139658 268911
rect 139606 268847 139658 268853
rect 139618 240292 139646 268847
rect 139714 267801 139742 270401
rect 139798 270237 139850 270243
rect 139798 270179 139850 270185
rect 139702 267795 139754 267801
rect 139702 267737 139754 267743
rect 139810 250189 139838 270179
rect 139798 250183 139850 250189
rect 139798 250125 139850 250131
rect 139906 250115 139934 270549
rect 140182 270311 140234 270317
rect 140182 270253 140234 270259
rect 140086 269867 140138 269873
rect 140086 269809 140138 269815
rect 139990 268757 140042 268763
rect 139990 268699 140042 268705
rect 139894 250109 139946 250115
rect 139894 250051 139946 250057
rect 140002 243677 140030 268699
rect 139990 243671 140042 243677
rect 139990 243613 140042 243619
rect 139618 240264 140030 240292
rect 139522 239968 139838 239996
rect 139426 233456 139646 233484
rect 139618 232744 139646 233456
rect 139426 232716 139646 232744
rect 139810 232744 139838 239968
rect 139810 232716 139934 232744
rect 139426 229340 139454 232716
rect 139906 229451 139934 232716
rect 140002 230265 140030 240264
rect 140098 235759 140126 269809
rect 140194 253149 140222 270253
rect 140374 270163 140426 270169
rect 140374 270105 140426 270111
rect 140278 270015 140330 270021
rect 140278 269957 140330 269963
rect 140182 253143 140234 253149
rect 140182 253085 140234 253091
rect 140182 250775 140234 250781
rect 140182 250717 140234 250723
rect 140194 240495 140222 250717
rect 140182 240489 140234 240495
rect 140182 240431 140234 240437
rect 140182 236197 140234 236203
rect 140182 236139 140234 236145
rect 140086 235753 140138 235759
rect 140086 235695 140138 235701
rect 140194 235167 140222 236139
rect 140182 235161 140234 235167
rect 140182 235103 140234 235109
rect 140290 230431 140318 269957
rect 140386 239237 140414 270105
rect 140374 239231 140426 239237
rect 140374 239173 140426 239179
rect 140482 239108 140510 270623
rect 140566 269201 140618 269207
rect 140566 269143 140618 269149
rect 140386 239080 140510 239108
rect 140278 230425 140330 230431
rect 140278 230367 140330 230373
rect 140002 230237 140318 230265
rect 139990 229463 140042 229469
rect 139906 229423 139990 229451
rect 139990 229405 140042 229411
rect 139426 229312 139934 229340
rect 139906 229229 139934 229312
rect 139990 229241 140042 229247
rect 139906 229201 139990 229229
rect 139990 229183 140042 229189
rect 140290 227619 140318 230237
rect 140386 229543 140414 239080
rect 140578 238960 140606 269143
rect 140758 269127 140810 269133
rect 140758 269069 140810 269075
rect 140662 268979 140714 268985
rect 140662 268921 140714 268927
rect 140482 238932 140606 238960
rect 140482 229691 140510 238932
rect 140566 238787 140618 238793
rect 140566 238729 140618 238735
rect 140470 229685 140522 229691
rect 140470 229627 140522 229633
rect 140374 229537 140426 229543
rect 140374 229479 140426 229485
rect 140578 229469 140606 238729
rect 140674 229839 140702 268921
rect 140770 229913 140798 269069
rect 140854 269053 140906 269059
rect 140854 268995 140906 269001
rect 140866 237609 140894 268995
rect 140950 268831 141002 268837
rect 140950 268773 141002 268779
rect 140962 238793 140990 268773
rect 140950 238787 141002 238793
rect 140950 238729 141002 238735
rect 140854 237603 140906 237609
rect 140854 237545 140906 237551
rect 141058 237480 141086 275488
rect 141922 269873 141950 275502
rect 141910 269867 141962 269873
rect 141910 269809 141962 269815
rect 141142 263059 141194 263065
rect 141142 263001 141194 263007
rect 141154 262917 141182 263001
rect 141142 262911 141194 262917
rect 141142 262853 141194 262859
rect 143170 258181 143198 275502
rect 144322 268245 144350 275502
rect 144310 268239 144362 268245
rect 144310 268181 144362 268187
rect 145570 260105 145598 275502
rect 146722 270021 146750 275502
rect 146710 270015 146762 270021
rect 146710 269957 146762 269963
rect 147970 268689 147998 275502
rect 147958 268683 148010 268689
rect 147958 268625 148010 268631
rect 146518 268239 146570 268245
rect 146518 268181 146570 268187
rect 145558 260099 145610 260105
rect 145558 260041 145610 260047
rect 143158 258175 143210 258181
rect 143158 258117 143210 258123
rect 141142 255881 141194 255887
rect 141142 255823 141194 255829
rect 141154 255739 141182 255823
rect 141142 255733 141194 255739
rect 141142 255675 141194 255681
rect 141526 253143 141578 253149
rect 141526 253085 141578 253091
rect 141142 252921 141194 252927
rect 141142 252863 141194 252869
rect 141154 250337 141182 252863
rect 141142 250331 141194 250337
rect 141142 250273 141194 250279
rect 141334 250183 141386 250189
rect 141334 250125 141386 250131
rect 141238 250109 141290 250115
rect 141238 250051 141290 250057
rect 141142 239231 141194 239237
rect 141142 239173 141194 239179
rect 140866 237452 141086 237480
rect 140758 229907 140810 229913
rect 140758 229849 140810 229855
rect 140662 229833 140714 229839
rect 140662 229775 140714 229781
rect 140566 229463 140618 229469
rect 140566 229405 140618 229411
rect 139990 227613 140042 227619
rect 139990 227555 140042 227561
rect 140278 227613 140330 227619
rect 140278 227555 140330 227561
rect 140002 213115 140030 227555
rect 140866 218739 140894 237452
rect 140950 237381 141002 237387
rect 140950 237323 141002 237329
rect 140962 229765 140990 237323
rect 141154 236296 141182 239173
rect 141058 236268 141182 236296
rect 141058 230524 141086 236268
rect 141250 236203 141278 250051
rect 141238 236197 141290 236203
rect 141238 236139 141290 236145
rect 141346 236111 141374 250125
rect 141430 240489 141482 240495
rect 141430 240431 141482 240437
rect 141250 236083 141374 236111
rect 141250 236037 141278 236083
rect 141442 236037 141470 240431
rect 141154 236009 141278 236037
rect 141346 236009 141470 236037
rect 141154 232651 141182 236009
rect 141142 232645 141194 232651
rect 141142 232587 141194 232593
rect 141058 230496 141278 230524
rect 141046 230425 141098 230431
rect 141046 230367 141098 230373
rect 140950 229759 141002 229765
rect 140950 229701 141002 229707
rect 141058 229636 141086 230367
rect 141058 229608 141182 229636
rect 141154 229543 141182 229608
rect 141142 229537 141194 229543
rect 141142 229479 141194 229485
rect 141250 229321 141278 230496
rect 141238 229315 141290 229321
rect 141238 229257 141290 229263
rect 140854 218733 140906 218739
rect 140854 218675 140906 218681
rect 141346 216001 141374 236009
rect 141538 235852 141566 253085
rect 142486 252995 142538 253001
rect 142486 252937 142538 252943
rect 142198 243671 142250 243677
rect 142198 243613 142250 243619
rect 141442 235824 141566 235852
rect 141442 229247 141470 235824
rect 141526 235753 141578 235759
rect 141526 235695 141578 235701
rect 141430 229241 141482 229247
rect 141430 229183 141482 229189
rect 141538 221773 141566 235695
rect 141910 235161 141962 235167
rect 141910 235103 141962 235109
rect 141718 232645 141770 232651
rect 141718 232587 141770 232593
rect 141526 221767 141578 221773
rect 141526 221709 141578 221715
rect 141334 215995 141386 216001
rect 141334 215937 141386 215943
rect 141730 215927 141758 232587
rect 141922 218887 141950 235103
rect 141910 218881 141962 218887
rect 141910 218823 141962 218829
rect 142210 218813 142238 243613
rect 142498 233317 142526 252937
rect 145366 250627 145418 250633
rect 145366 250569 145418 250575
rect 145378 250411 145406 250569
rect 145366 250405 145418 250411
rect 145366 250347 145418 250353
rect 144406 250331 144458 250337
rect 144406 250273 144458 250279
rect 144310 250257 144362 250263
rect 144310 250199 144362 250205
rect 144020 248150 144076 248159
rect 144020 248085 144076 248094
rect 144034 247821 144062 248085
rect 144022 247815 144074 247821
rect 144022 247757 144074 247763
rect 144116 246374 144172 246383
rect 144116 246309 144172 246318
rect 144020 245338 144076 245347
rect 144020 245273 144076 245282
rect 144034 244861 144062 245273
rect 144130 244935 144158 246309
rect 144118 244929 144170 244935
rect 144118 244871 144170 244877
rect 144022 244855 144074 244861
rect 144022 244797 144074 244803
rect 144020 242822 144076 242831
rect 144020 242757 144076 242766
rect 144034 242049 144062 242757
rect 144022 242043 144074 242049
rect 144022 241985 144074 241991
rect 144020 239122 144076 239131
rect 144020 239057 144022 239066
rect 144074 239057 144076 239066
rect 144022 239025 144074 239031
rect 144020 237938 144076 237947
rect 144020 237873 144076 237882
rect 144034 236573 144062 237873
rect 144022 236567 144074 236573
rect 144022 236509 144074 236515
rect 144116 234386 144172 234395
rect 144116 234321 144172 234330
rect 144020 233498 144076 233507
rect 144020 233433 144076 233442
rect 144034 233391 144062 233433
rect 144022 233385 144074 233391
rect 144022 233327 144074 233333
rect 144130 233317 144158 234321
rect 142486 233311 142538 233317
rect 142486 233253 142538 233259
rect 144118 233311 144170 233317
rect 144118 233253 144170 233259
rect 144020 231278 144076 231287
rect 144020 231213 144076 231222
rect 144034 230505 144062 231213
rect 144022 230499 144074 230505
rect 144022 230441 144074 230447
rect 144116 229502 144172 229511
rect 144116 229437 144172 229446
rect 144020 228910 144076 228919
rect 144020 228845 144076 228854
rect 144034 227619 144062 228845
rect 144130 227693 144158 229437
rect 144322 229099 144350 250199
rect 144418 244491 144446 250273
rect 145460 249334 145516 249343
rect 145460 249269 145516 249278
rect 145474 247747 145502 249269
rect 145462 247741 145514 247747
rect 145462 247683 145514 247689
rect 144406 244485 144458 244491
rect 144406 244427 144458 244433
rect 145748 242082 145804 242091
rect 145748 242017 145804 242026
rect 145762 241975 145790 242017
rect 145750 241969 145802 241975
rect 145750 241911 145802 241917
rect 145364 236162 145420 236171
rect 145364 236097 145420 236106
rect 144310 229093 144362 229099
rect 144310 229035 144362 229041
rect 144118 227687 144170 227693
rect 144118 227629 144170 227635
rect 144022 227613 144074 227619
rect 144022 227555 144074 227561
rect 144020 225062 144076 225071
rect 144020 224997 144076 225006
rect 144034 224733 144062 224997
rect 144022 224727 144074 224733
rect 144022 224669 144074 224675
rect 144020 224026 144076 224035
rect 144020 223961 144076 223970
rect 144034 221847 144062 223961
rect 144022 221841 144074 221847
rect 144022 221783 144074 221789
rect 144116 221362 144172 221371
rect 144116 221297 144172 221306
rect 144020 220030 144076 220039
rect 144020 219965 144076 219974
rect 144034 218961 144062 219965
rect 144130 219035 144158 221297
rect 144118 219029 144170 219035
rect 144118 218971 144170 218977
rect 144022 218955 144074 218961
rect 144022 218897 144074 218903
rect 142198 218807 142250 218813
rect 142198 218749 142250 218755
rect 144020 218106 144076 218115
rect 144020 218041 144022 218050
rect 144074 218041 144076 218050
rect 144022 218009 144074 218015
rect 141718 215921 141770 215927
rect 141718 215863 141770 215869
rect 144020 214406 144076 214415
rect 144020 214341 144076 214350
rect 144034 213263 144062 214341
rect 144022 213257 144074 213263
rect 144022 213199 144074 213205
rect 139990 213109 140042 213115
rect 139990 213051 140042 213057
rect 144020 210854 144076 210863
rect 144020 210789 144076 210798
rect 144034 210303 144062 210789
rect 144022 210297 144074 210303
rect 144022 210239 144074 210245
rect 144020 209078 144076 209087
rect 144020 209013 144076 209022
rect 144034 207417 144062 209013
rect 144022 207411 144074 207417
rect 144022 207353 144074 207359
rect 144980 203454 145036 203463
rect 144980 203389 145036 203398
rect 144994 201645 145022 203389
rect 144982 201639 145034 201645
rect 144982 201581 145034 201587
rect 144980 200642 145036 200651
rect 144980 200577 145036 200586
rect 144404 199458 144460 199467
rect 144404 199393 144460 199402
rect 144418 198759 144446 199393
rect 144994 198833 145022 200577
rect 144982 198827 145034 198833
rect 144982 198769 145034 198775
rect 144406 198753 144458 198759
rect 144406 198695 144458 198701
rect 145268 197682 145324 197691
rect 145268 197617 145324 197626
rect 144980 196202 145036 196211
rect 144980 196137 145036 196146
rect 47638 194535 47690 194541
rect 47638 194477 47690 194483
rect 144596 193982 144652 193991
rect 144596 193917 144652 193926
rect 43318 193499 43370 193505
rect 43318 193441 43370 193447
rect 144610 193135 144638 193917
rect 144598 193129 144650 193135
rect 144598 193071 144650 193077
rect 144308 192206 144364 192215
rect 144308 192141 144364 192150
rect 43126 191057 43178 191063
rect 43126 190999 43178 191005
rect 144322 190175 144350 192141
rect 144884 191022 144940 191031
rect 144884 190957 144940 190966
rect 144310 190169 144362 190175
rect 144310 190111 144362 190117
rect 42658 188168 42974 188196
rect 42658 187141 42686 188168
rect 42742 187875 42794 187881
rect 42742 187817 42794 187823
rect 42646 187135 42698 187141
rect 42646 187077 42698 187083
rect 42070 186691 42122 186697
rect 42070 186633 42122 186639
rect 42454 186691 42506 186697
rect 42454 186633 42506 186639
rect 42082 186184 42110 186633
rect 41780 185990 41836 185999
rect 41780 185925 41836 185934
rect 41794 185592 41822 185925
rect 41780 184214 41836 184223
rect 41780 184149 41836 184158
rect 41794 183742 41822 184149
rect 41780 183622 41836 183631
rect 41780 183557 41836 183566
rect 41794 183121 41822 183557
rect 41780 182882 41836 182891
rect 41780 182817 41836 182826
rect 41794 182484 41822 182817
rect 42754 177119 42782 187817
rect 144692 182734 144748 182743
rect 144692 182669 144748 182678
rect 144706 181591 144734 182669
rect 144694 181585 144746 181591
rect 144694 181527 144746 181533
rect 144898 181369 144926 190957
rect 144994 182923 145022 196137
rect 145172 187470 145228 187479
rect 145172 187405 145228 187414
rect 145076 184362 145132 184371
rect 145076 184297 145132 184306
rect 144982 182917 145034 182923
rect 144982 182859 145034 182865
rect 144886 181363 144938 181369
rect 144886 181305 144938 181311
rect 144884 180810 144940 180819
rect 144884 180745 144940 180754
rect 144020 179182 144076 179191
rect 144020 179117 144076 179126
rect 144034 178631 144062 179117
rect 144022 178625 144074 178631
rect 144022 178567 144074 178573
rect 144692 177850 144748 177859
rect 144692 177785 144748 177794
rect 42740 177110 42796 177119
rect 42740 177045 42796 177054
rect 144500 177110 144556 177119
rect 144500 177045 144556 177054
rect 144404 172374 144460 172383
rect 144404 172309 144460 172318
rect 144020 164678 144076 164687
rect 144020 164613 144076 164622
rect 144034 164201 144062 164613
rect 144022 164195 144074 164201
rect 144022 164137 144074 164143
rect 144308 163938 144364 163947
rect 144308 163873 144364 163882
rect 144212 162162 144268 162171
rect 144212 162097 144268 162106
rect 144226 161315 144254 162097
rect 144322 161463 144350 163873
rect 144310 161457 144362 161463
rect 144310 161399 144362 161405
rect 144214 161309 144266 161315
rect 144214 161251 144266 161257
rect 144308 160386 144364 160395
rect 144308 160321 144364 160330
rect 144116 158610 144172 158619
rect 144116 158545 144172 158554
rect 143926 139479 143978 139485
rect 143926 139421 143978 139427
rect 143938 138079 143966 139421
rect 144130 138172 144158 158545
rect 144322 158503 144350 160321
rect 144310 158497 144362 158503
rect 144310 158439 144362 158445
rect 144308 156242 144364 156251
rect 144308 156177 144364 156186
rect 144322 156061 144350 156177
rect 144310 156055 144362 156061
rect 144310 155997 144362 156003
rect 144212 155502 144268 155511
rect 144212 155437 144268 155446
rect 144226 149105 144254 155437
rect 144308 153726 144364 153735
rect 144308 153661 144364 153670
rect 144322 152731 144350 153661
rect 144310 152725 144362 152731
rect 144310 152667 144362 152673
rect 144308 150766 144364 150775
rect 144308 150701 144364 150710
rect 144322 149919 144350 150701
rect 144310 149913 144362 149919
rect 144310 149855 144362 149861
rect 144214 149099 144266 149105
rect 144214 149041 144266 149047
rect 144212 148990 144268 148999
rect 144212 148925 144268 148934
rect 144226 147107 144254 148925
rect 144308 147806 144364 147815
rect 144308 147741 144364 147750
rect 144214 147101 144266 147107
rect 144214 147043 144266 147049
rect 144322 147033 144350 147741
rect 144310 147027 144362 147033
rect 144310 146969 144362 146975
rect 144214 146953 144266 146959
rect 144214 146895 144266 146901
rect 144226 139485 144254 146895
rect 144308 145290 144364 145299
rect 144308 145225 144364 145234
rect 144322 144147 144350 145225
rect 144310 144141 144362 144147
rect 144310 144083 144362 144089
rect 144308 143514 144364 143523
rect 144308 143449 144364 143458
rect 144322 141187 144350 143449
rect 144310 141181 144362 141187
rect 144310 141123 144362 141129
rect 144308 140554 144364 140563
rect 144308 140489 144364 140498
rect 144214 139479 144266 139485
rect 144214 139421 144266 139427
rect 144212 139370 144268 139379
rect 144212 139305 144268 139314
rect 144226 138449 144254 139305
rect 144214 138443 144266 138449
rect 144214 138385 144266 138391
rect 144322 138375 144350 140489
rect 144310 138369 144362 138375
rect 144310 138311 144362 138317
rect 144418 138301 144446 172309
rect 144514 161167 144542 177045
rect 144596 170006 144652 170015
rect 144596 169941 144652 169950
rect 144502 161161 144554 161167
rect 144502 161103 144554 161109
rect 144500 157426 144556 157435
rect 144500 157361 144556 157370
rect 144514 155617 144542 157361
rect 144502 155611 144554 155617
rect 144502 155553 144554 155559
rect 144500 153134 144556 153143
rect 144500 153069 144556 153078
rect 144514 152805 144542 153069
rect 144502 152799 144554 152805
rect 144502 152741 144554 152747
rect 144500 151950 144556 151959
rect 144500 151885 144556 151894
rect 144514 149845 144542 151885
rect 144502 149839 144554 149845
rect 144502 149781 144554 149787
rect 144502 149099 144554 149105
rect 144502 149041 144554 149047
rect 144514 147181 144542 149041
rect 144502 147175 144554 147181
rect 144502 147117 144554 147123
rect 144500 147066 144556 147075
rect 144500 147001 144556 147010
rect 144514 146959 144542 147001
rect 144502 146953 144554 146959
rect 144502 146895 144554 146901
rect 144500 144402 144556 144411
rect 144500 144337 144556 144346
rect 144514 144073 144542 144337
rect 144502 144067 144554 144073
rect 144502 144009 144554 144015
rect 144500 142330 144556 142339
rect 144500 142265 144502 142274
rect 144554 142265 144556 142274
rect 144502 142233 144554 142239
rect 144500 138630 144556 138639
rect 144500 138565 144556 138574
rect 144514 138301 144542 138565
rect 144406 138295 144458 138301
rect 144406 138237 144458 138243
rect 144502 138295 144554 138301
rect 144502 138237 144554 138243
rect 144130 138144 144542 138172
rect 143926 138073 143978 138079
rect 143926 138015 143978 138021
rect 144310 138073 144362 138079
rect 144310 138015 144362 138021
rect 144406 138073 144458 138079
rect 144406 138015 144458 138021
rect 144212 137002 144268 137011
rect 144212 136937 144268 136946
rect 144116 135966 144172 135975
rect 144116 135901 144172 135910
rect 144130 135489 144158 135901
rect 144226 135563 144254 136937
rect 144214 135557 144266 135563
rect 144214 135499 144266 135505
rect 144118 135483 144170 135489
rect 144118 135425 144170 135431
rect 144116 135078 144172 135087
rect 144116 135013 144172 135022
rect 144020 132710 144076 132719
rect 144020 132645 144022 132654
rect 144074 132645 144076 132654
rect 144022 132613 144074 132619
rect 144130 132529 144158 135013
rect 144212 133894 144268 133903
rect 144212 133829 144268 133838
rect 144226 132603 144254 133829
rect 144214 132597 144266 132603
rect 144214 132539 144266 132545
rect 144118 132523 144170 132529
rect 144118 132465 144170 132471
rect 144116 130934 144172 130943
rect 144116 130869 144172 130878
rect 144130 129717 144158 130869
rect 144212 130194 144268 130203
rect 144212 130129 144268 130138
rect 144118 129711 144170 129717
rect 144118 129653 144170 129659
rect 144226 129643 144254 130129
rect 144214 129637 144266 129643
rect 144214 129579 144266 129585
rect 144116 128566 144172 128575
rect 144116 128501 144172 128510
rect 144130 126831 144158 128501
rect 144212 127382 144268 127391
rect 144212 127317 144268 127326
rect 144118 126825 144170 126831
rect 144118 126767 144170 126773
rect 144226 126757 144254 127317
rect 144214 126751 144266 126757
rect 144214 126693 144266 126699
rect 144020 126642 144076 126651
rect 144020 126577 144076 126586
rect 144034 124019 144062 126577
rect 144212 125458 144268 125467
rect 144212 125393 144268 125402
rect 144116 124274 144172 124283
rect 144116 124209 144172 124218
rect 144022 124013 144074 124019
rect 144022 123955 144074 123961
rect 144130 123945 144158 124209
rect 144226 124093 144254 125393
rect 144214 124087 144266 124093
rect 144214 124029 144266 124035
rect 144118 123939 144170 123945
rect 144118 123881 144170 123887
rect 144212 121906 144268 121915
rect 144212 121841 144268 121850
rect 144226 121059 144254 121841
rect 144214 121053 144266 121059
rect 144214 120995 144266 121001
rect 144116 120130 144172 120139
rect 144116 120065 144172 120074
rect 144020 118946 144076 118955
rect 144020 118881 144076 118890
rect 144034 118173 144062 118881
rect 144130 118247 144158 120065
rect 144214 118315 144266 118321
rect 144214 118257 144266 118263
rect 144118 118241 144170 118247
rect 144226 118215 144254 118257
rect 144118 118183 144170 118189
rect 144212 118206 144268 118215
rect 144022 118167 144074 118173
rect 144212 118141 144268 118150
rect 144022 118109 144074 118115
rect 144116 117022 144172 117031
rect 144116 116957 144172 116966
rect 144130 115287 144158 116957
rect 144212 115542 144268 115551
rect 144212 115477 144268 115486
rect 144226 115361 144254 115477
rect 144214 115355 144266 115361
rect 144214 115297 144266 115303
rect 144118 115281 144170 115287
rect 144118 115223 144170 115229
rect 144116 114210 144172 114219
rect 144116 114145 144172 114154
rect 144130 112401 144158 114145
rect 144212 113470 144268 113479
rect 144212 113405 144268 113414
rect 144226 112475 144254 113405
rect 144214 112469 144266 112475
rect 144214 112411 144266 112417
rect 144118 112395 144170 112401
rect 144118 112337 144170 112343
rect 144020 111694 144076 111703
rect 144020 111629 144076 111638
rect 144034 109589 144062 111629
rect 144116 110510 144172 110519
rect 144116 110445 144172 110454
rect 144022 109583 144074 109589
rect 144022 109525 144074 109531
rect 144130 109515 144158 110445
rect 144212 109770 144268 109779
rect 144212 109705 144268 109714
rect 144226 109663 144254 109705
rect 144214 109657 144266 109663
rect 144214 109599 144266 109605
rect 144118 109509 144170 109515
rect 144118 109451 144170 109457
rect 144212 106958 144268 106967
rect 144212 106893 144268 106902
rect 144226 106629 144254 106893
rect 144214 106623 144266 106629
rect 144214 106565 144266 106571
rect 144020 105774 144076 105783
rect 144020 105709 144076 105718
rect 144034 103743 144062 105709
rect 144116 105034 144172 105043
rect 144116 104969 144172 104978
rect 144130 103891 144158 104969
rect 144118 103885 144170 103891
rect 144118 103827 144170 103833
rect 144212 103850 144268 103859
rect 144212 103785 144214 103794
rect 144266 103785 144268 103794
rect 144214 103753 144266 103759
rect 144022 103737 144074 103743
rect 144022 103679 144074 103685
rect 144212 102074 144268 102083
rect 144212 102009 144268 102018
rect 144226 100857 144254 102009
rect 144214 100851 144266 100857
rect 144214 100793 144266 100799
rect 144212 100150 144268 100159
rect 144212 100085 144268 100094
rect 144226 97971 144254 100085
rect 144214 97965 144266 97971
rect 144214 97907 144266 97913
rect 144116 97338 144172 97347
rect 144116 97273 144172 97282
rect 144020 95414 144076 95423
rect 144020 95349 144076 95358
rect 143924 92306 143980 92315
rect 143924 92241 143980 92250
rect 143938 75031 143966 92241
rect 144034 75253 144062 95349
rect 144130 95159 144158 97273
rect 144212 96598 144268 96607
rect 144212 96533 144268 96542
rect 144118 95153 144170 95159
rect 144118 95095 144170 95101
rect 144226 95085 144254 96533
rect 144214 95079 144266 95085
rect 144214 95021 144266 95027
rect 144212 93638 144268 93647
rect 144212 93573 144214 93582
rect 144266 93573 144268 93582
rect 144214 93541 144266 93547
rect 144116 91862 144172 91871
rect 144116 91797 144172 91806
rect 144130 88296 144158 91797
rect 144212 90678 144268 90687
rect 144212 90613 144214 90622
rect 144266 90613 144268 90622
rect 144214 90581 144266 90587
rect 144212 89346 144268 89355
rect 144212 89281 144214 89290
rect 144266 89281 144268 89290
rect 144214 89249 144266 89255
rect 144130 88268 144254 88296
rect 144116 88162 144172 88171
rect 144116 88097 144172 88106
rect 144130 86575 144158 88097
rect 144226 87093 144254 88268
rect 144214 87087 144266 87093
rect 144214 87029 144266 87035
rect 144212 86978 144268 86987
rect 144212 86913 144268 86922
rect 144118 86569 144170 86575
rect 144118 86511 144170 86517
rect 144226 86501 144254 86913
rect 144214 86495 144266 86501
rect 144214 86437 144266 86443
rect 144118 86421 144170 86427
rect 144118 86363 144170 86369
rect 144130 85336 144158 86363
rect 144130 85308 144254 85336
rect 144116 85202 144172 85211
rect 144116 85137 144172 85146
rect 144130 83689 144158 85137
rect 144118 83683 144170 83689
rect 144118 83625 144170 83631
rect 144116 83426 144172 83435
rect 144116 83361 144172 83370
rect 144130 80729 144158 83361
rect 144118 80723 144170 80729
rect 144118 80665 144170 80671
rect 144116 79726 144172 79735
rect 144116 79661 144172 79670
rect 144130 77917 144158 79661
rect 144226 78657 144254 85308
rect 144214 78651 144266 78657
rect 144214 78593 144266 78599
rect 144212 78542 144268 78551
rect 144212 78477 144268 78486
rect 144118 77911 144170 77917
rect 144118 77853 144170 77859
rect 144226 77843 144254 78477
rect 144214 77837 144266 77843
rect 144214 77779 144266 77785
rect 144118 77763 144170 77769
rect 144118 77705 144170 77711
rect 144022 75247 144074 75253
rect 144022 75189 144074 75195
rect 144130 75124 144158 77705
rect 144212 77358 144268 77367
rect 144212 77293 144214 77302
rect 144266 77293 144268 77302
rect 144214 77261 144266 77267
rect 144212 75878 144268 75887
rect 144212 75813 144268 75822
rect 144226 75401 144254 75813
rect 144214 75395 144266 75401
rect 144214 75337 144266 75343
rect 144214 75247 144266 75253
rect 144214 75189 144266 75195
rect 144034 75096 144158 75124
rect 143926 75025 143978 75031
rect 143926 74967 143978 74973
rect 143924 73806 143980 73815
rect 143924 73741 143926 73750
rect 143978 73741 143980 73750
rect 143926 73709 143978 73715
rect 143924 72178 143980 72187
rect 143924 72113 143980 72122
rect 143938 72071 143966 72113
rect 143926 72065 143978 72071
rect 143926 72007 143978 72013
rect 143828 68330 143884 68339
rect 143828 68265 143884 68274
rect 143842 66299 143870 68265
rect 143924 67146 143980 67155
rect 143924 67081 143980 67090
rect 143938 66965 143966 67081
rect 143926 66959 143978 66965
rect 143926 66901 143978 66907
rect 143924 66850 143980 66859
rect 143924 66785 143926 66794
rect 143978 66785 143980 66794
rect 143926 66753 143978 66759
rect 143830 66293 143882 66299
rect 143830 66235 143882 66241
rect 143924 64778 143980 64787
rect 143924 64713 143980 64722
rect 143938 63413 143966 64713
rect 143926 63407 143978 63413
rect 143926 63349 143978 63355
rect 138166 60521 138218 60527
rect 138166 60463 138218 60469
rect 138178 40219 138206 60463
rect 143924 54714 143980 54723
rect 143924 54649 143980 54658
rect 143938 51277 143966 54649
rect 143926 51271 143978 51277
rect 143926 51213 143978 51219
rect 144034 49871 144062 75096
rect 144118 75025 144170 75031
rect 144118 74967 144170 74973
rect 144130 49945 144158 74967
rect 144226 54723 144254 75189
rect 144212 54714 144268 54723
rect 144212 54649 144268 54658
rect 144118 49939 144170 49945
rect 144118 49881 144170 49887
rect 144022 49865 144074 49871
rect 144022 49807 144074 49813
rect 144322 49797 144350 138015
rect 144418 51129 144446 138015
rect 144406 51123 144458 51129
rect 144406 51065 144458 51071
rect 144310 49791 144362 49797
rect 144310 49733 144362 49739
rect 144514 49575 144542 138144
rect 144610 51055 144638 169941
rect 144598 51049 144650 51055
rect 144598 50991 144650 50997
rect 144706 50241 144734 177785
rect 144788 173558 144844 173567
rect 144788 173493 144844 173502
rect 144802 50981 144830 173493
rect 144898 161260 144926 180745
rect 144980 175926 145036 175935
rect 144980 175861 145036 175870
rect 144994 175819 145022 175861
rect 144982 175813 145034 175819
rect 144982 175755 145034 175761
rect 144980 174298 145036 174307
rect 144980 174233 145036 174242
rect 144994 172859 145022 174233
rect 144982 172853 145034 172859
rect 144982 172795 145034 172801
rect 144980 170598 145036 170607
rect 144980 170533 145036 170542
rect 144994 169973 145022 170533
rect 144982 169967 145034 169973
rect 144982 169909 145034 169915
rect 144980 168674 145036 168683
rect 144980 168609 145036 168618
rect 144994 167901 145022 168609
rect 144982 167895 145034 167901
rect 144982 167837 145034 167843
rect 144980 167194 145036 167203
rect 144980 167129 145036 167138
rect 144994 167087 145022 167129
rect 144982 167081 145034 167087
rect 144982 167023 145034 167029
rect 144980 165862 145036 165871
rect 144980 165797 145036 165806
rect 144994 164275 145022 165797
rect 144982 164269 145034 164275
rect 144982 164211 145034 164217
rect 144980 161570 145036 161579
rect 144980 161505 145036 161514
rect 144994 161389 145022 161505
rect 144982 161383 145034 161389
rect 144982 161325 145034 161331
rect 144898 161232 145022 161260
rect 144886 161161 144938 161167
rect 144886 161103 144938 161109
rect 144790 50975 144842 50981
rect 144790 50917 144842 50923
rect 144694 50235 144746 50241
rect 144694 50177 144746 50183
rect 144898 50167 144926 161103
rect 144886 50161 144938 50167
rect 144886 50103 144938 50109
rect 144994 50093 145022 161232
rect 144982 50087 145034 50093
rect 144982 50029 145034 50035
rect 145090 50019 145118 184297
rect 145186 50759 145214 187405
rect 145174 50753 145226 50759
rect 145174 50695 145226 50701
rect 145282 50685 145310 197617
rect 145270 50679 145322 50685
rect 145270 50621 145322 50627
rect 145078 50013 145130 50019
rect 145078 49955 145130 49961
rect 145378 49649 145406 236097
rect 145460 232462 145516 232471
rect 145460 232397 145516 232406
rect 145366 49643 145418 49649
rect 145366 49585 145418 49591
rect 144502 49569 144554 49575
rect 144502 49511 144554 49517
rect 145474 49353 145502 232397
rect 146530 229987 146558 268181
rect 149122 260919 149150 275502
rect 150274 270095 150302 275502
rect 150262 270089 150314 270095
rect 150262 270031 150314 270037
rect 149686 268683 149738 268689
rect 149686 268625 149738 268631
rect 149398 263059 149450 263065
rect 149398 263001 149450 263007
rect 149410 262917 149438 263001
rect 149398 262911 149450 262917
rect 149398 262853 149450 262859
rect 149110 260913 149162 260919
rect 149110 260855 149162 260861
rect 146806 252847 146858 252853
rect 146806 252789 146858 252795
rect 146818 241901 146846 252789
rect 146902 252773 146954 252779
rect 146902 252715 146954 252721
rect 146806 241895 146858 241901
rect 146806 241837 146858 241843
rect 146914 239015 146942 252715
rect 148246 247741 148298 247747
rect 148246 247683 148298 247689
rect 146902 239009 146954 239015
rect 146902 238951 146954 238957
rect 147190 233237 147242 233243
rect 147190 233179 147242 233185
rect 147202 230431 147230 233179
rect 147190 230425 147242 230431
rect 147190 230367 147242 230373
rect 146518 229981 146570 229987
rect 146518 229923 146570 229929
rect 145556 227726 145612 227735
rect 145556 227661 145612 227670
rect 145570 51425 145598 227661
rect 145652 225950 145708 225959
rect 145652 225885 145708 225894
rect 145558 51419 145610 51425
rect 145558 51361 145610 51367
rect 145558 51271 145610 51277
rect 145558 51213 145610 51219
rect 145570 50315 145598 51213
rect 145558 50309 145610 50315
rect 145558 50251 145610 50257
rect 145462 49347 145514 49353
rect 145462 49289 145514 49295
rect 145666 49205 145694 225885
rect 145748 222842 145804 222851
rect 145748 222777 145804 222786
rect 145762 51351 145790 222777
rect 145844 219290 145900 219299
rect 145844 219225 145900 219234
rect 145750 51345 145802 51351
rect 145750 51287 145802 51293
rect 145858 51277 145886 219225
rect 145940 216330 145996 216339
rect 145940 216265 145996 216274
rect 145846 51271 145898 51277
rect 145846 51213 145898 51219
rect 145954 50907 145982 216265
rect 146516 215590 146572 215599
rect 146516 215525 146572 215534
rect 146036 213370 146092 213379
rect 146036 213305 146092 213314
rect 145942 50901 145994 50907
rect 145942 50843 145994 50849
rect 146050 50833 146078 213305
rect 146530 213189 146558 215525
rect 146518 213183 146570 213189
rect 146518 213125 146570 213131
rect 146132 211594 146188 211603
rect 146132 211529 146188 211538
rect 146038 50827 146090 50833
rect 146038 50769 146090 50775
rect 146146 49723 146174 211529
rect 146228 207894 146284 207903
rect 146228 207829 146284 207838
rect 146134 49717 146186 49723
rect 146134 49659 146186 49665
rect 146242 49501 146270 207829
rect 148054 207411 148106 207417
rect 148054 207353 148106 207359
rect 146804 207154 146860 207163
rect 146804 207089 146860 207098
rect 146324 206118 146380 206127
rect 146324 206053 146380 206062
rect 146230 49495 146282 49501
rect 146230 49437 146282 49443
rect 146338 49279 146366 206053
rect 146818 205197 146846 207089
rect 146806 205191 146858 205197
rect 146806 205133 146858 205139
rect 146804 204934 146860 204943
rect 146804 204869 146860 204878
rect 146818 204531 146846 204869
rect 146806 204525 146858 204531
rect 146806 204467 146858 204473
rect 146420 202418 146476 202427
rect 146420 202353 146476 202362
rect 146434 51203 146462 202353
rect 146708 198718 146764 198727
rect 146708 198653 146764 198662
rect 146516 190430 146572 190439
rect 146516 190365 146572 190374
rect 146530 183016 146558 190365
rect 146612 186286 146668 186295
rect 146612 186221 146668 186230
rect 146626 184403 146654 186221
rect 146614 184397 146666 184403
rect 146614 184339 146666 184345
rect 146530 182988 146654 183016
rect 146518 182917 146570 182923
rect 146518 182859 146570 182865
rect 146422 51197 146474 51203
rect 146422 51139 146474 51145
rect 146530 50611 146558 182859
rect 146518 50605 146570 50611
rect 146518 50547 146570 50553
rect 146626 50537 146654 182988
rect 146614 50531 146666 50537
rect 146614 50473 146666 50479
rect 146722 50463 146750 198653
rect 146804 194722 146860 194731
rect 146804 194657 146860 194666
rect 146818 193061 146846 194657
rect 146806 193055 146858 193061
rect 146806 192997 146858 193003
rect 146804 189246 146860 189255
rect 146804 189181 146860 189190
rect 146818 187289 146846 189181
rect 146806 187283 146858 187289
rect 146806 187225 146858 187231
rect 146804 185546 146860 185555
rect 146804 185481 146860 185490
rect 146818 184477 146846 185481
rect 146806 184471 146858 184477
rect 146806 184413 146858 184419
rect 146804 181994 146860 182003
rect 146804 181929 146860 181938
rect 146818 181517 146846 181929
rect 146806 181511 146858 181517
rect 146806 181453 146858 181459
rect 146806 181363 146858 181369
rect 146806 181305 146858 181311
rect 146710 50457 146762 50463
rect 146710 50399 146762 50405
rect 146818 50389 146846 181305
rect 147958 158497 148010 158503
rect 147958 158439 148010 158445
rect 147862 147101 147914 147107
rect 147862 147043 147914 147049
rect 147766 144141 147818 144147
rect 147766 144083 147818 144089
rect 147670 132671 147722 132677
rect 147670 132613 147722 132619
rect 147476 122498 147532 122507
rect 147476 122433 147532 122442
rect 147380 100890 147436 100899
rect 147380 100825 147436 100834
rect 147284 98522 147340 98531
rect 147284 98457 147340 98466
rect 146900 83870 146956 83879
rect 146900 83805 146902 83814
rect 146954 83805 146956 83814
rect 146902 83773 146954 83779
rect 146902 83535 146954 83541
rect 146902 83477 146954 83483
rect 146914 81067 146942 83477
rect 146996 82242 147052 82251
rect 146996 82177 146998 82186
rect 147050 82177 147052 82186
rect 146998 82145 147050 82151
rect 146900 81058 146956 81067
rect 146900 80993 146956 81002
rect 146900 74990 146956 74999
rect 146900 74925 146902 74934
rect 146954 74925 146956 74934
rect 146902 74893 146954 74899
rect 146996 71290 147052 71299
rect 146996 71225 147052 71234
rect 146900 70106 146956 70115
rect 146900 70041 146902 70050
rect 146954 70041 146956 70050
rect 146902 70009 146954 70015
rect 146900 64186 146956 64195
rect 146900 64121 146902 64130
rect 146954 64121 146956 64130
rect 146902 64089 146954 64095
rect 147010 63339 147038 71225
rect 147298 66151 147326 98457
rect 147394 66225 147422 100825
rect 147490 69111 147518 122433
rect 147572 108586 147628 108595
rect 147572 108521 147628 108530
rect 147478 69105 147530 69111
rect 147478 69047 147530 69053
rect 147382 66219 147434 66225
rect 147382 66161 147434 66167
rect 147286 66145 147338 66151
rect 147286 66087 147338 66093
rect 146998 63333 147050 63339
rect 146998 63275 147050 63281
rect 146996 62262 147052 62271
rect 146996 62197 147052 62206
rect 146900 61226 146956 61235
rect 146900 61161 146956 61170
rect 146914 60675 146942 61161
rect 146902 60669 146954 60675
rect 146902 60611 146954 60617
rect 147010 60601 147038 62197
rect 146998 60595 147050 60601
rect 146998 60537 147050 60543
rect 146806 50383 146858 50389
rect 146806 50325 146858 50331
rect 146326 49273 146378 49279
rect 146326 49215 146378 49221
rect 145654 49199 145706 49205
rect 145654 49141 145706 49147
rect 147586 48169 147614 108521
rect 147682 48243 147710 132613
rect 147670 48237 147722 48243
rect 147670 48179 147722 48185
rect 147574 48163 147626 48169
rect 147574 48105 147626 48111
rect 147778 46245 147806 144083
rect 147874 46541 147902 147043
rect 147862 46535 147914 46541
rect 147862 46477 147914 46483
rect 147970 46393 147998 158439
rect 148066 47767 148094 207353
rect 148150 161457 148202 161463
rect 148150 161399 148202 161405
rect 148162 48021 148190 161399
rect 148258 48655 148286 247683
rect 148438 244929 148490 244935
rect 148438 244871 148490 244877
rect 148342 213183 148394 213189
rect 148342 213125 148394 213131
rect 148244 48646 148300 48655
rect 148244 48581 148300 48590
rect 148150 48015 148202 48021
rect 148150 47957 148202 47963
rect 148052 47758 148108 47767
rect 148052 47693 148108 47702
rect 148354 47429 148382 213125
rect 148450 48507 148478 244871
rect 149590 244485 149642 244491
rect 149590 244427 149642 244433
rect 148630 241969 148682 241975
rect 148630 241911 148682 241917
rect 148534 193129 148586 193135
rect 148534 193071 148586 193077
rect 148436 48498 148492 48507
rect 148436 48433 148492 48442
rect 148546 47725 148574 193071
rect 148642 48359 148670 241911
rect 149602 239163 149630 244427
rect 149590 239157 149642 239163
rect 149590 239099 149642 239105
rect 148822 236567 148874 236573
rect 148822 236509 148874 236515
rect 148726 229019 148778 229025
rect 148726 228961 148778 228967
rect 148738 83541 148766 228961
rect 148726 83535 148778 83541
rect 148726 83477 148778 83483
rect 148628 48350 148684 48359
rect 148628 48285 148684 48294
rect 148534 47719 148586 47725
rect 148534 47661 148586 47667
rect 148834 47619 148862 236509
rect 149206 233385 149258 233391
rect 149206 233327 149258 233333
rect 148918 181585 148970 181591
rect 148918 181527 148970 181533
rect 148930 47651 148958 181527
rect 149014 175813 149066 175819
rect 149014 175755 149066 175761
rect 149026 77695 149054 175755
rect 149110 156055 149162 156061
rect 149110 155997 149162 156003
rect 149122 77769 149150 155997
rect 149110 77763 149162 77769
rect 149110 77705 149162 77711
rect 149014 77689 149066 77695
rect 149014 77631 149066 77637
rect 149218 48211 149246 233327
rect 149398 227687 149450 227693
rect 149398 227629 149450 227635
rect 149302 172853 149354 172859
rect 149302 172795 149354 172801
rect 149204 48202 149260 48211
rect 149204 48137 149260 48146
rect 148918 47645 148970 47651
rect 148820 47610 148876 47619
rect 148918 47587 148970 47593
rect 148820 47545 148876 47554
rect 148342 47423 148394 47429
rect 148342 47365 148394 47371
rect 149314 46689 149342 172795
rect 149410 48063 149438 227629
rect 149590 219029 149642 219035
rect 149590 218971 149642 218977
rect 149494 167081 149546 167087
rect 149494 167023 149546 167029
rect 149396 48054 149452 48063
rect 149396 47989 149452 47998
rect 149506 46837 149534 167023
rect 149602 47915 149630 218971
rect 149698 218665 149726 268625
rect 151426 267949 151454 275502
rect 152578 270169 152606 275502
rect 152566 270163 152618 270169
rect 152566 270105 152618 270111
rect 151414 267943 151466 267949
rect 151414 267885 151466 267891
rect 152566 267943 152618 267949
rect 152566 267885 152618 267891
rect 151126 242043 151178 242049
rect 151126 241985 151178 241991
rect 149782 239009 149834 239015
rect 149782 238951 149834 238957
rect 149794 230357 149822 238951
rect 149782 230351 149834 230357
rect 149782 230293 149834 230299
rect 149686 218659 149738 218665
rect 149686 218601 149738 218607
rect 149686 164269 149738 164275
rect 149686 164211 149738 164217
rect 149588 47906 149644 47915
rect 149588 47841 149644 47850
rect 149494 46831 149546 46837
rect 149494 46773 149546 46779
rect 149698 46763 149726 164211
rect 149782 93599 149834 93605
rect 149782 93541 149834 93547
rect 149794 77621 149822 93541
rect 151138 92125 151166 241985
rect 152086 241895 152138 241901
rect 152086 241837 152138 241843
rect 152098 230283 152126 241837
rect 152086 230277 152138 230283
rect 152086 230219 152138 230225
rect 152578 230061 152606 267885
rect 153826 258255 153854 275502
rect 154992 275488 155486 275516
rect 153814 258249 153866 258255
rect 153814 258191 153866 258197
rect 155350 239157 155402 239163
rect 155350 239099 155402 239105
rect 155362 230653 155390 239099
rect 155350 230647 155402 230653
rect 155350 230589 155402 230595
rect 152566 230055 152618 230061
rect 152566 229997 152618 230003
rect 155458 218591 155486 275488
rect 156226 260179 156254 275502
rect 157378 270243 157406 275502
rect 158626 270687 158654 275502
rect 158614 270681 158666 270687
rect 158614 270623 158666 270629
rect 159778 270391 159806 275502
rect 159766 270385 159818 270391
rect 159766 270327 159818 270333
rect 157366 270237 157418 270243
rect 157366 270179 157418 270185
rect 156214 260173 156266 260179
rect 156214 260115 156266 260121
rect 161026 258329 161054 275502
rect 162178 270687 162206 275502
rect 161206 270681 161258 270687
rect 161206 270623 161258 270629
rect 162166 270681 162218 270687
rect 162166 270623 162218 270629
rect 161014 258323 161066 258329
rect 161014 258265 161066 258271
rect 156886 230647 156938 230653
rect 156886 230589 156938 230595
rect 156898 228623 156926 230589
rect 161218 230135 161246 270623
rect 163426 270317 163454 275502
rect 164086 270681 164138 270687
rect 164086 270623 164138 270629
rect 163414 270311 163466 270317
rect 163414 270253 163466 270259
rect 161206 230129 161258 230135
rect 161206 230071 161258 230077
rect 156884 228614 156940 228623
rect 156884 228549 156940 228558
rect 155446 218585 155498 218591
rect 155446 218527 155498 218533
rect 159766 218067 159818 218073
rect 159766 218009 159818 218015
rect 154006 213257 154058 213263
rect 154006 213199 154058 213205
rect 151222 169967 151274 169973
rect 151222 169909 151274 169915
rect 151126 92119 151178 92125
rect 151126 92061 151178 92067
rect 151234 86427 151262 169909
rect 151318 138443 151370 138449
rect 151318 138385 151370 138391
rect 151222 86421 151274 86427
rect 151222 86363 151274 86369
rect 149782 77615 149834 77621
rect 149782 77557 149834 77563
rect 151126 74951 151178 74957
rect 151126 74893 151178 74899
rect 151138 63265 151166 74893
rect 151330 71701 151358 138385
rect 152662 92193 152714 92199
rect 152662 92135 152714 92141
rect 151318 71695 151370 71701
rect 151318 71637 151370 71643
rect 152674 65411 152702 92135
rect 154018 86353 154046 213199
rect 156886 205191 156938 205197
rect 156886 205133 156938 205139
rect 154102 149913 154154 149919
rect 154102 149855 154154 149861
rect 154006 86347 154058 86353
rect 154006 86289 154058 86295
rect 154114 74883 154142 149855
rect 156898 92051 156926 205133
rect 156982 167895 157034 167901
rect 156982 167837 157034 167843
rect 156886 92045 156938 92051
rect 156886 91987 156938 91993
rect 156994 83245 157022 167837
rect 157078 142291 157130 142297
rect 157078 142233 157130 142239
rect 156982 83239 157034 83245
rect 156982 83181 157034 83187
rect 155542 77319 155594 77325
rect 155542 77261 155594 77267
rect 154102 74877 154154 74883
rect 154102 74819 154154 74825
rect 152662 65405 152714 65411
rect 152662 65347 152714 65353
rect 155158 65405 155210 65411
rect 155158 65347 155210 65353
rect 151126 63259 151178 63265
rect 151126 63201 151178 63207
rect 155170 52184 155198 65347
rect 155554 63191 155582 77261
rect 157090 74809 157118 142233
rect 159778 86279 159806 218009
rect 164098 215853 164126 270623
rect 164578 270465 164606 275502
rect 165826 270687 165854 275502
rect 165814 270681 165866 270687
rect 165814 270623 165866 270629
rect 164566 270459 164618 270465
rect 164566 270401 164618 270407
rect 166882 269207 166910 275502
rect 166966 270681 167018 270687
rect 166966 270623 167018 270629
rect 166870 269201 166922 269207
rect 166870 269143 166922 269149
rect 166978 230209 167006 270623
rect 168034 261807 168062 275502
rect 169296 275488 169886 275516
rect 168022 261801 168074 261807
rect 168022 261743 168074 261749
rect 168406 233311 168458 233317
rect 168406 233253 168458 233259
rect 166966 230203 167018 230209
rect 166966 230145 167018 230151
rect 165526 218955 165578 218961
rect 165526 218897 165578 218903
rect 164086 215847 164138 215853
rect 164086 215789 164138 215795
rect 162646 198827 162698 198833
rect 162646 198769 162698 198775
rect 159862 152799 159914 152805
rect 159862 152741 159914 152747
rect 159766 86273 159818 86279
rect 159766 86215 159818 86221
rect 159766 75395 159818 75401
rect 159766 75337 159818 75343
rect 157078 74803 157130 74809
rect 157078 74745 157130 74751
rect 155542 63185 155594 63191
rect 155542 63127 155594 63133
rect 159094 60521 159146 60527
rect 159094 60463 159146 60469
rect 159106 56476 159134 60463
rect 159072 56448 159134 56476
rect 159778 52480 159806 75337
rect 159874 74661 159902 152741
rect 160246 90639 160298 90645
rect 160246 90581 160298 90587
rect 160054 82203 160106 82209
rect 160054 82145 160106 82151
rect 159862 74655 159914 74661
rect 159862 74597 159914 74603
rect 159958 73767 160010 73773
rect 159958 73709 160010 73715
rect 159862 70067 159914 70073
rect 159862 70009 159914 70015
rect 159874 52628 159902 70009
rect 159970 52757 159998 73709
rect 160066 63117 160094 82145
rect 160258 74735 160286 90581
rect 162658 86205 162686 198769
rect 162742 147027 162794 147033
rect 162742 146969 162794 146975
rect 162646 86199 162698 86205
rect 162646 86141 162698 86147
rect 162646 80723 162698 80729
rect 162646 80665 162698 80671
rect 160246 74729 160298 74735
rect 160246 74671 160298 74677
rect 160150 72065 160202 72071
rect 160150 72007 160202 72013
rect 160054 63111 160106 63117
rect 160054 63053 160106 63059
rect 160162 52905 160190 72007
rect 160246 66959 160298 66965
rect 160246 66901 160298 66907
rect 160258 53053 160286 66901
rect 160342 66811 160394 66817
rect 160342 66753 160394 66759
rect 160354 53201 160382 66753
rect 160438 64147 160490 64153
rect 160438 64089 160490 64095
rect 160450 53349 160478 64089
rect 160534 60669 160586 60675
rect 160534 60611 160586 60617
rect 160438 53343 160490 53349
rect 160438 53285 160490 53291
rect 160342 53195 160394 53201
rect 160342 53137 160394 53143
rect 160246 53047 160298 53053
rect 160246 52989 160298 52995
rect 160150 52899 160202 52905
rect 160150 52841 160202 52847
rect 159958 52751 160010 52757
rect 159958 52693 160010 52699
rect 160546 52683 160574 60611
rect 160534 52677 160586 52683
rect 159874 52609 159998 52628
rect 160534 52619 160586 52625
rect 159874 52603 160010 52609
rect 159874 52600 159958 52603
rect 159958 52545 160010 52551
rect 162658 52535 162686 80665
rect 162646 52529 162698 52535
rect 159778 52452 159998 52480
rect 162646 52471 162698 52477
rect 155170 52156 155424 52184
rect 159970 52017 159998 52452
rect 162754 52165 162782 146969
rect 163030 146953 163082 146959
rect 163030 146895 163082 146901
rect 162838 144067 162890 144073
rect 162838 144009 162890 144015
rect 162850 52313 162878 144009
rect 162934 138369 162986 138375
rect 162934 138311 162986 138317
rect 162946 52461 162974 138311
rect 163042 74587 163070 146895
rect 163126 89307 163178 89313
rect 163126 89249 163178 89255
rect 163030 74581 163082 74587
rect 163030 74523 163082 74529
rect 162934 52455 162986 52461
rect 162934 52397 162986 52403
rect 162838 52307 162890 52313
rect 162838 52249 162890 52255
rect 163138 52239 163166 89249
rect 163222 86569 163274 86575
rect 163222 86511 163274 86517
rect 163234 52387 163262 86511
rect 165538 86131 165566 218897
rect 165622 155611 165674 155617
rect 165622 155553 165674 155559
rect 165526 86125 165578 86131
rect 165526 86067 165578 86073
rect 163606 83831 163658 83837
rect 163606 83773 163658 83779
rect 163318 83683 163370 83689
rect 163318 83625 163370 83631
rect 163330 52831 163358 83625
rect 163414 77911 163466 77917
rect 163414 77853 163466 77859
rect 163426 52979 163454 77853
rect 163510 77837 163562 77843
rect 163510 77779 163562 77785
rect 163522 53497 163550 77779
rect 163618 63043 163646 83773
rect 165634 77547 165662 155553
rect 165718 103885 165770 103891
rect 165718 103827 165770 103833
rect 165622 77541 165674 77547
rect 165622 77483 165674 77489
rect 165730 66077 165758 103827
rect 168418 89239 168446 233253
rect 169858 228951 169886 275488
rect 170434 261067 170462 275502
rect 171682 269133 171710 275502
rect 172834 270687 172862 275502
rect 172822 270681 172874 270687
rect 172822 270623 172874 270629
rect 174082 270539 174110 275502
rect 174070 270533 174122 270539
rect 174070 270475 174122 270481
rect 171670 269127 171722 269133
rect 171670 269069 171722 269075
rect 175234 261881 175262 275502
rect 176482 270687 176510 275502
rect 175606 270681 175658 270687
rect 175606 270623 175658 270629
rect 176470 270681 176522 270687
rect 176470 270623 176522 270629
rect 175222 261875 175274 261881
rect 175222 261817 175274 261823
rect 170422 261061 170474 261067
rect 170422 261003 170474 261009
rect 169846 228945 169898 228951
rect 169846 228887 169898 228893
rect 174166 224727 174218 224733
rect 174166 224669 174218 224675
rect 171286 221841 171338 221847
rect 171286 221783 171338 221789
rect 168502 181511 168554 181517
rect 168502 181453 168554 181459
rect 168406 89233 168458 89239
rect 168406 89175 168458 89181
rect 168514 80655 168542 181453
rect 168598 115355 168650 115361
rect 168598 115297 168650 115303
rect 168502 80649 168554 80655
rect 168502 80591 168554 80597
rect 168610 69037 168638 115297
rect 171298 86057 171326 221783
rect 171382 161383 171434 161389
rect 171382 161325 171434 161331
rect 171286 86051 171338 86057
rect 171286 85993 171338 85999
rect 171394 77473 171422 161325
rect 171478 106623 171530 106629
rect 171478 106565 171530 106571
rect 171382 77467 171434 77473
rect 171382 77409 171434 77415
rect 168598 69031 168650 69037
rect 168598 68973 168650 68979
rect 167062 66293 167114 66299
rect 167062 66235 167114 66241
rect 165718 66071 165770 66077
rect 165718 66013 165770 66019
rect 164278 63407 164330 63413
rect 164278 63349 164330 63355
rect 163606 63037 163658 63043
rect 163606 62979 163658 62985
rect 164290 60379 164318 63349
rect 164278 60373 164330 60379
rect 164278 60315 164330 60321
rect 167074 60305 167102 66235
rect 171490 66003 171518 106565
rect 174178 89165 174206 224669
rect 175618 215779 175646 270623
rect 177634 261215 177662 275502
rect 178896 275488 179198 275516
rect 178486 270681 178538 270687
rect 178486 270623 178538 270629
rect 177622 261209 177674 261215
rect 177622 261151 177674 261157
rect 178498 228877 178526 270623
rect 179170 270539 179198 275488
rect 180034 270687 180062 275502
rect 180022 270681 180074 270687
rect 180022 270623 180074 270629
rect 179158 270533 179210 270539
rect 179158 270475 179210 270481
rect 181282 261141 181310 275502
rect 181556 273458 181612 273467
rect 181556 273393 181612 273402
rect 181570 273171 181598 273393
rect 181556 273162 181612 273171
rect 181556 273097 181612 273106
rect 181366 270681 181418 270687
rect 181366 270623 181418 270629
rect 181270 261135 181322 261141
rect 181270 261077 181322 261083
rect 178594 255813 178718 255832
rect 178582 255807 178730 255813
rect 178634 255804 178678 255807
rect 178582 255749 178634 255755
rect 178678 255749 178730 255755
rect 178486 228871 178538 228877
rect 178486 228813 178538 228819
rect 177046 227613 177098 227619
rect 177046 227555 177098 227561
rect 175606 215773 175658 215779
rect 175606 215715 175658 215721
rect 174262 161309 174314 161315
rect 174262 161251 174314 161257
rect 174166 89159 174218 89165
rect 174166 89101 174218 89107
rect 174274 77399 174302 161251
rect 174358 109657 174410 109663
rect 174358 109599 174410 109605
rect 174262 77393 174314 77399
rect 174262 77335 174314 77341
rect 171478 65997 171530 66003
rect 171478 65939 171530 65945
rect 174370 65929 174398 109599
rect 177058 89091 177086 227555
rect 181378 215705 181406 270623
rect 182434 267061 182462 275502
rect 183490 270687 183518 275502
rect 183478 270681 183530 270687
rect 183478 270623 183530 270629
rect 184246 270681 184298 270687
rect 184246 270623 184298 270629
rect 184342 270681 184394 270687
rect 184342 270623 184394 270629
rect 182422 267055 182474 267061
rect 182422 266997 182474 267003
rect 182326 250627 182378 250633
rect 182326 250569 182378 250575
rect 182338 247599 182366 250569
rect 182326 247593 182378 247599
rect 182326 247535 182378 247541
rect 184258 228803 184286 270623
rect 184354 269133 184382 270623
rect 184738 269133 184766 275502
rect 184342 269127 184394 269133
rect 184342 269069 184394 269075
rect 184726 269127 184778 269133
rect 184726 269069 184778 269075
rect 185890 261585 185918 275502
rect 185878 261579 185930 261585
rect 185878 261521 185930 261527
rect 184246 228797 184298 228803
rect 184246 228739 184298 228745
rect 181366 215699 181418 215705
rect 181366 215641 181418 215647
rect 187138 215631 187166 275502
rect 188290 268837 188318 275502
rect 189538 268985 189566 275502
rect 189526 268979 189578 268985
rect 189526 268921 189578 268927
rect 188278 268831 188330 268837
rect 188278 268773 188330 268779
rect 190690 268615 190718 275502
rect 190678 268609 190730 268615
rect 190678 268551 190730 268557
rect 191938 261511 191966 275502
rect 192886 268609 192938 268615
rect 192886 268551 192938 268557
rect 191926 261505 191978 261511
rect 191926 261447 191978 261453
rect 191446 247815 191498 247821
rect 191446 247757 191498 247763
rect 188566 239083 188618 239089
rect 188566 239025 188618 239031
rect 187126 215625 187178 215631
rect 187126 215567 187178 215573
rect 185686 210297 185738 210303
rect 185686 210239 185738 210245
rect 182806 204525 182858 204531
rect 182806 204467 182858 204473
rect 179926 201639 179978 201645
rect 179926 201581 179978 201587
rect 177142 178625 177194 178631
rect 177142 178567 177194 178573
rect 177046 89085 177098 89091
rect 177046 89027 177098 89033
rect 177154 80581 177182 178567
rect 177238 109583 177290 109589
rect 177238 109525 177290 109531
rect 177142 80575 177194 80581
rect 177142 80517 177194 80523
rect 174358 65923 174410 65929
rect 174358 65865 174410 65871
rect 177250 65855 177278 109525
rect 179938 89017 179966 201581
rect 180022 184471 180074 184477
rect 180022 184413 180074 184419
rect 179926 89011 179978 89017
rect 179926 88953 179978 88959
rect 180034 80507 180062 184413
rect 180118 118315 180170 118321
rect 180118 118257 180170 118263
rect 180022 80501 180074 80507
rect 180022 80443 180074 80449
rect 180130 68963 180158 118257
rect 182818 91829 182846 204467
rect 182902 184397 182954 184403
rect 182902 184339 182954 184345
rect 182806 91823 182858 91829
rect 182806 91765 182858 91771
rect 182914 80285 182942 184339
rect 182998 118241 183050 118247
rect 182998 118183 183050 118189
rect 182902 80279 182954 80285
rect 182902 80221 182954 80227
rect 180118 68957 180170 68963
rect 180118 68899 180170 68905
rect 183010 68815 183038 118183
rect 185698 91903 185726 210239
rect 185782 187283 185834 187289
rect 185782 187225 185834 187231
rect 185686 91897 185738 91903
rect 185686 91839 185738 91845
rect 185794 80433 185822 187225
rect 185878 124087 185930 124093
rect 185878 124029 185930 124035
rect 185782 80427 185834 80433
rect 185782 80369 185834 80375
rect 185890 68889 185918 124029
rect 188578 91977 188606 239025
rect 188662 190169 188714 190175
rect 188662 190111 188714 190117
rect 188566 91971 188618 91977
rect 188566 91913 188618 91919
rect 188674 83319 188702 190111
rect 188758 126825 188810 126831
rect 188758 126767 188810 126773
rect 188662 83313 188714 83319
rect 188662 83255 188714 83261
rect 188770 71775 188798 126767
rect 191458 94937 191486 247757
rect 192898 228655 192926 268551
rect 193090 261363 193118 275502
rect 194338 266543 194366 275502
rect 194326 266537 194378 266543
rect 194326 266479 194378 266485
rect 193078 261357 193130 261363
rect 193078 261299 193130 261305
rect 195490 261289 195518 275502
rect 196738 264101 196766 275502
rect 197890 264735 197918 275502
rect 197876 264726 197932 264735
rect 197876 264661 197932 264670
rect 196726 264095 196778 264101
rect 196726 264037 196778 264043
rect 199042 261437 199070 275502
rect 200194 264027 200222 275502
rect 201346 266469 201374 275502
rect 202594 269059 202622 275502
rect 202582 269053 202634 269059
rect 202582 268995 202634 269001
rect 201334 266463 201386 266469
rect 201334 266405 201386 266411
rect 200182 264021 200234 264027
rect 200182 263963 200234 263969
rect 203746 263879 203774 275502
rect 204310 269053 204362 269059
rect 204310 268995 204362 269001
rect 203734 263873 203786 263879
rect 203734 263815 203786 263821
rect 201622 261579 201674 261585
rect 201622 261521 201674 261527
rect 199030 261431 199082 261437
rect 199030 261373 199082 261379
rect 195478 261283 195530 261289
rect 195478 261225 195530 261231
rect 198740 260730 198796 260739
rect 198740 260665 198742 260674
rect 198794 260665 198796 260674
rect 198742 260633 198794 260639
rect 201634 258403 201662 261521
rect 201622 258397 201674 258403
rect 201622 258339 201674 258345
rect 200278 254919 200330 254925
rect 200278 254861 200330 254867
rect 200182 252625 200234 252631
rect 200182 252567 200234 252573
rect 200086 250035 200138 250041
rect 200086 249977 200138 249983
rect 197206 244855 197258 244861
rect 197206 244797 197258 244803
rect 194326 230499 194378 230505
rect 194326 230441 194378 230447
rect 192886 228649 192938 228655
rect 192886 228591 192938 228597
rect 191542 193055 191594 193061
rect 191542 192997 191594 193003
rect 191446 94931 191498 94937
rect 191446 94873 191498 94879
rect 191554 83393 191582 192997
rect 191638 129711 191690 129717
rect 191638 129653 191690 129659
rect 191542 83387 191594 83393
rect 191542 83329 191594 83335
rect 191650 71849 191678 129653
rect 194338 88943 194366 230441
rect 194422 164195 194474 164201
rect 194422 164137 194474 164143
rect 194326 88937 194378 88943
rect 194326 88879 194378 88885
rect 194434 83467 194462 164137
rect 194518 132597 194570 132603
rect 194518 132539 194570 132545
rect 194422 83461 194474 83467
rect 194422 83403 194474 83409
rect 194530 71923 194558 132539
rect 197218 95011 197246 244797
rect 200098 241920 200126 249977
rect 200002 241892 200126 241920
rect 200002 227619 200030 241892
rect 199990 227613 200042 227619
rect 199990 227555 200042 227561
rect 200086 227539 200138 227545
rect 200086 227481 200138 227487
rect 199796 222102 199852 222111
rect 199796 222037 199852 222046
rect 199700 221806 199756 221815
rect 198742 221767 198794 221773
rect 199700 221741 199756 221750
rect 198742 221709 198794 221715
rect 198754 219151 198782 221709
rect 198740 219142 198796 219151
rect 198740 219077 198796 219086
rect 199030 218881 199082 218887
rect 199030 218823 199082 218829
rect 198742 218807 198794 218813
rect 198742 218749 198794 218755
rect 198754 218707 198782 218749
rect 198838 218733 198890 218739
rect 198740 218698 198796 218707
rect 198838 218675 198890 218681
rect 198740 218633 198796 218642
rect 198742 218585 198794 218591
rect 198742 218527 198794 218533
rect 198754 216487 198782 218527
rect 198850 217523 198878 218675
rect 198934 218659 198986 218665
rect 198934 218601 198986 218607
rect 198836 217514 198892 217523
rect 198836 217449 198892 217458
rect 198946 217375 198974 218601
rect 199042 218115 199070 218823
rect 199028 218106 199084 218115
rect 199028 218041 199084 218050
rect 198932 217366 198988 217375
rect 198932 217301 198988 217310
rect 198740 216478 198796 216487
rect 198740 216413 198796 216422
rect 199030 215995 199082 216001
rect 199030 215937 199082 215943
rect 198934 215921 198986 215927
rect 198740 215886 198796 215895
rect 198934 215863 198986 215869
rect 198740 215821 198742 215830
rect 198794 215821 198796 215830
rect 198742 215789 198794 215795
rect 198838 215773 198890 215779
rect 198836 215738 198838 215747
rect 198890 215738 198892 215747
rect 198742 215699 198794 215705
rect 198836 215673 198892 215682
rect 198742 215641 198794 215647
rect 198754 214859 198782 215641
rect 198838 215625 198890 215631
rect 198838 215567 198890 215573
rect 198740 214850 198796 214859
rect 198740 214785 198796 214794
rect 198850 214267 198878 215567
rect 198836 214258 198892 214267
rect 198836 214193 198892 214202
rect 198946 214119 198974 215863
rect 198932 214110 198988 214119
rect 198932 214045 198988 214054
rect 199042 213231 199070 215937
rect 199028 213222 199084 213231
rect 199028 213157 199084 213166
rect 198742 213109 198794 213115
rect 198742 213051 198794 213057
rect 198754 212639 198782 213051
rect 198740 212630 198796 212639
rect 198740 212565 198796 212574
rect 197302 198753 197354 198759
rect 197302 198695 197354 198701
rect 197206 95005 197258 95011
rect 197206 94947 197258 94953
rect 197314 83541 197342 198695
rect 197398 135483 197450 135489
rect 197398 135425 197450 135431
rect 197302 83535 197354 83541
rect 197302 83477 197354 83483
rect 197410 71997 197438 135425
rect 198742 95005 198794 95011
rect 198742 94947 198794 94953
rect 198754 92463 198782 94947
rect 198934 94931 198986 94937
rect 198934 94873 198986 94879
rect 198836 93490 198892 93499
rect 198836 93425 198892 93434
rect 198740 92454 198796 92463
rect 198740 92389 198796 92398
rect 198850 92199 198878 93425
rect 198946 93351 198974 94873
rect 198932 93342 198988 93351
rect 198932 93277 198988 93286
rect 198838 92193 198890 92199
rect 198838 92135 198890 92141
rect 198742 92119 198794 92125
rect 198742 92061 198794 92067
rect 198754 91871 198782 92061
rect 199030 92045 199082 92051
rect 199030 91987 199082 91993
rect 198838 91897 198890 91903
rect 198740 91862 198796 91871
rect 198838 91839 198890 91845
rect 198740 91797 198796 91806
rect 198850 91131 198878 91839
rect 198934 91823 198986 91829
rect 198934 91765 198986 91771
rect 198836 91122 198892 91131
rect 198836 91057 198892 91066
rect 198946 90095 198974 91765
rect 199042 90243 199070 91987
rect 199126 91971 199178 91977
rect 199126 91913 199178 91919
rect 199138 91723 199166 91913
rect 199124 91714 199180 91723
rect 199124 91649 199180 91658
rect 199028 90234 199084 90243
rect 199028 90169 199084 90178
rect 198932 90086 198988 90095
rect 198932 90021 198988 90030
rect 198934 89233 198986 89239
rect 198934 89175 198986 89181
rect 198838 89085 198890 89091
rect 198740 89050 198796 89059
rect 198838 89027 198890 89033
rect 198740 88985 198742 88994
rect 198794 88985 198796 88994
rect 198742 88953 198794 88959
rect 198850 87875 198878 89027
rect 198946 88615 198974 89175
rect 199030 89159 199082 89165
rect 199030 89101 199082 89107
rect 198932 88606 198988 88615
rect 198932 88541 198988 88550
rect 198836 87866 198892 87875
rect 198836 87801 198892 87810
rect 199042 86987 199070 89101
rect 199222 88937 199274 88943
rect 199222 88879 199274 88885
rect 199234 88467 199262 88879
rect 199220 88458 199276 88467
rect 199220 88393 199276 88402
rect 199028 86978 199084 86987
rect 199028 86913 199084 86922
rect 199222 86421 199274 86427
rect 199222 86363 199274 86369
rect 199126 86347 199178 86353
rect 199126 86289 199178 86295
rect 198934 86273 198986 86279
rect 198836 86238 198892 86247
rect 198934 86215 198986 86221
rect 198836 86173 198892 86182
rect 198742 86125 198794 86131
rect 198740 86090 198742 86099
rect 198794 86090 198796 86099
rect 198850 86057 198878 86173
rect 198740 86025 198796 86034
rect 198838 86051 198890 86057
rect 198838 85993 198890 85999
rect 198946 85359 198974 86215
rect 199030 86199 199082 86205
rect 199030 86141 199082 86147
rect 198932 85350 198988 85359
rect 198932 85285 198988 85294
rect 199042 84619 199070 86141
rect 199138 85063 199166 86289
rect 199124 85054 199180 85063
rect 199124 84989 199180 84998
rect 199028 84610 199084 84619
rect 199028 84545 199084 84554
rect 199234 83731 199262 86363
rect 199220 83722 199276 83731
rect 199220 83657 199276 83666
rect 199510 83461 199562 83467
rect 199510 83403 199562 83409
rect 198838 83387 198890 83393
rect 198838 83329 198890 83335
rect 198740 83278 198796 83287
rect 198740 83213 198742 83222
rect 198794 83213 198796 83222
rect 198742 83181 198794 83187
rect 198850 81807 198878 83329
rect 198934 83313 198986 83319
rect 198934 83255 198986 83261
rect 198836 81798 198892 81807
rect 198836 81733 198892 81742
rect 198946 81363 198974 83255
rect 199522 82103 199550 83403
rect 199508 82094 199564 82103
rect 199508 82029 199564 82038
rect 198932 81354 198988 81363
rect 198932 81289 198988 81298
rect 198934 80649 198986 80655
rect 198934 80591 198986 80597
rect 198838 80501 198890 80507
rect 198740 80466 198796 80475
rect 198838 80443 198890 80449
rect 198740 80401 198742 80410
rect 198794 80401 198796 80410
rect 198742 80369 198794 80375
rect 198742 80279 198794 80285
rect 198742 80221 198794 80227
rect 198754 79883 198782 80221
rect 198740 79874 198796 79883
rect 198740 79809 198796 79818
rect 198850 79735 198878 80443
rect 198836 79726 198892 79735
rect 198836 79661 198892 79670
rect 198946 78847 198974 80591
rect 199030 80575 199082 80581
rect 199030 80517 199082 80523
rect 198932 78838 198988 78847
rect 198932 78773 198988 78782
rect 199042 78255 199070 80517
rect 199028 78246 199084 78255
rect 199028 78181 199084 78190
rect 199126 77763 199178 77769
rect 199126 77705 199178 77711
rect 198742 77689 198794 77695
rect 198740 77654 198742 77663
rect 198794 77654 198796 77663
rect 198740 77589 198796 77598
rect 198934 77615 198986 77621
rect 198934 77557 198986 77563
rect 198838 77467 198890 77473
rect 198838 77409 198890 77415
rect 198742 77393 198794 77399
rect 198742 77335 198794 77341
rect 198754 77219 198782 77335
rect 198740 77210 198796 77219
rect 198740 77145 198796 77154
rect 198850 76479 198878 77409
rect 198946 76627 198974 77557
rect 199030 77541 199082 77547
rect 199030 77483 199082 77489
rect 198932 76618 198988 76627
rect 198932 76553 198988 76562
rect 198836 76470 198892 76479
rect 198836 76405 198892 76414
rect 199042 75591 199070 77483
rect 199028 75582 199084 75591
rect 199028 75517 199084 75526
rect 199138 74999 199166 77705
rect 199124 74990 199180 74999
rect 199124 74925 199180 74934
rect 198934 74877 198986 74883
rect 198934 74819 198986 74825
rect 198742 74655 198794 74661
rect 198742 74597 198794 74603
rect 198754 74555 198782 74597
rect 198838 74581 198890 74587
rect 198740 74546 198796 74555
rect 198838 74523 198890 74529
rect 198740 74481 198796 74490
rect 198850 73371 198878 74523
rect 198946 73963 198974 74819
rect 199126 74803 199178 74809
rect 199126 74745 199178 74751
rect 199030 74729 199082 74735
rect 199030 74671 199082 74677
rect 198932 73954 198988 73963
rect 198932 73889 198988 73898
rect 198836 73362 198892 73371
rect 198836 73297 198892 73306
rect 199042 73223 199070 74671
rect 199028 73214 199084 73223
rect 199028 73149 199084 73158
rect 199138 72335 199166 74745
rect 199124 72326 199180 72335
rect 199124 72261 199180 72270
rect 197398 71991 197450 71997
rect 197398 71933 197450 71939
rect 194518 71917 194570 71923
rect 194518 71859 194570 71865
rect 199606 71917 199658 71923
rect 199606 71859 199658 71865
rect 191638 71843 191690 71849
rect 191638 71785 191690 71791
rect 198838 71843 198890 71849
rect 198838 71785 198890 71791
rect 188758 71769 188810 71775
rect 188758 71711 188810 71717
rect 198740 71734 198796 71743
rect 198740 71669 198742 71678
rect 198794 71669 198796 71678
rect 198742 71637 198794 71643
rect 198850 70115 198878 71785
rect 198934 71769 198986 71775
rect 198934 71711 198986 71717
rect 198836 70106 198892 70115
rect 198836 70041 198892 70050
rect 198946 69967 198974 71711
rect 199618 71003 199646 71859
rect 199604 70994 199660 71003
rect 199604 70929 199660 70938
rect 198932 69958 198988 69967
rect 198932 69893 198988 69902
rect 199030 69105 199082 69111
rect 199030 69047 199082 69053
rect 198934 68957 198986 68963
rect 198836 68922 198892 68931
rect 185878 68883 185930 68889
rect 198934 68899 198986 68905
rect 198836 68857 198838 68866
rect 185878 68825 185930 68831
rect 198890 68857 198892 68866
rect 198838 68825 198890 68831
rect 182998 68809 183050 68815
rect 182998 68751 183050 68757
rect 198742 68809 198794 68815
rect 198742 68751 198794 68757
rect 198754 68339 198782 68751
rect 198740 68330 198796 68339
rect 198740 68265 198796 68274
rect 198946 67747 198974 68899
rect 199042 68487 199070 69047
rect 199126 69031 199178 69037
rect 199126 68973 199178 68979
rect 199028 68478 199084 68487
rect 199028 68413 199084 68422
rect 198932 67738 198988 67747
rect 198932 67673 198988 67682
rect 199138 66859 199166 68973
rect 199124 66850 199180 66859
rect 199124 66785 199180 66794
rect 199126 66219 199178 66225
rect 199126 66161 199178 66167
rect 198932 66110 198988 66119
rect 198932 66045 198988 66054
rect 199030 66071 199082 66077
rect 198838 65997 198890 66003
rect 198740 65962 198796 65971
rect 198838 65939 198890 65945
rect 198740 65897 198742 65906
rect 198794 65897 198796 65906
rect 198742 65865 198794 65871
rect 177238 65849 177290 65855
rect 177238 65791 177290 65797
rect 198850 65231 198878 65939
rect 198946 65855 198974 66045
rect 199030 66013 199082 66019
rect 198934 65849 198986 65855
rect 198934 65791 198986 65797
rect 198836 65222 198892 65231
rect 198836 65157 198892 65166
rect 199042 64935 199070 66013
rect 199028 64926 199084 64935
rect 199028 64861 199084 64870
rect 199138 64491 199166 66161
rect 199222 66145 199274 66151
rect 199222 66087 199274 66093
rect 199124 64482 199180 64491
rect 199124 64417 199180 64426
rect 199234 63603 199262 66087
rect 199220 63594 199276 63603
rect 199220 63529 199276 63538
rect 199126 63333 199178 63339
rect 199126 63275 199178 63281
rect 199030 63259 199082 63265
rect 199030 63201 199082 63207
rect 198934 63185 198986 63191
rect 198740 63150 198796 63159
rect 198934 63127 198986 63133
rect 198740 63085 198796 63094
rect 198838 63111 198890 63117
rect 198754 63043 198782 63085
rect 198838 63053 198890 63059
rect 198742 63037 198794 63043
rect 198742 62979 198794 62985
rect 198850 62863 198878 63053
rect 198836 62854 198892 62863
rect 198836 62789 198892 62798
rect 198946 61975 198974 63127
rect 198932 61966 198988 61975
rect 198932 61901 198988 61910
rect 199042 61679 199070 63201
rect 199028 61670 199084 61679
rect 199028 61605 199084 61614
rect 199138 61235 199166 63275
rect 199124 61226 199180 61235
rect 199124 61161 199180 61170
rect 198934 60447 198986 60453
rect 198934 60389 198986 60395
rect 198838 60373 198890 60379
rect 198740 60338 198796 60347
rect 167062 60299 167114 60305
rect 198838 60315 198890 60321
rect 198740 60273 198742 60282
rect 167062 60241 167114 60247
rect 198794 60273 198796 60282
rect 198742 60241 198794 60247
rect 198850 59755 198878 60315
rect 198836 59746 198892 59755
rect 198836 59681 198892 59690
rect 198946 59607 198974 60389
rect 198932 59598 198988 59607
rect 198932 59533 198988 59542
rect 199714 53867 199742 221741
rect 199702 53861 199754 53867
rect 199702 53803 199754 53809
rect 199810 53571 199838 222037
rect 200098 221847 200126 227481
rect 199990 221841 200042 221847
rect 199990 221783 200042 221789
rect 200086 221841 200138 221847
rect 200086 221783 200138 221789
rect 200002 218610 200030 221783
rect 200194 221371 200222 252567
rect 200290 222111 200318 254861
rect 200374 252699 200426 252705
rect 200374 252641 200426 252647
rect 200276 222102 200332 222111
rect 200276 222037 200332 222046
rect 200180 221362 200236 221371
rect 200180 221297 200236 221306
rect 200386 220779 200414 252641
rect 200566 252551 200618 252557
rect 200566 252493 200618 252499
rect 200470 252477 200522 252483
rect 200470 252419 200522 252425
rect 200482 221815 200510 252419
rect 200468 221806 200524 221815
rect 200468 221741 200524 221750
rect 200372 220770 200428 220779
rect 200372 220705 200428 220714
rect 200578 219891 200606 252493
rect 204214 252033 204266 252039
rect 204214 251975 204266 251981
rect 200758 247593 200810 247599
rect 200758 247535 200810 247541
rect 200564 219882 200620 219891
rect 200564 219817 200620 219826
rect 200770 219743 200798 247535
rect 204226 241975 204254 251975
rect 204214 241969 204266 241975
rect 204214 241911 204266 241917
rect 204322 236055 204350 268995
rect 204994 267431 205022 275502
rect 204982 267425 205034 267431
rect 204982 267367 205034 267373
rect 206146 261585 206174 275502
rect 207284 273458 207340 273467
rect 207284 273393 207286 273402
rect 207338 273393 207340 273402
rect 207286 273361 207338 273367
rect 207394 263953 207422 275502
rect 208438 273419 208490 273425
rect 208438 273361 208490 273367
rect 208450 273319 208478 273361
rect 208436 273310 208492 273319
rect 208436 273245 208492 273254
rect 208546 267505 208574 275502
rect 209808 275488 210014 275516
rect 208534 267499 208586 267505
rect 208534 267441 208586 267447
rect 207382 263947 207434 263953
rect 207382 263889 207434 263895
rect 206134 261579 206186 261585
rect 206134 261521 206186 261527
rect 204406 253587 204458 253593
rect 204406 253529 204458 253535
rect 204310 236049 204362 236055
rect 204310 235991 204362 235997
rect 202580 228762 202636 228771
rect 202580 228697 202636 228706
rect 202594 227735 202622 228697
rect 202580 227726 202636 227735
rect 202580 227661 202636 227670
rect 204310 223839 204362 223845
rect 204310 223781 204362 223787
rect 201236 221362 201292 221371
rect 201236 221297 201292 221306
rect 201140 219882 201196 219891
rect 201140 219817 201196 219826
rect 200756 219734 200812 219743
rect 200756 219669 200812 219678
rect 200002 218582 200414 218610
rect 200386 202871 200414 218582
rect 200372 202862 200428 202871
rect 200372 202797 200428 202806
rect 200662 201565 200714 201571
rect 200662 201507 200714 201513
rect 200674 181517 200702 201507
rect 200770 187289 200798 219669
rect 200948 202862 201004 202871
rect 200948 202797 201004 202806
rect 200962 201571 200990 202797
rect 200950 201565 201002 201571
rect 200950 201507 201002 201513
rect 200758 187283 200810 187289
rect 200758 187225 200810 187231
rect 201046 187283 201098 187289
rect 201046 187225 201098 187231
rect 200662 181511 200714 181517
rect 200662 181453 200714 181459
rect 200854 181511 200906 181517
rect 200854 181453 200906 181459
rect 200866 181411 200894 181453
rect 200852 181402 200908 181411
rect 200852 181337 200908 181346
rect 200948 166898 201004 166907
rect 200948 166833 201004 166842
rect 200962 126799 200990 166833
rect 200756 126790 200812 126799
rect 200756 126725 200812 126734
rect 200948 126790 201004 126799
rect 200948 126725 201004 126734
rect 200770 120985 200798 126725
rect 201058 126683 201086 187225
rect 200854 126677 200906 126683
rect 200854 126619 200906 126625
rect 201046 126677 201098 126683
rect 201046 126619 201098 126625
rect 200866 120985 200894 126619
rect 200470 120979 200522 120985
rect 200470 120921 200522 120927
rect 200758 120979 200810 120985
rect 200758 120921 200810 120927
rect 200854 120979 200906 120985
rect 200854 120921 200906 120927
rect 201046 120979 201098 120985
rect 201046 120921 201098 120927
rect 200482 106555 200510 120921
rect 200470 106549 200522 106555
rect 200470 106491 200522 106497
rect 200662 106549 200714 106555
rect 200662 106491 200714 106497
rect 200674 54089 200702 106491
rect 201058 86427 201086 120921
rect 200854 86421 200906 86427
rect 200854 86363 200906 86369
rect 201046 86421 201098 86427
rect 201046 86363 201098 86369
rect 200758 83535 200810 83541
rect 200758 83477 200810 83483
rect 200770 82991 200798 83477
rect 200756 82982 200812 82991
rect 200756 82917 200812 82926
rect 200758 71991 200810 71997
rect 200758 71933 200810 71939
rect 200770 71595 200798 71933
rect 200756 71586 200812 71595
rect 200756 71521 200812 71530
rect 200866 66373 200894 86363
rect 200854 66367 200906 66373
rect 200854 66309 200906 66315
rect 201046 66293 201098 66299
rect 201046 66235 201098 66241
rect 201058 54163 201086 66235
rect 201046 54157 201098 54163
rect 201046 54099 201098 54105
rect 200662 54083 200714 54089
rect 200662 54025 200714 54031
rect 201154 54015 201182 219817
rect 201142 54009 201194 54015
rect 201142 53951 201194 53957
rect 201250 53719 201278 221297
rect 201332 220770 201388 220779
rect 201332 220705 201388 220714
rect 201346 60028 201374 220705
rect 202966 152725 203018 152731
rect 202966 152667 203018 152673
rect 202774 103811 202826 103817
rect 202774 103753 202826 103759
rect 202678 100851 202730 100857
rect 202678 100793 202730 100799
rect 202582 97965 202634 97971
rect 202582 97907 202634 97913
rect 202198 95153 202250 95159
rect 202198 95095 202250 95101
rect 201814 95079 201866 95085
rect 201814 95021 201866 95027
rect 201826 80729 201854 95021
rect 202210 86353 202238 95095
rect 202594 86575 202622 97907
rect 202582 86569 202634 86575
rect 202582 86511 202634 86517
rect 202390 86495 202442 86501
rect 202390 86437 202442 86443
rect 202198 86347 202250 86353
rect 202198 86289 202250 86295
rect 201814 80723 201866 80729
rect 201814 80665 201866 80671
rect 202102 80723 202154 80729
rect 202102 80665 202154 80671
rect 202006 61557 202058 61563
rect 202006 61499 202058 61505
rect 201346 60000 201470 60028
rect 201332 55602 201388 55611
rect 201332 55537 201388 55546
rect 201238 53713 201290 53719
rect 201238 53655 201290 53661
rect 199798 53565 199850 53571
rect 199798 53507 199850 53513
rect 163510 53491 163562 53497
rect 163510 53433 163562 53439
rect 163414 52973 163466 52979
rect 163414 52915 163466 52921
rect 163318 52825 163370 52831
rect 163318 52767 163370 52773
rect 163222 52381 163274 52387
rect 163222 52323 163274 52329
rect 163126 52233 163178 52239
rect 163126 52175 163178 52181
rect 162742 52159 162794 52165
rect 162742 52101 162794 52107
rect 159958 52011 160010 52017
rect 159958 51953 160010 51959
rect 149686 46757 149738 46763
rect 149686 46699 149738 46705
rect 161300 46722 161356 46731
rect 149302 46683 149354 46689
rect 161300 46657 161302 46666
rect 149302 46625 149354 46631
rect 161354 46657 161356 46666
rect 181364 46722 181420 46731
rect 181364 46657 181366 46666
rect 161302 46625 161354 46631
rect 181418 46657 181420 46666
rect 181366 46625 181418 46631
rect 147958 46387 148010 46393
rect 147958 46329 148010 46335
rect 147766 46239 147818 46245
rect 147766 46181 147818 46187
rect 201346 42175 201374 55537
rect 201442 53793 201470 60000
rect 201430 53787 201482 53793
rect 201430 53729 201482 53735
rect 201622 48237 201674 48243
rect 201622 48179 201674 48185
rect 201634 47503 201662 48179
rect 201622 47497 201674 47503
rect 201622 47439 201674 47445
rect 202018 46319 202046 61499
rect 202114 53423 202142 80665
rect 202294 61483 202346 61489
rect 202294 61425 202346 61431
rect 202198 61409 202250 61415
rect 202198 61351 202250 61357
rect 202102 53417 202154 53423
rect 202102 53359 202154 53365
rect 202006 46313 202058 46319
rect 202006 46255 202058 46261
rect 202210 46171 202238 61351
rect 202306 46467 202334 61425
rect 202402 48095 202430 86437
rect 202582 86347 202634 86353
rect 202582 86289 202634 86295
rect 202486 61335 202538 61341
rect 202486 61277 202538 61283
rect 202390 48089 202442 48095
rect 202390 48031 202442 48037
rect 202498 46615 202526 61277
rect 202594 48983 202622 86289
rect 202582 48977 202634 48983
rect 202582 48919 202634 48925
rect 202690 48909 202718 100793
rect 202678 48903 202730 48909
rect 202678 48845 202730 48851
rect 202786 48835 202814 103753
rect 202870 103737 202922 103743
rect 202870 103679 202922 103685
rect 202882 53391 202910 103679
rect 202978 61489 203006 152667
rect 203062 149839 203114 149845
rect 203062 149781 203114 149787
rect 203074 61563 203102 149781
rect 203158 141181 203210 141187
rect 203158 141123 203210 141129
rect 203062 61557 203114 61563
rect 203062 61499 203114 61505
rect 202966 61483 203018 61489
rect 202966 61425 203018 61431
rect 203170 61360 203198 141123
rect 203254 138295 203306 138301
rect 203254 138237 203306 138243
rect 202978 61332 203198 61360
rect 203266 61341 203294 138237
rect 203350 135409 203402 135415
rect 203350 135351 203402 135357
rect 203362 61415 203390 135351
rect 203446 129637 203498 129643
rect 203446 129579 203498 129585
rect 203350 61409 203402 61415
rect 203350 61351 203402 61357
rect 203254 61335 203306 61341
rect 202868 53382 202924 53391
rect 202868 53317 202924 53326
rect 202978 51573 203006 61332
rect 203254 61277 203306 61283
rect 203458 61212 203486 129579
rect 203542 126751 203594 126757
rect 203542 126693 203594 126699
rect 203074 61184 203486 61212
rect 203074 52799 203102 61184
rect 203554 61064 203582 126693
rect 203734 124013 203786 124019
rect 203734 123955 203786 123961
rect 203638 123939 203690 123945
rect 203638 123881 203690 123887
rect 203170 61036 203582 61064
rect 203060 52790 203116 52799
rect 203060 52725 203116 52734
rect 203170 52651 203198 61036
rect 203254 60891 203306 60897
rect 203650 60842 203678 123881
rect 203746 60897 203774 123955
rect 203830 121053 203882 121059
rect 203830 120995 203882 121001
rect 203254 60833 203306 60839
rect 203156 52642 203212 52651
rect 203156 52577 203212 52586
rect 202966 51567 203018 51573
rect 202966 51509 203018 51515
rect 202774 48829 202826 48835
rect 202774 48771 202826 48777
rect 203266 47873 203294 60833
rect 203362 60814 203678 60842
rect 203734 60891 203786 60897
rect 203734 60833 203786 60839
rect 203362 47947 203390 60814
rect 203842 60768 203870 120995
rect 203926 118167 203978 118173
rect 203926 118109 203978 118115
rect 203458 60740 203870 60768
rect 203458 48243 203486 60740
rect 203938 60620 203966 118109
rect 204022 115281 204074 115287
rect 204022 115223 204074 115229
rect 204034 62271 204062 115223
rect 204118 112469 204170 112475
rect 204118 112411 204170 112417
rect 204020 62262 204076 62271
rect 204020 62197 204076 62206
rect 203554 60592 203966 60620
rect 203554 53539 203582 60592
rect 204130 60324 204158 112411
rect 204214 109509 204266 109515
rect 204214 109451 204266 109457
rect 203746 60296 204158 60324
rect 203540 53530 203596 53539
rect 203540 53465 203596 53474
rect 203746 48465 203774 60296
rect 204226 60176 204254 109451
rect 203842 60148 204254 60176
rect 203842 48539 203870 60148
rect 204322 60028 204350 223781
rect 203938 60000 204350 60028
rect 203938 52947 203966 60000
rect 204418 59880 204446 253529
rect 204502 252403 204554 252409
rect 204502 252345 204554 252351
rect 204514 230103 204542 252345
rect 204694 252329 204746 252335
rect 204694 252271 204746 252277
rect 204598 252107 204650 252113
rect 204598 252049 204650 252055
rect 204500 230094 204556 230103
rect 204500 230029 204556 230038
rect 204610 228729 204638 252049
rect 204598 228723 204650 228729
rect 204598 228665 204650 228671
rect 204706 228600 204734 252271
rect 204886 252255 204938 252261
rect 204886 252197 204938 252203
rect 204790 252181 204842 252187
rect 204790 252123 204842 252129
rect 204514 228572 204734 228600
rect 204514 227767 204542 228572
rect 204694 228353 204746 228359
rect 204694 228295 204746 228301
rect 204502 227761 204554 227767
rect 204502 227703 204554 227709
rect 204514 223253 204542 227703
rect 204502 223247 204554 223253
rect 204502 223189 204554 223195
rect 204502 223099 204554 223105
rect 204502 223041 204554 223047
rect 204322 59852 204446 59880
rect 204022 59115 204074 59121
rect 204022 59057 204074 59063
rect 203924 52938 203980 52947
rect 203924 52873 203980 52882
rect 204034 51592 204062 59057
rect 204118 57339 204170 57345
rect 204118 57281 204170 57287
rect 204130 53275 204158 57281
rect 204214 56303 204266 56309
rect 204214 56245 204266 56251
rect 204118 53269 204170 53275
rect 204118 53211 204170 53217
rect 204226 52924 204254 56245
rect 204322 53645 204350 59852
rect 204404 58118 204460 58127
rect 204404 58053 204460 58062
rect 204310 53639 204362 53645
rect 204310 53581 204362 53587
rect 204310 53417 204362 53423
rect 204310 53359 204362 53365
rect 204322 53095 204350 53359
rect 204418 53127 204446 58053
rect 204514 57345 204542 223041
rect 204598 207411 204650 207417
rect 204598 207353 204650 207359
rect 204610 58696 204638 207353
rect 204706 58867 204734 228295
rect 204802 227619 204830 252123
rect 204898 230524 204926 252197
rect 207382 241969 207434 241975
rect 207382 241911 207434 241917
rect 204898 230496 205118 230524
rect 204884 230390 204940 230399
rect 204884 230325 204940 230334
rect 204790 227613 204842 227619
rect 204790 227555 204842 227561
rect 204802 58973 204830 227555
rect 204898 222976 204926 230325
rect 204980 230094 205036 230103
rect 204980 230029 205036 230038
rect 204994 227693 205022 230029
rect 205090 228359 205118 230496
rect 205460 230242 205516 230251
rect 205460 230177 205516 230186
rect 205078 228353 205130 228359
rect 205078 228295 205130 228301
rect 204982 227687 205034 227693
rect 204982 227629 205034 227635
rect 204994 223105 205022 227629
rect 205474 224035 205502 230177
rect 205846 228723 205898 228729
rect 205846 228665 205898 228671
rect 205460 224026 205516 224035
rect 205460 223961 205516 223970
rect 205474 223554 205502 223961
rect 205858 223887 205886 228665
rect 206614 228353 206666 228359
rect 206614 228295 206666 228301
rect 206230 227613 206282 227619
rect 206230 227555 206282 227561
rect 205844 223878 205900 223887
rect 205844 223813 205900 223822
rect 205858 223554 205886 223813
rect 206242 223554 206270 227555
rect 206626 223554 206654 228295
rect 206902 227761 206954 227767
rect 206902 227703 206954 227709
rect 206914 223864 206942 227703
rect 207286 227687 207338 227693
rect 207286 227629 207338 227635
rect 207298 223864 207326 227629
rect 207394 223993 207422 241911
rect 209986 235981 210014 275488
rect 210946 268837 210974 275502
rect 212194 268911 212222 275502
rect 212182 268905 212234 268911
rect 212182 268847 212234 268853
rect 212950 268905 213002 268911
rect 212950 268847 213002 268853
rect 210934 268831 210986 268837
rect 210934 268773 210986 268779
rect 212962 238835 212990 268847
rect 213046 268831 213098 268837
rect 213046 268773 213098 268779
rect 212948 238826 213004 238835
rect 212948 238761 213004 238770
rect 209974 235975 210026 235981
rect 209974 235917 210026 235923
rect 213058 234987 213086 268773
rect 213346 260327 213374 275502
rect 214498 264175 214526 275502
rect 215746 267579 215774 275502
rect 215734 267573 215786 267579
rect 215734 267515 215786 267521
rect 214486 264169 214538 264175
rect 214486 264111 214538 264117
rect 216802 260401 216830 275502
rect 218050 260623 218078 275502
rect 219202 268911 219230 275502
rect 219190 268905 219242 268911
rect 219190 268847 219242 268853
rect 218038 260617 218090 260623
rect 218038 260559 218090 260565
rect 218710 260617 218762 260623
rect 218806 260617 218858 260623
rect 218710 260559 218762 260565
rect 218804 260582 218806 260591
rect 218858 260582 218860 260591
rect 216790 260395 216842 260401
rect 216790 260337 216842 260343
rect 213334 260321 213386 260327
rect 213334 260263 213386 260269
rect 218722 255832 218750 260559
rect 218804 260517 218860 260526
rect 220450 260401 220478 275502
rect 221494 268905 221546 268911
rect 221494 268847 221546 268853
rect 218806 260395 218858 260401
rect 218806 260337 218858 260343
rect 220438 260395 220490 260401
rect 220438 260337 220490 260343
rect 218422 255807 218474 255813
rect 218422 255749 218474 255755
rect 218626 255804 218750 255832
rect 218818 255813 218846 260337
rect 218806 255807 218858 255813
rect 218434 249153 218462 255749
rect 218626 249172 218654 255804
rect 218806 255749 218858 255755
rect 218902 255733 218954 255739
rect 218902 255675 218954 255681
rect 218914 255517 218942 255675
rect 218902 255511 218954 255517
rect 218902 255453 218954 255459
rect 218422 249147 218474 249153
rect 218626 249144 218750 249172
rect 218422 249089 218474 249095
rect 218722 239015 218750 249144
rect 218806 249147 218858 249153
rect 218806 249089 218858 249095
rect 218710 239009 218762 239015
rect 218710 238951 218762 238957
rect 218818 236129 218846 249089
rect 221506 238539 221534 268847
rect 221602 266913 221630 275502
rect 222850 268837 222878 275502
rect 224016 275488 224606 275516
rect 222838 268831 222890 268837
rect 222838 268773 222890 268779
rect 221590 266907 221642 266913
rect 221590 266849 221642 266855
rect 221686 262985 221738 262991
rect 221782 262985 221834 262991
rect 221738 262933 221782 262936
rect 221686 262927 221834 262933
rect 221698 262908 221822 262927
rect 221492 238530 221548 238539
rect 221492 238465 221548 238474
rect 218806 236123 218858 236129
rect 218806 236065 218858 236071
rect 224578 235759 224606 275488
rect 225250 268911 225278 275502
rect 225238 268905 225290 268911
rect 225238 268847 225290 268853
rect 226402 268689 226430 275502
rect 227350 268905 227402 268911
rect 227350 268847 227402 268853
rect 226390 268683 226442 268689
rect 226390 268625 226442 268631
rect 227362 238941 227390 268847
rect 227650 268837 227678 275502
rect 227638 268831 227690 268837
rect 227638 268773 227690 268779
rect 227446 268683 227498 268689
rect 227446 268625 227498 268631
rect 227350 238935 227402 238941
rect 227350 238877 227402 238883
rect 227458 238391 227486 268625
rect 228802 263731 228830 275502
rect 229954 266765 229982 275502
rect 230134 268831 230186 268837
rect 230134 268773 230186 268779
rect 229942 266759 229994 266765
rect 229942 266701 229994 266707
rect 228790 263725 228842 263731
rect 228790 263667 228842 263673
rect 230146 250559 230174 268773
rect 231202 261955 231230 275502
rect 232354 263657 232382 275502
rect 233506 266839 233534 275502
rect 234658 268837 234686 275502
rect 235920 275488 236030 275516
rect 234646 268831 234698 268837
rect 234646 268773 234698 268779
rect 235894 268831 235946 268837
rect 235894 268773 235946 268779
rect 233494 266833 233546 266839
rect 233494 266775 233546 266781
rect 232342 263651 232394 263657
rect 232342 263593 232394 263599
rect 231190 261949 231242 261955
rect 231190 261891 231242 261897
rect 234070 261875 234122 261881
rect 234070 261817 234122 261823
rect 233206 261801 233258 261807
rect 233206 261743 233258 261749
rect 233218 258477 233246 261743
rect 234082 258551 234110 261817
rect 234070 258545 234122 258551
rect 234070 258487 234122 258493
rect 233206 258471 233258 258477
rect 233206 258413 233258 258419
rect 230134 250553 230186 250559
rect 230134 250495 230186 250501
rect 235906 247673 235934 268773
rect 236002 266987 236030 275488
rect 235990 266981 236042 266987
rect 235990 266923 236042 266929
rect 237058 263255 237086 275502
rect 237044 263246 237100 263255
rect 236194 263204 236318 263232
rect 236194 263139 236222 263204
rect 236182 263133 236234 263139
rect 236182 263075 236234 263081
rect 236290 263065 236318 263204
rect 237044 263181 237100 263190
rect 236278 263059 236330 263065
rect 236278 263001 236330 263007
rect 238306 261881 238334 275502
rect 239458 263805 239486 275502
rect 240706 267653 240734 275502
rect 241666 275488 241872 275516
rect 240694 267647 240746 267653
rect 240694 267589 240746 267595
rect 239446 263799 239498 263805
rect 239446 263741 239498 263747
rect 238294 261875 238346 261881
rect 238294 261817 238346 261823
rect 235894 247667 235946 247673
rect 235894 247609 235946 247615
rect 241666 244787 241694 275488
rect 243106 264249 243134 275502
rect 244258 267727 244286 275502
rect 244246 267721 244298 267727
rect 244246 267663 244298 267669
rect 243094 264243 243146 264249
rect 243094 264185 243146 264191
rect 245410 261955 245438 275502
rect 246658 264323 246686 275502
rect 247810 267801 247838 275502
rect 247892 273606 247948 273615
rect 247892 273541 247948 273550
rect 247906 273319 247934 273541
rect 247892 273310 247948 273319
rect 247892 273245 247948 273254
rect 247798 267795 247850 267801
rect 247798 267737 247850 267743
rect 246646 264317 246698 264323
rect 246646 264259 246698 264265
rect 249058 262029 249086 275502
rect 250114 264397 250142 275502
rect 251362 264989 251390 275502
rect 252514 268837 252542 275502
rect 252502 268831 252554 268837
rect 252502 268773 252554 268779
rect 253366 268831 253418 268837
rect 253366 268773 253418 268779
rect 251350 264983 251402 264989
rect 251350 264925 251402 264931
rect 250102 264391 250154 264397
rect 250102 264333 250154 264339
rect 249046 262023 249098 262029
rect 249046 261965 249098 261971
rect 245398 261949 245450 261955
rect 245398 261891 245450 261897
rect 241654 244781 241706 244787
rect 241654 244723 241706 244729
rect 253378 244713 253406 268773
rect 253762 264545 253790 275502
rect 254914 266321 254942 275502
rect 254902 266315 254954 266321
rect 254902 266257 254954 266263
rect 253750 264539 253802 264545
rect 253750 264481 253802 264487
rect 256162 262103 256190 275502
rect 256342 273345 256394 273351
rect 256340 273310 256342 273319
rect 256394 273310 256396 273319
rect 256340 273245 256396 273254
rect 256918 267129 256970 267135
rect 256918 267071 256970 267077
rect 256930 266839 256958 267071
rect 256918 266833 256970 266839
rect 256918 266775 256970 266781
rect 257314 264693 257342 275502
rect 258562 266247 258590 275502
rect 259714 268837 259742 275502
rect 259702 268831 259754 268837
rect 259702 268773 259754 268779
rect 258550 266241 258602 266247
rect 258550 266183 258602 266189
rect 257302 264687 257354 264693
rect 257302 264629 257354 264635
rect 260866 264619 260894 275502
rect 262006 268831 262058 268837
rect 262006 268773 262058 268779
rect 260854 264613 260906 264619
rect 260854 264555 260906 264561
rect 256150 262097 256202 262103
rect 256150 262039 256202 262045
rect 259318 255955 259370 255961
rect 259318 255897 259370 255903
rect 259330 255684 259358 255897
rect 259234 255665 259358 255684
rect 259222 255659 259358 255665
rect 259274 255656 259358 255659
rect 259222 255601 259274 255607
rect 253366 244707 253418 244713
rect 253366 244649 253418 244655
rect 262018 244639 262046 268773
rect 262114 266173 262142 275502
rect 262102 266167 262154 266173
rect 262102 266109 262154 266115
rect 262102 263133 262154 263139
rect 262294 263133 262346 263139
rect 262154 263081 262294 263084
rect 262102 263075 262346 263081
rect 262114 263056 262334 263075
rect 263266 260623 263294 275502
rect 264514 264767 264542 275502
rect 265666 265877 265694 275502
rect 266818 268837 266846 275502
rect 266806 268831 266858 268837
rect 266806 268773 266858 268779
rect 267766 268831 267818 268837
rect 267766 268773 267818 268779
rect 265654 265871 265706 265877
rect 265654 265813 265706 265819
rect 264502 264761 264554 264767
rect 264502 264703 264554 264709
rect 263254 260617 263306 260623
rect 263254 260559 263306 260565
rect 262006 244633 262058 244639
rect 262006 244575 262058 244581
rect 267778 244565 267806 268773
rect 267970 264841 267998 275502
rect 267958 264835 268010 264841
rect 267958 264777 268010 264783
rect 269218 260253 269246 275502
rect 270370 260549 270398 275502
rect 271618 264915 271646 275502
rect 272770 266025 272798 275502
rect 274018 268837 274046 275502
rect 274006 268831 274058 268837
rect 274006 268773 274058 268779
rect 272758 266019 272810 266025
rect 272758 265961 272810 265967
rect 271606 264909 271658 264915
rect 271606 264851 271658 264857
rect 275170 263583 275198 275502
rect 276322 268689 276350 275502
rect 276404 273754 276460 273763
rect 276404 273689 276460 273698
rect 276418 273351 276446 273689
rect 276406 273345 276458 273351
rect 276406 273287 276458 273293
rect 276406 268831 276458 268837
rect 276406 268773 276458 268779
rect 276310 268683 276362 268689
rect 276310 268625 276362 268631
rect 275158 263577 275210 263583
rect 275158 263519 275210 263525
rect 270358 260543 270410 260549
rect 270358 260485 270410 260491
rect 269206 260247 269258 260253
rect 269206 260189 269258 260195
rect 267766 244559 267818 244565
rect 267766 244501 267818 244507
rect 276418 244491 276446 268773
rect 277078 261801 277130 261807
rect 277078 261743 277130 261749
rect 277090 254999 277118 261743
rect 277570 260475 277598 275502
rect 277846 267129 277898 267135
rect 277846 267071 277898 267077
rect 277858 266839 277886 267071
rect 277942 267055 277994 267061
rect 277942 266997 277994 267003
rect 277846 266833 277898 266839
rect 277846 266775 277898 266781
rect 277846 266611 277898 266617
rect 277846 266553 277898 266559
rect 277558 260469 277610 260475
rect 277558 260411 277610 260417
rect 277858 258699 277886 266553
rect 277846 258693 277898 258699
rect 277846 258635 277898 258641
rect 277954 258625 277982 266997
rect 278722 263361 278750 275502
rect 279970 265803 279998 275502
rect 281122 268319 281150 275502
rect 282384 275488 282974 275516
rect 282166 273789 282218 273795
rect 282164 273754 282166 273763
rect 282218 273754 282220 273763
rect 282164 273689 282220 273698
rect 281110 268313 281162 268319
rect 281110 268255 281162 268261
rect 282838 267055 282890 267061
rect 282838 266997 282890 267003
rect 282262 266685 282314 266691
rect 282262 266627 282314 266633
rect 279958 265797 280010 265803
rect 279958 265739 280010 265745
rect 278710 263355 278762 263361
rect 278710 263297 278762 263303
rect 279478 260987 279530 260993
rect 279478 260929 279530 260935
rect 279382 260691 279434 260697
rect 279382 260633 279434 260639
rect 279394 260605 279422 260633
rect 279490 260605 279518 260929
rect 279394 260577 279518 260605
rect 282274 258773 282302 266627
rect 282466 266460 282686 266488
rect 282466 259532 282494 266460
rect 282658 266395 282686 266460
rect 282550 266389 282602 266395
rect 282550 266331 282602 266337
rect 282646 266389 282698 266395
rect 282646 266331 282698 266337
rect 282370 259504 282494 259532
rect 282262 258767 282314 258773
rect 282262 258709 282314 258715
rect 277942 258619 277994 258625
rect 277942 258561 277994 258567
rect 282262 257731 282314 257737
rect 282262 257673 282314 257679
rect 277078 254993 277130 254999
rect 277078 254935 277130 254941
rect 282274 245028 282302 257673
rect 282370 248931 282398 259504
rect 282454 259359 282506 259365
rect 282454 259301 282506 259307
rect 282358 248925 282410 248931
rect 282358 248867 282410 248873
rect 282358 247667 282410 247673
rect 282358 247609 282410 247615
rect 282370 245347 282398 247609
rect 282356 245338 282412 245347
rect 282356 245273 282412 245282
rect 282274 245000 282398 245028
rect 282166 244855 282218 244861
rect 282166 244797 282218 244803
rect 276406 244485 276458 244491
rect 276406 244427 276458 244433
rect 282178 243548 282206 244797
rect 282262 244781 282314 244787
rect 282260 244746 282262 244755
rect 282314 244746 282316 244755
rect 282260 244681 282316 244690
rect 282262 244633 282314 244639
rect 282262 244575 282314 244581
rect 282274 243719 282302 244575
rect 282260 243710 282316 243719
rect 282260 243645 282316 243654
rect 282178 243520 282302 243548
rect 227444 238382 227500 238391
rect 227444 238317 227500 238326
rect 224566 235753 224618 235759
rect 224566 235695 224618 235701
rect 213044 234978 213100 234987
rect 213044 234913 213100 234922
rect 207862 230425 207914 230431
rect 207862 230367 207914 230373
rect 208052 230390 208108 230399
rect 207766 230351 207818 230357
rect 207766 230293 207818 230299
rect 207778 227767 207806 230293
rect 207766 227761 207818 227767
rect 207766 227703 207818 227709
rect 207778 226699 207806 227703
rect 207874 227693 207902 230367
rect 208052 230325 208108 230334
rect 208436 230390 208492 230399
rect 208436 230325 208492 230334
rect 207862 227687 207914 227693
rect 207862 227629 207914 227635
rect 207874 226847 207902 227629
rect 207860 226838 207916 226847
rect 207860 226773 207916 226782
rect 207764 226690 207820 226699
rect 207764 226625 207820 226634
rect 207382 223987 207434 223993
rect 207382 223929 207434 223935
rect 208066 223887 208094 230325
rect 208150 230277 208202 230283
rect 208150 230219 208202 230225
rect 208162 227545 208190 230219
rect 208150 227539 208202 227545
rect 208150 227481 208202 227487
rect 208162 226551 208190 227481
rect 208148 226542 208204 226551
rect 208148 226477 208204 226486
rect 208450 223887 208478 230325
rect 212470 230203 212522 230209
rect 212470 230145 212522 230151
rect 212086 230129 212138 230135
rect 212086 230071 212138 230077
rect 211702 230055 211754 230061
rect 211702 229997 211754 230003
rect 211030 229981 211082 229987
rect 211030 229923 211082 229929
rect 209494 229907 209546 229913
rect 209494 229849 209546 229855
rect 208822 229759 208874 229765
rect 208822 229701 208874 229707
rect 208052 223878 208108 223887
rect 206914 223836 206990 223864
rect 207298 223836 207374 223864
rect 206962 223554 206990 223836
rect 207346 223554 207374 223836
rect 207670 223839 207722 223845
rect 208052 223813 208108 223822
rect 208436 223878 208492 223887
rect 208436 223813 208492 223822
rect 207670 223781 207722 223787
rect 207682 223554 207710 223781
rect 208066 223554 208094 223813
rect 208450 223554 208478 223813
rect 208834 223554 208862 229701
rect 209110 229685 209162 229691
rect 209110 229627 209162 229633
rect 209122 223864 209150 229627
rect 209506 223864 209534 229849
rect 209878 229833 209930 229839
rect 209878 229775 209930 229781
rect 209122 223836 209198 223864
rect 209506 223836 209582 223864
rect 209170 223554 209198 223836
rect 209554 223554 209582 223836
rect 209890 223554 209918 229775
rect 210646 229611 210698 229617
rect 210646 229553 210698 229559
rect 210262 229537 210314 229543
rect 210262 229479 210314 229485
rect 210274 223554 210302 229479
rect 210658 223554 210686 229553
rect 211042 223554 211070 229923
rect 211318 229389 211370 229395
rect 211318 229331 211370 229337
rect 211330 223864 211358 229331
rect 211714 223864 211742 229997
rect 211330 223836 211406 223864
rect 211714 223836 211790 223864
rect 211378 223554 211406 223836
rect 211762 223554 211790 223836
rect 212098 223554 212126 230071
rect 212482 223554 212510 230145
rect 215062 229463 215114 229469
rect 215062 229405 215114 229411
rect 213910 229315 213962 229321
rect 213910 229257 213962 229263
rect 212854 228945 212906 228951
rect 212854 228887 212906 228893
rect 212866 223554 212894 228887
rect 213238 228871 213290 228877
rect 213238 228813 213290 228819
rect 213250 223554 213278 228813
rect 213526 228797 213578 228803
rect 213526 228739 213578 228745
rect 213538 223864 213566 228739
rect 213922 223864 213950 229257
rect 214678 229241 214730 229247
rect 214678 229183 214730 229189
rect 214294 228723 214346 228729
rect 214294 228665 214346 228671
rect 213538 223836 213614 223864
rect 213922 223836 213998 223864
rect 213586 223554 213614 223836
rect 213970 223554 213998 223836
rect 214306 223554 214334 228665
rect 214690 223554 214718 229183
rect 215074 223554 215102 229405
rect 215446 229167 215498 229173
rect 215446 229109 215498 229115
rect 215458 223554 215486 229109
rect 282274 229099 282302 243520
rect 282370 242387 282398 245000
rect 282466 244639 282494 259301
rect 282562 257631 282590 266331
rect 282742 265871 282794 265877
rect 282742 265813 282794 265819
rect 282548 257622 282604 257631
rect 282548 257557 282604 257566
rect 282550 256843 282602 256849
rect 282550 256785 282602 256791
rect 282454 244633 282506 244639
rect 282454 244575 282506 244581
rect 282454 244485 282506 244491
rect 282454 244427 282506 244433
rect 282466 242535 282494 244427
rect 282452 242526 282508 242535
rect 282452 242461 282508 242470
rect 282356 242378 282412 242387
rect 282356 242313 282412 242322
rect 282562 237831 282590 256785
rect 282646 256103 282698 256109
rect 282646 256045 282698 256051
rect 282658 244861 282686 256045
rect 282754 250855 282782 265813
rect 282850 253339 282878 266997
rect 282946 263287 282974 275488
rect 283426 268467 283454 275502
rect 284386 275488 284688 275516
rect 283510 272161 283562 272167
rect 283510 272103 283562 272109
rect 283414 268461 283466 268467
rect 283414 268403 283466 268409
rect 283126 265057 283178 265063
rect 283126 264999 283178 265005
rect 282934 263281 282986 263287
rect 282934 263223 282986 263229
rect 282934 254549 282986 254555
rect 282934 254491 282986 254497
rect 282836 253330 282892 253339
rect 282836 253265 282892 253274
rect 282838 253217 282890 253223
rect 282838 253159 282890 253165
rect 282742 250849 282794 250855
rect 282742 250791 282794 250797
rect 282742 250553 282794 250559
rect 282742 250495 282794 250501
rect 282754 249639 282782 250495
rect 282740 249630 282796 249639
rect 282740 249565 282796 249574
rect 282850 249468 282878 253159
rect 282754 249440 282878 249468
rect 282754 245305 282782 249440
rect 282946 249320 282974 254491
rect 283030 253291 283082 253297
rect 283030 253233 283082 253239
rect 282850 249292 282974 249320
rect 282742 245299 282794 245305
rect 282742 245241 282794 245247
rect 282742 245151 282794 245157
rect 282742 245093 282794 245099
rect 282646 244855 282698 244861
rect 282646 244797 282698 244803
rect 282646 244633 282698 244639
rect 282646 244575 282698 244581
rect 282550 237825 282602 237831
rect 282550 237767 282602 237773
rect 282658 231171 282686 244575
rect 282646 231165 282698 231171
rect 282646 231107 282698 231113
rect 215734 229093 215786 229099
rect 215734 229035 215786 229041
rect 282262 229093 282314 229099
rect 282262 229035 282314 229041
rect 215746 223864 215774 229035
rect 282754 228581 282782 245093
rect 282850 229469 282878 249292
rect 283042 249172 283070 253233
rect 283138 251003 283166 264999
rect 283318 264465 283370 264471
rect 283318 264407 283370 264413
rect 283222 255363 283274 255369
rect 283222 255305 283274 255311
rect 283126 250997 283178 251003
rect 283126 250939 283178 250945
rect 283126 250849 283178 250855
rect 283126 250791 283178 250797
rect 282946 249144 283070 249172
rect 282838 229463 282890 229469
rect 282838 229405 282890 229411
rect 282946 229173 282974 249144
rect 283138 249024 283166 250791
rect 283042 248996 283166 249024
rect 283042 244732 283070 248996
rect 283124 248890 283180 248899
rect 283124 248825 283180 248834
rect 283138 244880 283166 248825
rect 283234 245028 283262 255305
rect 283330 251151 283358 264407
rect 283414 255067 283466 255073
rect 283414 255009 283466 255015
rect 283318 251145 283370 251151
rect 283318 251087 283370 251093
rect 283318 250997 283370 251003
rect 283318 250939 283370 250945
rect 283330 245157 283358 250939
rect 283318 245151 283370 245157
rect 283318 245093 283370 245099
rect 283234 245000 283358 245028
rect 283138 244852 283262 244880
rect 283042 244704 283166 244732
rect 283030 244559 283082 244565
rect 283030 244501 283082 244507
rect 283042 243127 283070 244501
rect 283028 243118 283084 243127
rect 283028 243053 283084 243062
rect 283138 233317 283166 244704
rect 283126 233311 283178 233317
rect 283126 233253 283178 233259
rect 283234 233169 283262 244852
rect 283222 233163 283274 233169
rect 283222 233105 283274 233111
rect 283330 230283 283358 245000
rect 283426 232799 283454 255009
rect 283522 233243 283550 272103
rect 283700 266798 283756 266807
rect 283700 266733 283756 266742
rect 283606 256399 283658 256405
rect 283606 256341 283658 256347
rect 283510 233237 283562 233243
rect 283510 233179 283562 233185
rect 283414 232793 283466 232799
rect 283414 232735 283466 232741
rect 283318 230277 283370 230283
rect 283318 230219 283370 230225
rect 282934 229167 282986 229173
rect 282934 229109 282986 229115
rect 282742 228575 282794 228581
rect 282742 228517 282794 228523
rect 283618 228507 283646 256341
rect 283714 251267 283742 266733
rect 283796 266502 283852 266511
rect 283796 266437 283852 266446
rect 283700 251258 283756 251267
rect 283700 251193 283756 251202
rect 283702 251145 283754 251151
rect 283702 251087 283754 251093
rect 283714 238719 283742 251087
rect 283810 250231 283838 266437
rect 283892 266354 283948 266363
rect 283892 266289 283948 266298
rect 283796 250222 283852 250231
rect 283796 250157 283852 250166
rect 283906 249047 283934 266289
rect 284386 257737 284414 275488
rect 285622 267129 285674 267135
rect 285622 267071 285674 267077
rect 284566 259285 284618 259291
rect 284566 259227 284618 259233
rect 284374 257731 284426 257737
rect 284374 257673 284426 257679
rect 284086 255955 284138 255961
rect 284086 255897 284138 255903
rect 283990 254475 284042 254481
rect 283990 254417 284042 254423
rect 283892 249038 283948 249047
rect 283892 248973 283948 248982
rect 283894 248925 283946 248931
rect 283894 248867 283946 248873
rect 283798 244855 283850 244861
rect 283798 244797 283850 244803
rect 283702 238713 283754 238719
rect 283702 238655 283754 238661
rect 283606 228501 283658 228507
rect 283606 228443 283658 228449
rect 283810 228137 283838 244797
rect 283906 238867 283934 248867
rect 283894 238861 283946 238867
rect 283894 238803 283946 238809
rect 284002 230357 284030 254417
rect 283990 230351 284042 230357
rect 283990 230293 284042 230299
rect 284098 228951 284126 255897
rect 284182 255289 284234 255295
rect 284182 255231 284234 255237
rect 284194 229247 284222 255231
rect 284278 254253 284330 254259
rect 284278 254195 284330 254201
rect 284290 244861 284318 254195
rect 284374 252847 284426 252853
rect 284374 252789 284426 252795
rect 284278 244855 284330 244861
rect 284278 244797 284330 244803
rect 284278 244707 284330 244713
rect 284278 244649 284330 244655
rect 284290 244163 284318 244649
rect 284276 244154 284332 244163
rect 284276 244089 284332 244098
rect 284278 244041 284330 244047
rect 284278 243983 284330 243989
rect 284182 229241 284234 229247
rect 284182 229183 284234 229189
rect 284086 228945 284138 228951
rect 284086 228887 284138 228893
rect 284290 228359 284318 243983
rect 284386 235685 284414 252789
rect 284374 235679 284426 235685
rect 284374 235621 284426 235627
rect 284578 231467 284606 259227
rect 285238 256547 285290 256553
rect 285238 256489 285290 256495
rect 285142 256473 285194 256479
rect 285142 256415 285194 256421
rect 284854 254031 284906 254037
rect 284854 253973 284906 253979
rect 284866 236869 284894 253973
rect 285046 253735 285098 253741
rect 285046 253677 285098 253683
rect 284950 253661 285002 253667
rect 284950 253603 285002 253609
rect 284962 241499 284990 253603
rect 284948 241490 285004 241499
rect 284948 241425 285004 241434
rect 285058 238645 285086 253677
rect 285046 238639 285098 238645
rect 285046 238581 285098 238587
rect 284854 236863 284906 236869
rect 284854 236805 284906 236811
rect 285154 236795 285182 256415
rect 285250 238201 285278 256489
rect 285334 256029 285386 256035
rect 285334 255971 285386 255977
rect 285238 238195 285290 238201
rect 285238 238137 285290 238143
rect 285142 236789 285194 236795
rect 285142 236731 285194 236737
rect 284566 231461 284618 231467
rect 284566 231403 284618 231409
rect 285346 230209 285374 255971
rect 285430 254697 285482 254703
rect 285430 254639 285482 254645
rect 285442 235907 285470 254639
rect 285526 254623 285578 254629
rect 285526 254565 285578 254571
rect 285430 235901 285482 235907
rect 285430 235843 285482 235849
rect 285538 235833 285566 254565
rect 285634 247821 285662 267071
rect 285826 263435 285854 275502
rect 286198 268387 286250 268393
rect 286198 268329 286250 268335
rect 285814 263429 285866 263435
rect 285814 263371 285866 263377
rect 286006 259581 286058 259587
rect 286006 259523 286058 259529
rect 285910 256769 285962 256775
rect 285910 256711 285962 256717
rect 285814 256621 285866 256627
rect 285814 256563 285866 256569
rect 285718 253883 285770 253889
rect 285718 253825 285770 253831
rect 285622 247815 285674 247821
rect 285622 247757 285674 247763
rect 285622 247667 285674 247673
rect 285622 247609 285674 247615
rect 285526 235827 285578 235833
rect 285526 235769 285578 235775
rect 285334 230203 285386 230209
rect 285334 230145 285386 230151
rect 285634 228729 285662 247609
rect 285730 230431 285758 253825
rect 285826 247544 285854 256563
rect 285922 248159 285950 256711
rect 285908 248150 285964 248159
rect 285908 248085 285964 248094
rect 286018 247840 286046 259523
rect 286102 259433 286154 259439
rect 286102 259375 286154 259381
rect 285922 247812 286046 247840
rect 285922 247673 285950 247812
rect 286006 247741 286058 247747
rect 286006 247683 286058 247689
rect 285910 247667 285962 247673
rect 285910 247609 285962 247615
rect 285826 247516 285950 247544
rect 285812 247262 285868 247271
rect 285812 247197 285868 247206
rect 285826 236943 285854 247197
rect 285814 236937 285866 236943
rect 285814 236879 285866 236885
rect 285922 231763 285950 247516
rect 286018 238275 286046 247683
rect 286006 238269 286058 238275
rect 286006 238211 286058 238217
rect 285910 231757 285962 231763
rect 285910 231699 285962 231705
rect 286114 231689 286142 259375
rect 286210 233391 286238 268329
rect 286582 266611 286634 266617
rect 286582 266553 286634 266559
rect 286390 262763 286442 262769
rect 286390 262705 286442 262711
rect 286294 255511 286346 255517
rect 286294 255453 286346 255459
rect 286198 233385 286250 233391
rect 286198 233327 286250 233333
rect 286102 231683 286154 231689
rect 286102 231625 286154 231631
rect 285718 230425 285770 230431
rect 285718 230367 285770 230373
rect 286306 228877 286334 255453
rect 286402 233095 286430 262705
rect 286486 256695 286538 256701
rect 286486 256637 286538 256643
rect 286390 233089 286442 233095
rect 286390 233031 286442 233037
rect 286294 228871 286346 228877
rect 286294 228813 286346 228819
rect 286498 228803 286526 256637
rect 286594 238497 286622 266553
rect 286870 265945 286922 265951
rect 286870 265887 286922 265893
rect 286774 265427 286826 265433
rect 286774 265369 286826 265375
rect 286678 259507 286730 259513
rect 286678 259449 286730 259455
rect 286582 238491 286634 238497
rect 286582 238433 286634 238439
rect 286690 231541 286718 259449
rect 286786 238349 286814 265369
rect 286882 238423 286910 265887
rect 287074 265507 287102 275502
rect 288226 268541 288254 275502
rect 288214 268535 288266 268541
rect 288214 268477 288266 268483
rect 288022 268461 288074 268467
rect 288022 268403 288074 268409
rect 288034 268245 288062 268403
rect 288022 268239 288074 268245
rect 288022 268181 288074 268187
rect 289270 266685 289322 266691
rect 289270 266627 289322 266633
rect 287926 266093 287978 266099
rect 287926 266035 287978 266041
rect 287158 265723 287210 265729
rect 287158 265665 287210 265671
rect 287062 265501 287114 265507
rect 287062 265443 287114 265449
rect 287170 256720 287198 265665
rect 287938 265655 287966 266035
rect 287926 265649 287978 265655
rect 287926 265591 287978 265597
rect 288790 261505 288842 261511
rect 288790 261447 288842 261453
rect 287074 256692 287198 256720
rect 286966 255215 287018 255221
rect 286966 255157 287018 255163
rect 286870 238417 286922 238423
rect 286870 238359 286922 238365
rect 286774 238343 286826 238349
rect 286774 238285 286826 238291
rect 286678 231535 286730 231541
rect 286678 231477 286730 231483
rect 286978 231097 287006 255157
rect 287074 238571 287102 256692
rect 288022 255881 288074 255887
rect 288022 255823 288074 255829
rect 287830 255141 287882 255147
rect 287830 255083 287882 255089
rect 287254 254179 287306 254185
rect 287254 254121 287306 254127
rect 287158 253957 287210 253963
rect 287158 253899 287210 253905
rect 287062 238565 287114 238571
rect 287062 238507 287114 238513
rect 287170 236203 287198 253899
rect 287266 236499 287294 254121
rect 287350 254105 287402 254111
rect 287350 254047 287402 254053
rect 287362 237609 287390 254047
rect 287638 253513 287690 253519
rect 287638 253455 287690 253461
rect 287446 253143 287498 253149
rect 287446 253085 287498 253091
rect 287350 237603 287402 237609
rect 287350 237545 287402 237551
rect 287254 236493 287306 236499
rect 287254 236435 287306 236441
rect 287458 236277 287486 253085
rect 287542 252995 287594 253001
rect 287542 252937 287594 252943
rect 287554 236425 287582 252937
rect 287650 237017 287678 253455
rect 287734 253069 287786 253075
rect 287842 253043 287870 255083
rect 287926 253365 287978 253371
rect 287926 253307 287978 253313
rect 287734 253011 287786 253017
rect 287828 253034 287884 253043
rect 287638 237011 287690 237017
rect 287638 236953 287690 236959
rect 287746 236647 287774 253011
rect 287828 252969 287884 252978
rect 287830 252921 287882 252927
rect 287830 252863 287882 252869
rect 287734 236641 287786 236647
rect 287734 236583 287786 236589
rect 287842 236573 287870 252863
rect 287938 237757 287966 253307
rect 288034 249343 288062 255823
rect 288598 255585 288650 255591
rect 288598 255527 288650 255533
rect 288118 254919 288170 254925
rect 288118 254861 288170 254867
rect 288020 249334 288076 249343
rect 288020 249269 288076 249278
rect 288130 248339 288158 254861
rect 288212 253922 288268 253931
rect 288212 253857 288268 253866
rect 288226 248751 288254 253857
rect 288310 253809 288362 253815
rect 288310 253751 288362 253757
rect 288212 248742 288268 248751
rect 288212 248677 288268 248686
rect 288322 248413 288350 253751
rect 288502 253439 288554 253445
rect 288502 253381 288554 253387
rect 288514 252983 288542 253381
rect 288418 252955 288542 252983
rect 288418 252724 288446 252955
rect 288418 252696 288542 252724
rect 288514 251119 288542 252696
rect 288500 251110 288556 251119
rect 288500 251045 288556 251054
rect 288404 249334 288460 249343
rect 288404 249269 288460 249278
rect 288310 248407 288362 248413
rect 288310 248349 288362 248355
rect 288118 248333 288170 248339
rect 288118 248275 288170 248281
rect 288212 248298 288268 248307
rect 288212 248233 288268 248242
rect 288022 248185 288074 248191
rect 288022 248127 288074 248133
rect 288034 247803 288062 248127
rect 288034 247775 288158 247803
rect 288020 242230 288076 242239
rect 288020 242165 288076 242174
rect 288034 237979 288062 242165
rect 288130 239607 288158 247775
rect 288118 239601 288170 239607
rect 288118 239543 288170 239549
rect 288226 239533 288254 248233
rect 288310 247667 288362 247673
rect 288310 247609 288362 247615
rect 288322 244787 288350 247609
rect 288310 244781 288362 244787
rect 288310 244723 288362 244729
rect 288310 244559 288362 244565
rect 288310 244501 288362 244507
rect 288322 242049 288350 244501
rect 288418 242239 288446 249269
rect 288500 248890 288556 248899
rect 288500 248825 288556 248834
rect 288514 248307 288542 248825
rect 288500 248298 288556 248307
rect 288500 248233 288556 248242
rect 288404 242230 288460 242239
rect 288404 242165 288460 242174
rect 288310 242043 288362 242049
rect 288310 241985 288362 241991
rect 288310 241821 288362 241827
rect 288310 241763 288362 241769
rect 288214 239527 288266 239533
rect 288214 239469 288266 239475
rect 288022 237973 288074 237979
rect 288022 237915 288074 237921
rect 288322 237905 288350 241763
rect 288404 240306 288460 240315
rect 288404 240241 288460 240250
rect 288418 239237 288446 240241
rect 288610 239681 288638 255527
rect 288802 252872 288830 261447
rect 288886 261209 288938 261215
rect 288886 261151 288938 261157
rect 288898 258847 288926 261151
rect 288886 258841 288938 258847
rect 288886 258783 288938 258789
rect 288886 256251 288938 256257
rect 288886 256193 288938 256199
rect 288898 253043 288926 256193
rect 289172 254810 289228 254819
rect 289172 254745 289228 254754
rect 289186 253043 289214 254745
rect 288884 253034 288940 253043
rect 288884 252969 288940 252978
rect 289172 253034 289228 253043
rect 289172 252969 289228 252978
rect 289282 252872 289310 266627
rect 289474 263213 289502 275502
rect 290626 268467 290654 275502
rect 290914 275488 291792 275516
rect 290614 268461 290666 268467
rect 290614 268403 290666 268409
rect 289556 267094 289612 267103
rect 289556 267029 289612 267038
rect 289462 263207 289514 263213
rect 289462 263149 289514 263155
rect 289462 255659 289514 255665
rect 289462 255601 289514 255607
rect 289474 253043 289502 255601
rect 289460 253034 289516 253043
rect 289460 252969 289516 252978
rect 288802 252844 288926 252872
rect 288898 252724 288926 252844
rect 288864 252696 288926 252724
rect 289234 252844 289310 252872
rect 289234 252710 289262 252844
rect 289570 252724 289598 267029
rect 289940 266946 289996 266955
rect 289940 266881 289996 266890
rect 289570 252696 289632 252724
rect 289954 252710 289982 266881
rect 290324 266650 290380 266659
rect 290324 266585 290380 266594
rect 290338 252710 290366 266585
rect 290708 265910 290764 265919
rect 290708 265845 290764 265854
rect 290722 252710 290750 265845
rect 290914 253667 290942 275488
rect 291092 265762 291148 265771
rect 291092 265697 291148 265706
rect 290998 253883 291050 253889
rect 290998 253825 291050 253831
rect 291010 253667 291038 253825
rect 290902 253661 290954 253667
rect 290902 253603 290954 253609
rect 290998 253661 291050 253667
rect 290998 253603 291050 253609
rect 291106 252724 291134 265697
rect 293026 263139 293054 275502
rect 294178 265285 294206 275502
rect 295426 268763 295454 275502
rect 295414 268757 295466 268763
rect 295414 268699 295466 268705
rect 294166 265279 294218 265285
rect 294166 265221 294218 265227
rect 293014 263133 293066 263139
rect 293014 263075 293066 263081
rect 296578 262843 296606 275502
rect 297826 272241 297854 275502
rect 297814 272235 297866 272241
rect 297814 272177 297866 272183
rect 298978 268837 299006 275502
rect 299446 273789 299498 273795
rect 299444 273754 299446 273763
rect 299498 273754 299500 273763
rect 299444 273689 299500 273698
rect 298966 268831 299018 268837
rect 298966 268773 299018 268779
rect 299542 268757 299594 268763
rect 299542 268699 299594 268705
rect 299158 268535 299210 268541
rect 299158 268477 299210 268483
rect 298774 268313 298826 268319
rect 298774 268255 298826 268261
rect 296566 262837 296618 262843
rect 296566 262779 296618 262785
rect 296950 262097 297002 262103
rect 291476 262062 291532 262071
rect 296950 262039 297002 262045
rect 291476 261997 291532 262006
rect 296566 262023 296618 262029
rect 291490 252872 291518 261997
rect 296566 261965 296618 261971
rect 296182 261949 296234 261955
rect 291764 261914 291820 261923
rect 296182 261891 296234 261897
rect 291764 261849 291820 261858
rect 295798 261875 295850 261881
rect 291072 252696 291134 252724
rect 291442 252844 291518 252872
rect 291442 252710 291470 252844
rect 291778 252724 291806 261849
rect 295798 261817 295850 261823
rect 292148 261766 292204 261775
rect 292148 261701 292204 261710
rect 291778 252696 291840 252724
rect 292162 252710 292190 261701
rect 292532 261618 292588 261627
rect 292532 261553 292588 261562
rect 292546 252710 292574 261553
rect 292916 261470 292972 261479
rect 292916 261405 292972 261414
rect 292930 252710 292958 261405
rect 293300 261322 293356 261331
rect 293300 261257 293356 261266
rect 293110 256103 293162 256109
rect 293110 256045 293162 256051
rect 293206 256103 293258 256109
rect 293206 256045 293258 256051
rect 293122 255739 293150 256045
rect 293110 255733 293162 255739
rect 293110 255675 293162 255681
rect 293218 253339 293246 256045
rect 293204 253330 293260 253339
rect 293204 253265 293260 253274
rect 293314 252724 293342 261257
rect 293972 261174 294028 261183
rect 293972 261109 294028 261118
rect 293590 254993 293642 254999
rect 293590 254935 293642 254941
rect 293602 252872 293630 254935
rect 293602 252844 293678 252872
rect 293280 252696 293342 252724
rect 293650 252710 293678 252844
rect 293986 252724 294014 261109
rect 294356 261026 294412 261035
rect 294356 260961 294412 260970
rect 293986 252696 294048 252724
rect 294370 252710 294398 260961
rect 294740 260878 294796 260887
rect 294740 260813 294796 260822
rect 294754 252710 294782 260813
rect 295124 260730 295180 260739
rect 295124 260665 295180 260674
rect 295138 252710 295166 260665
rect 295508 260582 295564 260591
rect 295508 260517 295564 260526
rect 295318 254845 295370 254851
rect 295318 254787 295370 254793
rect 295330 253043 295358 254787
rect 295316 253034 295372 253043
rect 295316 252969 295372 252978
rect 295522 252724 295550 260517
rect 295810 252872 295838 261817
rect 295810 252844 295886 252872
rect 295488 252696 295550 252724
rect 295858 252710 295886 252844
rect 296194 252724 296222 261891
rect 296578 255943 296606 261965
rect 296290 255915 296606 255943
rect 296290 253057 296318 255915
rect 296290 253029 296606 253057
rect 296194 252696 296256 252724
rect 296578 252710 296606 253029
rect 296962 252710 296990 262039
rect 297334 261283 297386 261289
rect 297334 261225 297386 261231
rect 297346 252710 297374 261225
rect 297718 260617 297770 260623
rect 297718 260559 297770 260565
rect 297730 252724 297758 260559
rect 298006 260543 298058 260549
rect 298006 260485 298058 260491
rect 298018 252872 298046 260485
rect 298390 260469 298442 260475
rect 298390 260411 298442 260417
rect 298294 254253 298346 254259
rect 298294 254195 298346 254201
rect 298306 253889 298334 254195
rect 298294 253883 298346 253889
rect 298294 253825 298346 253831
rect 298018 252844 298094 252872
rect 297696 252696 297758 252724
rect 298066 252710 298094 252844
rect 298402 252724 298430 260411
rect 298402 252696 298464 252724
rect 298786 252710 298814 268255
rect 299170 252710 299198 268477
rect 299446 260987 299498 260993
rect 299446 260929 299498 260935
rect 299458 260697 299486 260929
rect 299446 260691 299498 260697
rect 299446 260633 299498 260639
rect 299554 252710 299582 268699
rect 300130 262695 300158 275502
rect 300310 268831 300362 268837
rect 300310 268773 300362 268779
rect 300406 268831 300458 268837
rect 300406 268773 300458 268779
rect 300118 262689 300170 262695
rect 300118 262631 300170 262637
rect 299926 261431 299978 261437
rect 299926 261373 299978 261379
rect 299638 260691 299690 260697
rect 299638 260633 299690 260639
rect 299650 260443 299678 260633
rect 299636 260434 299692 260443
rect 299636 260369 299692 260378
rect 299938 252724 299966 261373
rect 300322 253020 300350 268773
rect 300418 268393 300446 268773
rect 300982 268757 301034 268763
rect 300982 268699 301034 268705
rect 300406 268387 300458 268393
rect 300406 268329 300458 268335
rect 300598 268387 300650 268393
rect 300598 268329 300650 268335
rect 300406 256177 300458 256183
rect 300406 256119 300458 256125
rect 300418 255961 300446 256119
rect 300406 255955 300458 255961
rect 300406 255897 300458 255903
rect 300502 255955 300554 255961
rect 300502 255897 300554 255903
rect 300514 255739 300542 255897
rect 300502 255733 300554 255739
rect 300502 255675 300554 255681
rect 299904 252696 299966 252724
rect 300274 252992 300350 253020
rect 300274 252710 300302 252992
rect 300610 252724 300638 268329
rect 300788 256734 300844 256743
rect 300788 256669 300844 256678
rect 300802 256405 300830 256669
rect 300790 256399 300842 256405
rect 300790 256341 300842 256347
rect 300886 255881 300938 255887
rect 300706 255813 300830 255832
rect 300886 255823 300938 255829
rect 300694 255807 300830 255813
rect 300746 255804 300830 255807
rect 300694 255749 300746 255755
rect 300802 255739 300830 255804
rect 300790 255733 300842 255739
rect 300790 255675 300842 255681
rect 300898 253297 300926 255823
rect 300886 253291 300938 253297
rect 300886 253233 300938 253239
rect 300610 252696 300672 252724
rect 300994 252710 301022 268699
rect 301282 265211 301310 275502
rect 302324 273754 302380 273763
rect 302324 273689 302380 273698
rect 302338 273467 302366 273689
rect 302324 273458 302380 273467
rect 302324 273393 302380 273402
rect 302434 268393 302462 275502
rect 302422 268387 302474 268393
rect 302422 268329 302474 268335
rect 301846 268165 301898 268171
rect 301846 268107 301898 268113
rect 301750 268091 301802 268097
rect 301750 268033 301802 268039
rect 301366 268017 301418 268023
rect 301366 267959 301418 267965
rect 301270 265205 301322 265211
rect 301270 265147 301322 265153
rect 301078 255437 301130 255443
rect 301078 255379 301130 255385
rect 301090 254481 301118 255379
rect 301078 254475 301130 254481
rect 301078 254417 301130 254423
rect 301378 252710 301406 267959
rect 301762 252710 301790 268033
rect 301858 262177 301886 268107
rect 303682 262621 303710 275502
rect 304930 268319 304958 275502
rect 306082 268763 306110 275502
rect 306070 268757 306122 268763
rect 306070 268699 306122 268705
rect 304918 268313 304970 268319
rect 304918 268255 304970 268261
rect 303670 262615 303722 262621
rect 303670 262557 303722 262563
rect 307234 262473 307262 275502
rect 308482 272315 308510 275502
rect 308470 272309 308522 272315
rect 308470 272251 308522 272257
rect 308002 268541 308222 268560
rect 307990 268535 308234 268541
rect 308042 268532 308182 268535
rect 307990 268477 308042 268483
rect 308182 268477 308234 268483
rect 309634 268023 309662 275502
rect 310678 268609 310730 268615
rect 310678 268551 310730 268557
rect 310690 268467 310718 268551
rect 310678 268461 310730 268467
rect 310678 268403 310730 268409
rect 309622 268017 309674 268023
rect 309622 267959 309674 267965
rect 310882 262547 310910 275502
rect 310870 262541 310922 262547
rect 310870 262483 310922 262489
rect 307222 262467 307274 262473
rect 307222 262409 307274 262415
rect 312034 262399 312062 275502
rect 313282 268097 313310 275502
rect 313270 268091 313322 268097
rect 313270 268033 313322 268039
rect 312404 264430 312460 264439
rect 312404 264365 312460 264374
rect 312418 264101 312446 264365
rect 312406 264095 312458 264101
rect 312406 264037 312458 264043
rect 314326 263651 314378 263657
rect 314326 263593 314378 263599
rect 312022 262393 312074 262399
rect 312022 262335 312074 262341
rect 314338 262251 314366 263593
rect 314434 262325 314462 275502
rect 315682 268393 315710 275502
rect 315670 268387 315722 268393
rect 315670 268329 315722 268335
rect 316738 268171 316766 275502
rect 316726 268165 316778 268171
rect 316726 268107 316778 268113
rect 317986 265748 318014 275502
rect 317986 265720 318590 265748
rect 318178 264980 318494 265008
rect 318070 264835 318122 264841
rect 318070 264777 318122 264783
rect 318082 263731 318110 264777
rect 318178 264693 318206 264980
rect 318262 264909 318314 264915
rect 318262 264851 318314 264857
rect 318166 264687 318218 264693
rect 318166 264629 318218 264635
rect 318070 263725 318122 263731
rect 318070 263667 318122 263673
rect 318166 263503 318218 263509
rect 318166 263445 318218 263451
rect 318178 263287 318206 263445
rect 318166 263281 318218 263287
rect 318166 263223 318218 263229
rect 318274 262917 318302 264851
rect 318466 264693 318494 264980
rect 318454 264687 318506 264693
rect 318454 264629 318506 264635
rect 318454 264095 318506 264101
rect 318454 264037 318506 264043
rect 318466 263583 318494 264037
rect 318562 263583 318590 265720
rect 318646 264613 318698 264619
rect 318646 264555 318698 264561
rect 318658 264439 318686 264555
rect 318644 264430 318700 264439
rect 318644 264365 318700 264374
rect 318454 263577 318506 263583
rect 318454 263519 318506 263525
rect 318550 263577 318602 263583
rect 318550 263519 318602 263525
rect 319138 263287 319166 275502
rect 319906 275488 320304 275516
rect 319702 273789 319754 273795
rect 319700 273754 319702 273763
rect 319754 273754 319756 273763
rect 319700 273689 319756 273698
rect 319906 267672 319934 275488
rect 319810 267644 319934 267672
rect 319126 263281 319178 263287
rect 319126 263223 319178 263229
rect 318262 262911 318314 262917
rect 318262 262853 318314 262859
rect 314422 262319 314474 262325
rect 314422 262261 314474 262267
rect 314326 262245 314378 262251
rect 314326 262187 314378 262193
rect 301846 262171 301898 262177
rect 301846 262113 301898 262119
rect 302038 262171 302090 262177
rect 302038 262113 302090 262119
rect 302050 262085 302078 262113
rect 301954 262057 302078 262085
rect 310294 262097 310346 262103
rect 301954 253020 301982 262057
rect 310294 262039 310346 262045
rect 310102 261949 310154 261955
rect 310102 261891 310154 261897
rect 303190 261727 303242 261733
rect 303190 261669 303242 261675
rect 302806 261283 302858 261289
rect 302806 261225 302858 261231
rect 302614 261209 302666 261215
rect 302614 261151 302666 261157
rect 302422 261135 302474 261141
rect 302422 261077 302474 261083
rect 302434 259069 302462 261077
rect 302518 261061 302570 261067
rect 302518 261003 302570 261009
rect 302422 259063 302474 259069
rect 302422 259005 302474 259011
rect 302530 258921 302558 261003
rect 302518 258915 302570 258921
rect 302518 258857 302570 258863
rect 302626 253020 302654 261151
rect 301954 252992 302126 253020
rect 302098 252710 302126 252992
rect 302482 252992 302654 253020
rect 302482 252710 302510 252992
rect 302818 252724 302846 261225
rect 302818 252696 302880 252724
rect 303202 252710 303230 261669
rect 303958 261653 304010 261659
rect 303958 261595 304010 261601
rect 303574 260839 303626 260845
rect 303574 260781 303626 260787
rect 303586 252710 303614 260781
rect 303970 252710 303998 261595
rect 305014 261579 305066 261585
rect 305014 261521 305066 261527
rect 304726 260691 304778 260697
rect 304726 260633 304778 260639
rect 304342 259655 304394 259661
rect 304342 259597 304394 259603
rect 304354 252724 304382 259597
rect 304738 252872 304766 260633
rect 304320 252696 304382 252724
rect 304690 252844 304766 252872
rect 304690 252710 304718 252844
rect 305026 252724 305054 261521
rect 305494 260913 305546 260919
rect 305494 260855 305546 260861
rect 305686 260913 305738 260919
rect 305686 260855 305738 260861
rect 305398 260173 305450 260179
rect 305398 260115 305450 260121
rect 305302 260099 305354 260105
rect 305302 260041 305354 260047
rect 305314 259217 305342 260041
rect 305302 259211 305354 259217
rect 305302 259153 305354 259159
rect 305410 259143 305438 260115
rect 305398 259137 305450 259143
rect 305398 259079 305450 259085
rect 305506 258995 305534 260855
rect 305590 260765 305642 260771
rect 305590 260707 305642 260713
rect 305494 258989 305546 258995
rect 305494 258931 305546 258937
rect 305602 257737 305630 260707
rect 305590 257731 305642 257737
rect 305590 257673 305642 257679
rect 305698 256424 305726 260855
rect 305782 260765 305834 260771
rect 305782 260707 305834 260713
rect 305410 256396 305726 256424
rect 305026 252696 305088 252724
rect 305410 252710 305438 256396
rect 305794 252710 305822 260707
rect 308758 260691 308810 260697
rect 308758 260633 308810 260639
rect 308374 260173 308426 260179
rect 308374 260115 308426 260121
rect 307990 260099 308042 260105
rect 307990 260041 308042 260047
rect 307222 260025 307274 260031
rect 307222 259967 307274 259973
rect 306934 259877 306986 259883
rect 306934 259819 306986 259825
rect 306550 259803 306602 259809
rect 306550 259745 306602 259751
rect 306166 259729 306218 259735
rect 306166 259671 306218 259677
rect 306178 252710 306206 259671
rect 306562 252724 306590 259745
rect 306946 252909 306974 259819
rect 306528 252696 306590 252724
rect 306898 252881 306974 252909
rect 306898 252710 306926 252881
rect 307234 252724 307262 259967
rect 307606 259951 307658 259957
rect 307606 259893 307658 259899
rect 307234 252696 307296 252724
rect 307618 252710 307646 259893
rect 308002 252710 308030 260041
rect 308386 252710 308414 260115
rect 308770 252724 308798 260633
rect 309814 260469 309866 260475
rect 309140 260434 309196 260443
rect 309814 260411 309866 260417
rect 309140 260369 309196 260378
rect 309046 260321 309098 260327
rect 309046 260263 309098 260269
rect 309058 252872 309086 260263
rect 309154 257663 309182 260369
rect 309430 260321 309482 260327
rect 309430 260263 309482 260269
rect 309142 257657 309194 257663
rect 309142 257599 309194 257605
rect 309058 252844 309134 252872
rect 308736 252696 308798 252724
rect 309106 252710 309134 252844
rect 309442 252724 309470 260263
rect 309442 252696 309504 252724
rect 309826 252710 309854 260411
rect 310114 254481 310142 261891
rect 310198 260543 310250 260549
rect 310198 260485 310250 260491
rect 310102 254475 310154 254481
rect 310102 254417 310154 254423
rect 310210 252710 310238 260485
rect 310306 254833 310334 262039
rect 311350 262023 311402 262029
rect 311350 261965 311402 261971
rect 310868 256734 310924 256743
rect 310868 256669 310924 256678
rect 310882 256405 310910 256669
rect 310964 256586 311020 256595
rect 310964 256521 311020 256530
rect 310870 256399 310922 256405
rect 310870 256341 310922 256347
rect 310978 256331 311006 256521
rect 310966 256325 311018 256331
rect 310966 256267 311018 256273
rect 310390 256177 310442 256183
rect 310442 256137 310718 256165
rect 310390 256119 310442 256125
rect 310582 256103 310634 256109
rect 310582 256045 310634 256051
rect 310594 255961 310622 256045
rect 310582 255955 310634 255961
rect 310690 255943 310718 256137
rect 310918 255955 310970 255961
rect 310690 255915 310918 255943
rect 310582 255897 310634 255903
rect 310918 255897 310970 255903
rect 310774 255585 310826 255591
rect 310870 255585 310922 255591
rect 310826 255533 310870 255536
rect 310774 255527 310922 255533
rect 310786 255508 310910 255527
rect 310306 254805 310622 254833
rect 310594 252710 310622 254805
rect 310966 254475 311018 254481
rect 310966 254417 311018 254423
rect 310978 252724 311006 254417
rect 311362 252872 311390 261965
rect 311638 261875 311690 261881
rect 311638 261817 311690 261823
rect 310944 252696 311006 252724
rect 311314 252844 311390 252872
rect 311314 252710 311342 252844
rect 311650 252724 311678 261817
rect 312022 261801 312074 261807
rect 312022 261743 312074 261749
rect 311650 252696 311712 252724
rect 312034 252710 312062 261743
rect 312790 261579 312842 261585
rect 312790 261521 312842 261527
rect 312406 260987 312458 260993
rect 312406 260929 312458 260935
rect 312418 252710 312446 260929
rect 312802 252710 312830 261521
rect 313558 261505 313610 261511
rect 313558 261447 313610 261453
rect 313270 260691 313322 260697
rect 313270 260633 313322 260639
rect 313282 260401 313310 260633
rect 313174 260395 313226 260401
rect 313174 260337 313226 260343
rect 313270 260395 313322 260401
rect 313270 260337 313322 260343
rect 313186 252724 313214 260337
rect 313570 252872 313598 261447
rect 314518 261283 314570 261289
rect 314518 261225 314570 261231
rect 313846 261061 313898 261067
rect 313846 261003 313898 261009
rect 313152 252696 313214 252724
rect 313522 252844 313598 252872
rect 313522 252710 313550 252844
rect 313858 252724 313886 261003
rect 314530 256572 314558 261225
rect 314614 261135 314666 261141
rect 314614 261077 314666 261083
rect 314242 256544 314558 256572
rect 313858 252696 313920 252724
rect 314242 252710 314270 256544
rect 314626 252710 314654 261077
rect 314996 260138 315052 260147
rect 314996 260073 315052 260082
rect 315010 252710 315038 260073
rect 319028 256882 319084 256891
rect 319028 256817 319084 256826
rect 317972 256734 318028 256743
rect 317972 256669 318028 256678
rect 317204 256586 317260 256595
rect 317204 256521 317260 256530
rect 316822 254771 316874 254777
rect 316822 254713 316874 254719
rect 316054 254475 316106 254481
rect 316054 254417 316106 254423
rect 315382 254253 315434 254259
rect 315382 254195 315434 254201
rect 315394 252724 315422 254195
rect 315668 254070 315724 254079
rect 315668 254005 315724 254014
rect 315682 253020 315710 254005
rect 315682 252992 315758 253020
rect 315360 252696 315422 252724
rect 315730 252710 315758 252992
rect 316066 252724 316094 254417
rect 316724 254070 316780 254079
rect 316724 254005 316780 254014
rect 316436 253774 316492 253783
rect 316436 253709 316492 253718
rect 316066 252696 316128 252724
rect 316450 252710 316478 253709
rect 316738 253593 316766 254005
rect 316726 253587 316778 253593
rect 316726 253529 316778 253535
rect 316834 252710 316862 254713
rect 317218 252710 317246 256521
rect 317590 254327 317642 254333
rect 317590 254269 317642 254275
rect 317602 252724 317630 254269
rect 317986 252872 318014 256669
rect 318262 254401 318314 254407
rect 318262 254343 318314 254349
rect 317568 252696 317630 252724
rect 317938 252844 318014 252872
rect 317938 252710 317966 252844
rect 318274 252724 318302 254343
rect 318644 253478 318700 253487
rect 318644 253413 318700 253422
rect 318274 252696 318336 252724
rect 318658 252710 318686 253413
rect 319042 252710 319070 256817
rect 319700 256142 319756 256151
rect 319700 256077 319756 256086
rect 319714 254227 319742 256077
rect 319810 255092 319838 267644
rect 321538 262177 321566 275502
rect 322690 267991 322718 275502
rect 322676 267982 322732 267991
rect 322676 267917 322732 267926
rect 321526 262171 321578 262177
rect 321526 262113 321578 262119
rect 323938 261215 323966 275502
rect 325090 264915 325118 275502
rect 326338 267875 326366 275502
rect 327202 275488 327504 275516
rect 326326 267869 326378 267875
rect 326326 267811 326378 267817
rect 325078 264909 325130 264915
rect 325078 264851 325130 264857
rect 325462 263059 325514 263065
rect 325462 263001 325514 263007
rect 324118 261283 324170 261289
rect 324118 261225 324170 261231
rect 323926 261209 323978 261215
rect 323926 261151 323978 261157
rect 324130 261067 324158 261225
rect 324118 261061 324170 261067
rect 324118 261003 324170 261009
rect 325474 257293 325502 263001
rect 326326 261579 326378 261585
rect 326326 261521 326378 261527
rect 326038 261431 326090 261437
rect 326038 261373 326090 261379
rect 325462 257287 325514 257293
rect 325462 257229 325514 257235
rect 322004 257030 322060 257039
rect 322004 256965 322060 256974
rect 320180 256882 320236 256891
rect 320180 256817 320236 256826
rect 319810 255064 319934 255092
rect 319798 254993 319850 254999
rect 319798 254935 319850 254941
rect 319700 254218 319756 254227
rect 319700 254153 319756 254162
rect 319412 253774 319468 253783
rect 319412 253709 319468 253718
rect 319426 252710 319454 253709
rect 319810 252724 319838 254935
rect 319906 254925 319934 255064
rect 319894 254919 319946 254925
rect 319894 254861 319946 254867
rect 320194 252872 320222 256817
rect 320468 256142 320524 256151
rect 320468 256077 320524 256086
rect 319776 252696 319838 252724
rect 320146 252844 320222 252872
rect 320146 252710 320174 252844
rect 320482 252724 320510 256077
rect 321622 254919 321674 254925
rect 321622 254861 321674 254867
rect 320854 254845 320906 254851
rect 320854 254787 320906 254793
rect 320482 252696 320544 252724
rect 320866 252710 320894 254787
rect 321236 254218 321292 254227
rect 321236 254153 321292 254162
rect 321250 252710 321278 254153
rect 321634 252710 321662 254861
rect 322018 252724 322046 256965
rect 322294 256917 322346 256923
rect 322294 256859 322346 256865
rect 322306 255665 322334 256859
rect 325654 256843 325706 256849
rect 325654 256785 325706 256791
rect 322498 256396 322814 256424
rect 322390 256325 322442 256331
rect 322390 256267 322442 256273
rect 322402 255665 322430 256267
rect 322498 256257 322526 256396
rect 322582 256325 322634 256331
rect 322582 256267 322634 256273
rect 322486 256251 322538 256257
rect 322486 256193 322538 256199
rect 322294 255659 322346 255665
rect 322294 255601 322346 255607
rect 322390 255659 322442 255665
rect 322390 255601 322442 255607
rect 322390 254845 322442 254851
rect 322390 254787 322442 254793
rect 322402 252872 322430 254787
rect 322594 254671 322622 256267
rect 322678 256251 322730 256257
rect 322678 256193 322730 256199
rect 322580 254662 322636 254671
rect 322580 254597 322636 254606
rect 322580 254070 322636 254079
rect 322580 254005 322636 254014
rect 322594 253815 322622 254005
rect 322690 253931 322718 256193
rect 322676 253922 322732 253931
rect 322676 253857 322732 253866
rect 322486 253809 322538 253815
rect 322486 253751 322538 253757
rect 322582 253809 322634 253815
rect 322582 253751 322634 253757
rect 322498 253593 322526 253751
rect 322486 253587 322538 253593
rect 322486 253529 322538 253535
rect 322786 252872 322814 256396
rect 324214 255659 324266 255665
rect 324214 255601 324266 255607
rect 323828 254218 323884 254227
rect 323828 254153 323884 254162
rect 323444 254070 323500 254079
rect 323444 254005 323500 254014
rect 323062 253587 323114 253593
rect 323062 253529 323114 253535
rect 321984 252696 322046 252724
rect 322354 252844 322430 252872
rect 322738 252844 322814 252872
rect 322354 252710 322382 252844
rect 322738 252710 322766 252844
rect 323074 252710 323102 253529
rect 323458 252710 323486 254005
rect 323842 252710 323870 254153
rect 324226 252724 324254 255601
rect 324884 254662 324940 254671
rect 324884 254597 324940 254606
rect 324500 254366 324556 254375
rect 324500 254301 324556 254310
rect 324514 253020 324542 254301
rect 324514 252992 324590 253020
rect 324192 252696 324254 252724
rect 324562 252710 324590 252992
rect 324898 252724 324926 254597
rect 325268 254366 325324 254375
rect 325268 254301 325324 254310
rect 324898 252696 324960 252724
rect 325282 252710 325310 254301
rect 325666 252710 325694 256785
rect 326050 252710 326078 261373
rect 326338 260993 326366 261521
rect 326422 261061 326474 261067
rect 326422 261003 326474 261009
rect 326326 260987 326378 260993
rect 326326 260929 326378 260935
rect 326434 252724 326462 261003
rect 326806 260987 326858 260993
rect 326806 260929 326858 260935
rect 326818 252872 326846 260929
rect 327092 260286 327148 260295
rect 327092 260221 327148 260230
rect 326400 252696 326462 252724
rect 326770 252844 326846 252872
rect 326770 252710 326798 252844
rect 327106 252724 327134 260221
rect 327202 256923 327230 275488
rect 328738 268023 328766 275502
rect 328726 268017 328778 268023
rect 328726 267959 328778 267965
rect 328054 267869 328106 267875
rect 328054 267811 328106 267817
rect 327862 265575 327914 265581
rect 327862 265517 327914 265523
rect 327476 260434 327532 260443
rect 327476 260369 327532 260378
rect 327190 256917 327242 256923
rect 327190 256859 327242 256865
rect 327106 252696 327168 252724
rect 327490 252710 327518 260369
rect 327874 252710 327902 265517
rect 328066 263065 328094 267811
rect 328246 265649 328298 265655
rect 328246 265591 328298 265597
rect 328054 263059 328106 263065
rect 328054 263001 328106 263007
rect 328258 252710 328286 265591
rect 329302 265353 329354 265359
rect 329302 265295 329354 265301
rect 329204 265022 329260 265031
rect 329204 264957 329260 264966
rect 329218 264841 329246 264957
rect 329206 264835 329258 264841
rect 329206 264777 329258 264783
rect 328630 260691 328682 260697
rect 328630 260633 328682 260639
rect 328642 252724 328670 260633
rect 329014 256843 329066 256849
rect 329014 256785 329066 256791
rect 329026 252872 329054 256785
rect 328608 252696 328670 252724
rect 328978 252844 329054 252872
rect 328978 252710 329006 252844
rect 329314 252724 329342 265295
rect 329890 265137 329918 275502
rect 329878 265131 329930 265137
rect 329878 265073 329930 265079
rect 329410 264980 330206 265008
rect 329410 264915 329438 264980
rect 329398 264909 329450 264915
rect 329398 264851 329450 264857
rect 329494 264909 329546 264915
rect 329494 264851 329546 264857
rect 329506 264027 329534 264851
rect 329494 264021 329546 264027
rect 329494 263963 329546 263969
rect 329590 264021 329642 264027
rect 329590 263963 329642 263969
rect 329602 263583 329630 263963
rect 330178 263657 330206 264980
rect 330740 263986 330796 263995
rect 330740 263921 330796 263930
rect 330070 263651 330122 263657
rect 330070 263593 330122 263599
rect 330166 263651 330218 263657
rect 330166 263593 330218 263599
rect 329590 263577 329642 263583
rect 329590 263519 329642 263525
rect 329686 263577 329738 263583
rect 329686 263519 329738 263525
rect 329314 252696 329376 252724
rect 329698 252710 329726 263519
rect 330082 252710 330110 263593
rect 330452 262654 330508 262663
rect 330452 262589 330508 262598
rect 330466 252710 330494 262589
rect 330754 257367 330782 263921
rect 330932 263690 330988 263699
rect 330932 263625 330988 263634
rect 330836 262802 330892 262811
rect 330836 262737 330892 262746
rect 330742 257361 330794 257367
rect 330742 257303 330794 257309
rect 330850 252724 330878 262737
rect 330946 256923 330974 263625
rect 331042 261363 331070 275502
rect 332290 268097 332318 275502
rect 333442 268171 333470 275502
rect 333430 268165 333482 268171
rect 333430 268107 333482 268113
rect 332278 268091 332330 268097
rect 332278 268033 332330 268039
rect 333718 264761 333770 264767
rect 333718 264703 333770 264709
rect 333730 264619 333758 264703
rect 333718 264613 333770 264619
rect 332660 264578 332716 264587
rect 333718 264555 333770 264561
rect 332660 264513 332716 264522
rect 331124 263838 331180 263847
rect 331124 263773 331180 263782
rect 331030 261357 331082 261363
rect 331030 261299 331082 261305
rect 331138 257441 331166 263773
rect 331510 262985 331562 262991
rect 331510 262927 331562 262933
rect 331126 257435 331178 257441
rect 331126 257377 331178 257383
rect 331222 257139 331274 257145
rect 331222 257081 331274 257087
rect 330934 256917 330986 256923
rect 330934 256859 330986 256865
rect 331234 252872 331262 257081
rect 330816 252696 330878 252724
rect 331186 252844 331262 252872
rect 331186 252710 331214 252844
rect 331522 252724 331550 262927
rect 332276 262506 332332 262515
rect 332276 262441 332332 262450
rect 331894 257509 331946 257515
rect 331894 257451 331946 257457
rect 331522 252696 331584 252724
rect 331906 252710 331934 257451
rect 332290 252710 332318 262441
rect 332674 252710 332702 264513
rect 333044 264430 333100 264439
rect 333044 264365 333100 264374
rect 333058 252724 333086 264365
rect 333428 264282 333484 264291
rect 333428 264217 333484 264226
rect 333238 263577 333290 263583
rect 333238 263519 333290 263525
rect 333250 263287 333278 263519
rect 333142 263281 333194 263287
rect 333142 263223 333194 263229
rect 333238 263281 333290 263287
rect 333238 263223 333290 263229
rect 333154 257219 333182 263223
rect 333142 257213 333194 257219
rect 333142 257155 333194 257161
rect 333442 252872 333470 264217
rect 333716 264134 333772 264143
rect 333716 264069 333772 264078
rect 333526 263059 333578 263065
rect 333526 263001 333578 263007
rect 333622 263059 333674 263065
rect 333622 263001 333674 263007
rect 333538 257293 333566 263001
rect 333634 257515 333662 263001
rect 333622 257509 333674 257515
rect 333622 257451 333674 257457
rect 333526 257287 333578 257293
rect 333526 257229 333578 257235
rect 333024 252696 333086 252724
rect 333394 252844 333470 252872
rect 333394 252710 333422 252844
rect 333730 252724 333758 264069
rect 334004 263542 334060 263551
rect 334004 263477 334060 263486
rect 334018 257483 334046 263477
rect 334102 262245 334154 262251
rect 334102 262187 334154 262193
rect 334004 257474 334060 257483
rect 334004 257409 334060 257418
rect 333730 252696 333792 252724
rect 334114 252710 334142 262187
rect 334594 261733 334622 275502
rect 335842 268245 335870 275502
rect 335830 268239 335882 268245
rect 335830 268181 335882 268187
rect 336994 267209 337022 275502
rect 337282 275488 338160 275516
rect 339408 275488 339518 275516
rect 336982 267203 337034 267209
rect 336982 267145 337034 267151
rect 335254 264539 335306 264545
rect 335254 264481 335306 264487
rect 335266 264175 335294 264481
rect 335254 264169 335306 264175
rect 335254 264111 335306 264117
rect 335350 264169 335402 264175
rect 335350 264111 335402 264117
rect 335362 263861 335390 264111
rect 335636 263986 335692 263995
rect 335636 263921 335692 263930
rect 334882 263833 335390 263861
rect 334882 263583 334910 263833
rect 335350 263651 335402 263657
rect 335350 263593 335402 263599
rect 334870 263577 334922 263583
rect 334870 263519 334922 263525
rect 334582 261727 334634 261733
rect 334582 261669 334634 261675
rect 334484 259990 334540 259999
rect 334484 259925 334540 259934
rect 334498 252710 334526 259925
rect 334870 257509 334922 257515
rect 334870 257451 334922 257457
rect 334882 252710 334910 257451
rect 335362 252872 335390 263593
rect 335650 252872 335678 263921
rect 335924 263838 335980 263847
rect 335924 263773 335980 263782
rect 335266 252844 335390 252872
rect 335602 252844 335678 252872
rect 335266 252724 335294 252844
rect 335232 252696 335294 252724
rect 335602 252710 335630 252844
rect 335938 252724 335966 263773
rect 336308 263690 336364 263699
rect 336308 263625 336364 263634
rect 335938 252696 336000 252724
rect 336322 252710 336350 263625
rect 336692 263542 336748 263551
rect 336692 263477 336748 263486
rect 336706 252710 336734 263477
rect 337078 262171 337130 262177
rect 337078 262113 337130 262119
rect 337090 252710 337118 262113
rect 337282 255591 337310 275488
rect 339490 267857 339518 275488
rect 339766 273789 339818 273795
rect 339766 273731 339818 273737
rect 339778 273615 339806 273731
rect 339764 273606 339820 273615
rect 339764 273541 339820 273550
rect 339766 268017 339818 268023
rect 339764 267982 339766 267991
rect 339818 267982 339820 267991
rect 339764 267917 339820 267926
rect 339574 267869 339626 267875
rect 339490 267829 339574 267857
rect 339574 267811 339626 267817
rect 339766 267203 339818 267209
rect 339766 267145 339818 267151
rect 337366 266981 337418 266987
rect 337366 266923 337418 266929
rect 337270 255585 337322 255591
rect 337270 255527 337322 255533
rect 337378 252872 337406 266923
rect 338708 265022 338764 265031
rect 338708 264957 338764 264966
rect 338050 264388 338654 264416
rect 338050 264175 338078 264388
rect 338626 264323 338654 264388
rect 338518 264317 338570 264323
rect 338518 264259 338570 264265
rect 338614 264317 338666 264323
rect 338614 264259 338666 264265
rect 338134 264243 338186 264249
rect 338134 264185 338186 264191
rect 338038 264169 338090 264175
rect 338038 264111 338090 264117
rect 337750 263799 337802 263805
rect 337750 263741 337802 263747
rect 337846 263799 337898 263805
rect 337846 263741 337898 263747
rect 337460 255994 337516 256003
rect 337460 255929 337516 255938
rect 337474 254671 337502 255929
rect 337460 254662 337516 254671
rect 337460 254597 337516 254606
rect 337762 252872 337790 263741
rect 337858 257145 337886 263741
rect 337846 257139 337898 257145
rect 337846 257081 337898 257087
rect 337378 252844 337502 252872
rect 337762 252844 337838 252872
rect 337474 252724 337502 252844
rect 337440 252696 337502 252724
rect 337810 252710 337838 252844
rect 338146 252724 338174 264185
rect 338230 264021 338282 264027
rect 338422 264021 338474 264027
rect 338282 263969 338422 263972
rect 338230 263963 338474 263969
rect 338242 263944 338462 263963
rect 338326 253809 338378 253815
rect 338326 253751 338378 253757
rect 338338 253593 338366 253751
rect 338326 253587 338378 253593
rect 338326 253529 338378 253535
rect 338146 252696 338208 252724
rect 338530 252710 338558 264259
rect 338722 263953 338750 264957
rect 339574 264687 339626 264693
rect 339574 264629 339626 264635
rect 339286 264613 339338 264619
rect 339286 264555 339338 264561
rect 338902 264391 338954 264397
rect 338902 264333 338954 264339
rect 338710 263947 338762 263953
rect 338710 263889 338762 263895
rect 338914 252710 338942 264333
rect 339298 252710 339326 264555
rect 339586 252872 339614 264629
rect 339778 264249 339806 267145
rect 339958 264835 340010 264841
rect 339958 264777 340010 264783
rect 339766 264243 339818 264249
rect 339766 264185 339818 264191
rect 339670 263725 339722 263731
rect 339670 263667 339722 263673
rect 339682 257515 339710 263667
rect 339670 257509 339722 257515
rect 339670 257451 339722 257457
rect 339970 252872 339998 264777
rect 340342 264761 340394 264767
rect 340342 264703 340394 264709
rect 339586 252844 339710 252872
rect 339970 252844 340046 252872
rect 339682 252724 339710 252844
rect 339648 252696 339710 252724
rect 340018 252710 340046 252844
rect 340354 252724 340382 264703
rect 340546 264101 340574 275502
rect 341686 264317 341738 264323
rect 341686 264259 341738 264265
rect 340534 264095 340586 264101
rect 340534 264037 340586 264043
rect 340726 263947 340778 263953
rect 340726 263889 340778 263895
rect 340354 252696 340416 252724
rect 340738 252710 340766 263889
rect 341110 263577 341162 263583
rect 341110 263519 341162 263525
rect 341122 252710 341150 263519
rect 341494 262911 341546 262917
rect 341494 262853 341546 262859
rect 341506 252710 341534 262853
rect 341698 253020 341726 264259
rect 341794 260845 341822 275502
rect 342070 268757 342122 268763
rect 342070 268699 342122 268705
rect 342082 268245 342110 268699
rect 342070 268239 342122 268245
rect 342070 268181 342122 268187
rect 342550 263503 342602 263509
rect 342550 263445 342602 263451
rect 342166 263355 342218 263361
rect 342166 263297 342218 263303
rect 341782 260839 341834 260845
rect 341782 260781 341834 260787
rect 341878 260839 341930 260845
rect 341878 260781 341930 260787
rect 341890 256849 341918 260781
rect 341878 256843 341930 256849
rect 341878 256785 341930 256791
rect 341698 252992 341870 253020
rect 341842 252710 341870 252992
rect 342178 252872 342206 263297
rect 342178 252844 342254 252872
rect 342226 252710 342254 252844
rect 342562 252724 342590 263445
rect 342838 263429 342890 263435
rect 342838 263371 342890 263377
rect 342850 256868 342878 263371
rect 342946 256997 342974 275502
rect 344208 275488 344606 275516
rect 344578 268139 344606 275488
rect 345058 275488 345360 275516
rect 344564 268130 344620 268139
rect 344564 268065 344620 268074
rect 344374 264909 344426 264915
rect 344374 264851 344426 264857
rect 343318 263207 343370 263213
rect 343318 263149 343370 263155
rect 342934 256991 342986 256997
rect 342934 256933 342986 256939
rect 342850 256840 342974 256868
rect 342562 252696 342624 252724
rect 342946 252710 342974 256840
rect 343330 252710 343358 263149
rect 343702 263133 343754 263139
rect 343702 263075 343754 263081
rect 343714 252710 343742 263075
rect 344086 262837 344138 262843
rect 344086 262779 344138 262785
rect 344098 252724 344126 262779
rect 344386 252872 344414 264851
rect 344758 262689 344810 262695
rect 344758 262631 344810 262637
rect 344386 252844 344462 252872
rect 344064 252696 344126 252724
rect 344434 252710 344462 252844
rect 344770 252724 344798 262631
rect 345058 254671 345086 275488
rect 346486 264021 346538 264027
rect 346486 263963 346538 263969
rect 345142 262615 345194 262621
rect 345142 262557 345194 262563
rect 345044 254662 345100 254671
rect 345044 254597 345100 254606
rect 344770 252696 344832 252724
rect 345154 252710 345182 262557
rect 345910 262541 345962 262547
rect 345910 262483 345962 262489
rect 345526 262467 345578 262473
rect 345526 262409 345578 262415
rect 345538 252710 345566 262409
rect 345922 252710 345950 262483
rect 346294 262319 346346 262325
rect 346294 262261 346346 262267
rect 346306 252724 346334 262261
rect 346498 253020 346526 263963
rect 346594 257071 346622 275502
rect 347542 267943 347594 267949
rect 347542 267885 347594 267891
rect 347350 264391 347402 264397
rect 347350 264333 347402 264339
rect 346966 262245 347018 262251
rect 346966 262187 347018 262193
rect 346582 257065 346634 257071
rect 346582 257007 346634 257013
rect 346498 252992 346670 253020
rect 346272 252696 346334 252724
rect 346642 252710 346670 252992
rect 346978 252724 347006 262187
rect 346978 252696 347040 252724
rect 347362 252710 347390 264333
rect 347554 259976 347582 267885
rect 347746 264027 347774 275502
rect 348404 273458 348460 273467
rect 348596 273458 348652 273467
rect 348460 273416 348596 273444
rect 348404 273393 348460 273402
rect 348596 273393 348652 273402
rect 348790 268757 348842 268763
rect 348790 268699 348842 268705
rect 348406 268313 348458 268319
rect 348406 268255 348458 268261
rect 348212 268130 348268 268139
rect 348118 268091 348170 268097
rect 348212 268065 348214 268074
rect 348118 268033 348170 268039
rect 348266 268065 348268 268074
rect 348214 268033 348266 268039
rect 347734 264021 347786 264027
rect 347734 263963 347786 263969
rect 347554 259948 347774 259976
rect 347746 252710 347774 259948
rect 348130 252710 348158 268033
rect 348418 268023 348446 268255
rect 348406 268017 348458 268023
rect 348406 267959 348458 267965
rect 348502 266981 348554 266987
rect 348502 266923 348554 266929
rect 348514 266025 348542 266923
rect 348502 266019 348554 266025
rect 348502 265961 348554 265967
rect 348502 263873 348554 263879
rect 348502 263815 348554 263821
rect 348514 252724 348542 263815
rect 348802 253020 348830 268699
rect 348898 261659 348926 275502
rect 350064 275488 350366 275516
rect 349270 267869 349322 267875
rect 349270 267811 349322 267817
rect 348886 261653 348938 261659
rect 348886 261595 348938 261601
rect 349282 253020 349310 267811
rect 349942 257065 349994 257071
rect 349942 257007 349994 257013
rect 349558 256991 349610 256997
rect 349558 256933 349610 256939
rect 348802 252992 348878 253020
rect 348480 252696 348542 252724
rect 348850 252710 348878 252992
rect 349234 252992 349310 253020
rect 349234 252710 349262 252992
rect 349570 252710 349598 256933
rect 349954 252710 349982 257007
rect 350338 252710 350366 275488
rect 351298 267283 351326 275502
rect 351490 275488 352464 275516
rect 351286 267277 351338 267283
rect 351286 267219 351338 267225
rect 351094 257361 351146 257367
rect 351094 257303 351146 257309
rect 350710 257139 350762 257145
rect 350710 257081 350762 257087
rect 350722 252724 350750 257081
rect 351106 252872 351134 257303
rect 351490 257187 351518 275488
rect 352918 267203 352970 267209
rect 352918 267145 352970 267151
rect 352150 264169 352202 264175
rect 352150 264111 352202 264117
rect 351476 257178 351532 257187
rect 351476 257113 351532 257122
rect 351766 256991 351818 256997
rect 351766 256933 351818 256939
rect 351382 253809 351434 253815
rect 351382 253751 351434 253757
rect 350688 252696 350750 252724
rect 351058 252844 351134 252872
rect 351058 252710 351086 252844
rect 351394 252724 351422 253751
rect 351394 252696 351456 252724
rect 351778 252710 351806 256933
rect 352162 252710 352190 264111
rect 352534 263873 352586 263879
rect 352534 263815 352586 263821
rect 352546 252710 352574 263815
rect 352930 252724 352958 267145
rect 353302 261653 353354 261659
rect 353302 261595 353354 261601
rect 353314 252872 353342 261595
rect 353602 257145 353630 275502
rect 354850 267357 354878 275502
rect 354838 267351 354890 267357
rect 354838 267293 354890 267299
rect 355798 262689 355850 262695
rect 355798 262631 355850 262637
rect 355510 262615 355562 262621
rect 355510 262557 355562 262563
rect 355126 262541 355178 262547
rect 355126 262483 355178 262489
rect 354742 262467 354794 262473
rect 354742 262409 354794 262415
rect 353974 262319 354026 262325
rect 353974 262261 354026 262267
rect 353686 262245 353738 262251
rect 353686 262187 353738 262193
rect 353590 257139 353642 257145
rect 353590 257081 353642 257087
rect 353698 252872 353726 262187
rect 352896 252696 352958 252724
rect 353266 252844 353342 252872
rect 353602 252844 353726 252872
rect 353266 252710 353294 252844
rect 353602 252724 353630 252844
rect 353602 252696 353664 252724
rect 353986 252710 354014 262261
rect 354262 261357 354314 261363
rect 354262 261299 354314 261305
rect 354274 259587 354302 261299
rect 354262 259581 354314 259587
rect 354262 259523 354314 259529
rect 354454 259581 354506 259587
rect 354454 259523 354506 259529
rect 354466 253464 354494 259523
rect 354370 253436 354494 253464
rect 354370 252710 354398 253436
rect 354754 252710 354782 262409
rect 355138 252724 355166 262483
rect 355522 253020 355550 262557
rect 355104 252696 355166 252724
rect 355474 252992 355550 253020
rect 355474 252710 355502 252992
rect 355810 252724 355838 262631
rect 356002 259661 356030 275502
rect 357264 275488 357470 275516
rect 356182 264539 356234 264545
rect 356182 264481 356234 264487
rect 355990 259655 356042 259661
rect 355990 259597 356042 259603
rect 355810 252696 355872 252724
rect 356194 252710 356222 264481
rect 357334 263133 357386 263139
rect 357334 263075 357386 263081
rect 356950 262837 357002 262843
rect 356950 262779 357002 262785
rect 356566 259655 356618 259661
rect 356566 259597 356618 259603
rect 356578 252710 356606 259597
rect 356962 252710 356990 262779
rect 357346 252724 357374 263075
rect 357442 257367 357470 275488
rect 358402 268097 358430 275502
rect 359362 275488 359664 275516
rect 358486 268831 358538 268837
rect 358486 268773 358538 268779
rect 358390 268091 358442 268097
rect 358390 268033 358442 268039
rect 358498 268023 358526 268773
rect 358486 268017 358538 268023
rect 358486 267959 358538 267965
rect 359158 263503 359210 263509
rect 359158 263445 359210 263451
rect 358774 263429 358826 263435
rect 358774 263371 358826 263377
rect 358390 263355 358442 263361
rect 358390 263297 358442 263303
rect 358006 263281 358058 263287
rect 358006 263223 358058 263229
rect 357718 263207 357770 263213
rect 357718 263149 357770 263155
rect 357430 257361 357482 257367
rect 357430 257303 357482 257309
rect 357730 252872 357758 263149
rect 357312 252696 357374 252724
rect 357682 252844 357758 252872
rect 357682 252710 357710 252844
rect 358018 252724 358046 263223
rect 358018 252696 358080 252724
rect 358402 252710 358430 263297
rect 358486 257361 358538 257367
rect 358486 257303 358538 257309
rect 358498 256849 358526 257303
rect 358486 256843 358538 256849
rect 358486 256785 358538 256791
rect 358786 252710 358814 263371
rect 359170 252710 359198 263445
rect 359362 255707 359390 275488
rect 360214 266907 360266 266913
rect 360214 266849 360266 266855
rect 359542 264909 359594 264915
rect 359542 264851 359594 264857
rect 359348 255698 359404 255707
rect 359348 255633 359404 255642
rect 359554 252724 359582 264851
rect 359926 264835 359978 264841
rect 359926 264777 359978 264783
rect 359938 252872 359966 264777
rect 360022 264095 360074 264101
rect 360022 264037 360074 264043
rect 360034 257145 360062 264037
rect 360022 257139 360074 257145
rect 360022 257081 360074 257087
rect 359520 252696 359582 252724
rect 359890 252844 359966 252872
rect 359890 252710 359918 252844
rect 360226 252724 360254 266849
rect 360598 264687 360650 264693
rect 360598 264629 360650 264635
rect 360226 252696 360288 252724
rect 360610 252710 360638 264629
rect 360802 253815 360830 275502
rect 362050 266913 362078 275502
rect 362038 266907 362090 266913
rect 362038 266849 362090 266855
rect 360982 264761 361034 264767
rect 360982 264703 361034 264709
rect 360790 253809 360842 253815
rect 360790 253751 360842 253757
rect 360994 252710 361022 264703
rect 361366 264613 361418 264619
rect 361366 264555 361418 264561
rect 361378 252710 361406 264555
rect 361750 264539 361802 264545
rect 361750 264481 361802 264487
rect 361762 252724 361790 264481
rect 362134 264391 362186 264397
rect 362134 264333 362186 264339
rect 362146 252872 362174 264333
rect 363202 260623 363230 275502
rect 364246 268757 364298 268763
rect 364246 268699 364298 268705
rect 363190 260617 363242 260623
rect 363190 260559 363242 260565
rect 362806 256103 362858 256109
rect 362806 256045 362858 256051
rect 362422 253661 362474 253667
rect 362422 253603 362474 253609
rect 361728 252696 361790 252724
rect 362098 252844 362174 252872
rect 362098 252710 362126 252844
rect 362434 252724 362462 253603
rect 362434 252696 362496 252724
rect 362818 252710 362846 256045
rect 363190 256029 363242 256035
rect 363190 255971 363242 255977
rect 363202 252710 363230 255971
rect 363958 255955 364010 255961
rect 363958 255897 364010 255903
rect 363574 255511 363626 255517
rect 363574 255453 363626 255459
rect 363586 252710 363614 255453
rect 363970 252724 363998 255897
rect 364258 255536 364286 268699
rect 364354 256997 364382 275502
rect 364438 268831 364490 268837
rect 364438 268773 364490 268779
rect 364342 256991 364394 256997
rect 364342 256933 364394 256939
rect 364450 255559 364478 268773
rect 365602 267875 365630 275502
rect 366658 268837 366686 275502
rect 366646 268831 366698 268837
rect 366646 268773 366698 268779
rect 365590 267869 365642 267875
rect 365590 267811 365642 267817
rect 367906 267135 367934 275502
rect 368566 268165 368618 268171
rect 368566 268107 368618 268113
rect 368578 267949 368606 268107
rect 368566 267943 368618 267949
rect 368566 267885 368618 267891
rect 367894 267129 367946 267135
rect 367894 267071 367946 267077
rect 368566 266981 368618 266987
rect 368566 266923 368618 266929
rect 368578 266025 368606 266923
rect 368566 266019 368618 266025
rect 368566 265961 368618 265967
rect 368662 264243 368714 264249
rect 368662 264185 368714 264191
rect 368470 264021 368522 264027
rect 368470 263963 368522 263969
rect 366838 262393 366890 262399
rect 366838 262335 366890 262341
rect 366262 261653 366314 261659
rect 366262 261595 366314 261601
rect 366274 261363 366302 261595
rect 366166 261357 366218 261363
rect 366166 261299 366218 261305
rect 366262 261357 366314 261363
rect 366262 261299 366314 261305
rect 365590 256843 365642 256849
rect 365590 256785 365642 256791
rect 365602 256627 365630 256785
rect 365878 256695 365930 256701
rect 365878 256637 365930 256643
rect 365590 256621 365642 256627
rect 365590 256563 365642 256569
rect 365398 255881 365450 255887
rect 365398 255823 365450 255829
rect 364436 255550 364492 255559
rect 364258 255508 364382 255536
rect 364246 255437 364298 255443
rect 364354 255411 364382 255508
rect 364436 255485 364492 255494
rect 364246 255379 364298 255385
rect 364340 255402 364396 255411
rect 364258 252872 364286 255379
rect 364340 255337 364396 255346
rect 364630 255363 364682 255369
rect 364630 255305 364682 255311
rect 364258 252844 364334 252872
rect 363936 252696 363998 252724
rect 364306 252710 364334 252844
rect 364642 252724 364670 255305
rect 365014 255289 365066 255295
rect 365014 255231 365066 255237
rect 364642 252696 364704 252724
rect 365026 252710 365054 255231
rect 365410 252710 365438 255823
rect 365890 254352 365918 256637
rect 365794 254324 365918 254352
rect 365794 252710 365822 254324
rect 366178 252724 366206 261299
rect 366850 256923 366878 262335
rect 367124 258806 367180 258815
rect 367124 258741 367180 258750
rect 366838 256917 366890 256923
rect 366838 256859 366890 256865
rect 366838 256769 366890 256775
rect 366838 256711 366890 256717
rect 366454 255141 366506 255147
rect 366454 255083 366506 255089
rect 366466 252872 366494 255083
rect 366466 252844 366542 252872
rect 366144 252696 366206 252724
rect 366514 252710 366542 252844
rect 366850 252724 366878 256711
rect 367138 256701 367166 258741
rect 367796 258658 367852 258667
rect 367796 258593 367852 258602
rect 367604 258510 367660 258519
rect 367604 258445 367660 258454
rect 367126 256695 367178 256701
rect 367126 256637 367178 256643
rect 367618 256627 367646 258445
rect 367810 256849 367838 258593
rect 367798 256843 367850 256849
rect 367798 256785 367850 256791
rect 368482 256775 368510 263963
rect 368566 263577 368618 263583
rect 368566 263519 368618 263525
rect 368578 263065 368606 263519
rect 368566 263059 368618 263065
rect 368566 263001 368618 263007
rect 368674 256997 368702 264185
rect 369058 262769 369086 275502
rect 370306 268763 370334 275502
rect 370294 268757 370346 268763
rect 370294 268699 370346 268705
rect 371458 264471 371486 275502
rect 372502 267795 372554 267801
rect 372502 267737 372554 267743
rect 372598 267795 372650 267801
rect 372598 267737 372650 267743
rect 372514 267135 372542 267737
rect 372610 267357 372638 267737
rect 372598 267351 372650 267357
rect 372598 267293 372650 267299
rect 372502 267129 372554 267135
rect 372502 267071 372554 267077
rect 372706 267061 372734 275502
rect 373570 275488 373872 275516
rect 372694 267055 372746 267061
rect 372694 266997 372746 267003
rect 373078 266537 373130 266543
rect 373078 266479 373130 266485
rect 371446 264465 371498 264471
rect 371446 264407 371498 264413
rect 369046 262763 369098 262769
rect 369046 262705 369098 262711
rect 369430 259507 369482 259513
rect 369430 259449 369482 259455
rect 369046 259359 369098 259365
rect 369046 259301 369098 259307
rect 368662 256991 368714 256997
rect 368662 256933 368714 256939
rect 368374 256769 368426 256775
rect 368374 256711 368426 256717
rect 368470 256769 368522 256775
rect 368470 256711 368522 256717
rect 367510 256621 367562 256627
rect 367510 256563 367562 256569
rect 367606 256621 367658 256627
rect 367606 256563 367658 256569
rect 367522 254204 367550 256563
rect 367990 255215 368042 255221
rect 367990 255157 368042 255163
rect 367522 254176 367646 254204
rect 367222 253513 367274 253519
rect 367222 253455 367274 253461
rect 366850 252696 366912 252724
rect 367234 252710 367262 253455
rect 367618 252710 367646 254176
rect 368002 252710 368030 255157
rect 368386 252724 368414 256711
rect 368662 255067 368714 255073
rect 368662 255009 368714 255015
rect 368674 252872 368702 255009
rect 368674 252844 368750 252872
rect 368352 252696 368414 252724
rect 368722 252710 368750 252844
rect 369058 252724 369086 259301
rect 369058 252696 369120 252724
rect 369442 252710 369470 259449
rect 370870 259433 370922 259439
rect 370870 259375 370922 259381
rect 370292 258362 370348 258371
rect 370292 258297 370348 258306
rect 369814 256473 369866 256479
rect 369814 256415 369866 256421
rect 369826 252710 369854 256415
rect 370306 256405 370334 258297
rect 370198 256399 370250 256405
rect 370198 256341 370250 256347
rect 370294 256399 370346 256405
rect 370294 256341 370346 256347
rect 370210 252710 370238 256341
rect 370582 253365 370634 253371
rect 370582 253307 370634 253313
rect 370594 252724 370622 253307
rect 370882 252872 370910 259375
rect 371444 258954 371500 258963
rect 371444 258889 371500 258898
rect 371458 256479 371486 258889
rect 371446 256473 371498 256479
rect 371446 256415 371498 256421
rect 371254 253217 371306 253223
rect 371254 253159 371306 253165
rect 370882 252844 370958 252872
rect 370560 252696 370622 252724
rect 370930 252710 370958 252844
rect 371266 252724 371294 253159
rect 372406 253143 372458 253149
rect 372406 253085 372458 253091
rect 371638 253069 371690 253075
rect 371638 253011 371690 253017
rect 371266 252696 371328 252724
rect 371650 252710 371678 253011
rect 372022 252921 372074 252927
rect 372022 252863 372074 252869
rect 372034 252710 372062 252863
rect 372418 252710 372446 253085
rect 372742 252995 372794 253001
rect 372742 252937 372794 252943
rect 372754 252710 372782 252937
rect 373090 252872 373118 266479
rect 373570 260919 373598 275488
rect 374806 266537 374858 266543
rect 374806 266479 374858 266485
rect 374818 266321 374846 266479
rect 374806 266315 374858 266321
rect 374806 266257 374858 266263
rect 374902 266315 374954 266321
rect 374902 266257 374954 266263
rect 374914 265137 374942 266257
rect 374902 265131 374954 265137
rect 374902 265073 374954 265079
rect 374230 264465 374282 264471
rect 374230 264407 374282 264413
rect 373846 261727 373898 261733
rect 373846 261669 373898 261675
rect 373558 260913 373610 260919
rect 373558 260855 373610 260861
rect 373462 260617 373514 260623
rect 373462 260559 373514 260565
rect 373090 252844 373166 252872
rect 373138 252710 373166 252844
rect 373474 252724 373502 260559
rect 373474 252696 373536 252724
rect 373858 252710 373886 261669
rect 374242 252710 374270 264407
rect 374998 264243 375050 264249
rect 374998 264185 375050 264191
rect 374614 261653 374666 261659
rect 374614 261595 374666 261601
rect 374626 252710 374654 261595
rect 375010 252724 375038 264185
rect 375106 263879 375134 275502
rect 376258 268763 376286 275502
rect 377520 275488 377822 275516
rect 377494 268831 377546 268837
rect 377494 268773 377546 268779
rect 376246 268757 376298 268763
rect 376246 268699 376298 268705
rect 377206 268757 377258 268763
rect 377206 268699 377258 268705
rect 376726 268165 376778 268171
rect 376726 268107 376778 268113
rect 376738 267875 376766 268107
rect 377218 268023 377246 268699
rect 377206 268017 377258 268023
rect 377206 267959 377258 267965
rect 376726 267869 376778 267875
rect 376726 267811 376778 267817
rect 377206 266759 377258 266765
rect 377206 266701 377258 266707
rect 375190 265501 375242 265507
rect 375242 265461 375422 265489
rect 375190 265443 375242 265449
rect 375394 265433 375422 265461
rect 375382 265427 375434 265433
rect 375382 265369 375434 265375
rect 375382 264317 375434 264323
rect 375382 264259 375434 264265
rect 375094 263873 375146 263879
rect 375094 263815 375146 263821
rect 375394 252872 375422 264259
rect 375670 264169 375722 264175
rect 375670 264111 375722 264117
rect 374976 252696 375038 252724
rect 375346 252844 375422 252872
rect 375346 252710 375374 252844
rect 375682 252724 375710 264111
rect 376054 264095 376106 264101
rect 376054 264037 376106 264043
rect 375682 252696 375744 252724
rect 376066 252710 376094 264037
rect 376438 264021 376490 264027
rect 376438 263963 376490 263969
rect 376450 252710 376478 263963
rect 376822 263873 376874 263879
rect 376822 263815 376874 263821
rect 376834 252710 376862 263815
rect 377218 252724 377246 266701
rect 377506 266691 377534 268773
rect 377494 266685 377546 266691
rect 377494 266627 377546 266633
rect 377590 263947 377642 263953
rect 377590 263889 377642 263895
rect 377602 252872 377630 263889
rect 377794 255263 377822 275488
rect 378562 275488 378672 275516
rect 379522 275488 379824 275516
rect 380770 275488 381072 275516
rect 378454 270755 378506 270761
rect 378454 270697 378506 270703
rect 378166 268757 378218 268763
rect 378166 268699 378218 268705
rect 378178 268319 378206 268699
rect 378166 268313 378218 268319
rect 378166 268255 378218 268261
rect 378466 268097 378494 270697
rect 378562 268153 378590 275488
rect 379522 270761 379550 275488
rect 379510 270755 379562 270761
rect 379510 270697 379562 270703
rect 378934 268239 378986 268245
rect 378934 268181 378986 268187
rect 378562 268125 378686 268153
rect 378454 268091 378506 268097
rect 378454 268033 378506 268039
rect 378550 267721 378602 267727
rect 378550 267663 378602 267669
rect 378358 267647 378410 267653
rect 378358 267589 378410 267595
rect 378070 266463 378122 266469
rect 378070 266405 378122 266411
rect 378166 266463 378218 266469
rect 378166 266405 378218 266411
rect 378082 265211 378110 266405
rect 378178 266025 378206 266405
rect 378166 266019 378218 266025
rect 378166 265961 378218 265967
rect 378070 265205 378122 265211
rect 378070 265147 378122 265153
rect 377878 259507 377930 259513
rect 377878 259449 377930 259455
rect 377780 255254 377836 255263
rect 377780 255189 377836 255198
rect 377184 252696 377246 252724
rect 377554 252844 377630 252872
rect 377554 252710 377582 252844
rect 377890 252724 377918 259449
rect 378370 259439 378398 267589
rect 378562 266987 378590 267663
rect 378550 266981 378602 266987
rect 378550 266923 378602 266929
rect 378550 266685 378602 266691
rect 378550 266627 378602 266633
rect 378562 266247 378590 266627
rect 378658 266617 378686 268125
rect 378946 268023 378974 268181
rect 380182 268165 380234 268171
rect 380180 268130 380182 268139
rect 380234 268130 380236 268139
rect 380180 268065 380236 268074
rect 378934 268017 378986 268023
rect 378934 267959 378986 267965
rect 379990 267721 380042 267727
rect 379990 267663 380042 267669
rect 378742 267647 378794 267653
rect 378742 267589 378794 267595
rect 378754 267283 378782 267589
rect 380002 267505 380030 267663
rect 379990 267499 380042 267505
rect 379990 267441 380042 267447
rect 380086 267499 380138 267505
rect 380086 267441 380138 267447
rect 378838 267351 378890 267357
rect 378838 267293 378890 267299
rect 378742 267277 378794 267283
rect 378742 267219 378794 267225
rect 378850 266913 378878 267293
rect 379798 267277 379850 267283
rect 379798 267219 379850 267225
rect 378838 266907 378890 266913
rect 378838 266849 378890 266855
rect 378742 266833 378794 266839
rect 378742 266775 378794 266781
rect 379222 266833 379274 266839
rect 379222 266775 379274 266781
rect 378646 266611 378698 266617
rect 378646 266553 378698 266559
rect 378550 266241 378602 266247
rect 378550 266183 378602 266189
rect 378754 266099 378782 266775
rect 378838 266611 378890 266617
rect 378838 266553 378890 266559
rect 378742 266093 378794 266099
rect 378742 266035 378794 266041
rect 378850 266025 378878 266553
rect 379030 266167 379082 266173
rect 379030 266109 379082 266115
rect 378838 266019 378890 266025
rect 378838 265961 378890 265967
rect 378646 265797 378698 265803
rect 378646 265739 378698 265745
rect 378658 265211 378686 265739
rect 378550 265205 378602 265211
rect 378550 265147 378602 265153
rect 378646 265205 378698 265211
rect 378646 265147 378698 265153
rect 378562 265008 378590 265147
rect 378562 264980 378878 265008
rect 378358 259433 378410 259439
rect 378358 259375 378410 259381
rect 378262 259359 378314 259365
rect 378262 259301 378314 259307
rect 377890 252696 377952 252724
rect 378274 252710 378302 259301
rect 378452 257326 378508 257335
rect 378452 257261 378508 257270
rect 378466 256923 378494 257261
rect 378742 257065 378794 257071
rect 378658 257013 378742 257016
rect 378658 257007 378794 257013
rect 378658 256988 378782 257007
rect 378850 256997 378878 264980
rect 378838 256991 378890 256997
rect 378454 256917 378506 256923
rect 378454 256859 378506 256865
rect 378550 256843 378602 256849
rect 378550 256785 378602 256791
rect 378562 256479 378590 256785
rect 378550 256473 378602 256479
rect 378550 256415 378602 256421
rect 378658 252710 378686 256988
rect 378838 256933 378890 256939
rect 379042 252710 379070 266109
rect 379126 266019 379178 266025
rect 379126 265961 379178 265967
rect 379138 259365 379166 265961
rect 379126 259359 379178 259365
rect 379126 259301 379178 259307
rect 379234 257071 379262 266775
rect 379414 266241 379466 266247
rect 379414 266183 379466 266189
rect 379222 257065 379274 257071
rect 379222 257007 379274 257013
rect 379426 252724 379454 266183
rect 379810 252872 379838 267219
rect 379392 252696 379454 252724
rect 379762 252844 379838 252872
rect 379762 252710 379790 252844
rect 380098 252724 380126 267441
rect 380470 260913 380522 260919
rect 380470 260855 380522 260861
rect 380098 252696 380160 252724
rect 380482 252710 380510 260855
rect 380770 260771 380798 275488
rect 382210 267209 382238 275502
rect 383362 268097 383390 275502
rect 384034 275488 384528 275516
rect 383350 268091 383402 268097
rect 383350 268033 383402 268039
rect 383158 267277 383210 267283
rect 383158 267219 383210 267225
rect 382198 267203 382250 267209
rect 382198 267145 382250 267151
rect 382006 267129 382058 267135
rect 382006 267071 382058 267077
rect 381238 266759 381290 266765
rect 381238 266701 381290 266707
rect 380758 260765 380810 260771
rect 380758 260707 380810 260713
rect 380854 260765 380906 260771
rect 380854 260707 380906 260713
rect 380866 252710 380894 260707
rect 381250 252710 381278 266701
rect 381622 266093 381674 266099
rect 381622 266035 381674 266041
rect 381634 252724 381662 266035
rect 382018 252872 382046 267071
rect 382198 267055 382250 267061
rect 382198 266997 382250 267003
rect 382294 267055 382346 267061
rect 382294 266997 382346 267003
rect 382210 265475 382238 266997
rect 382196 265466 382252 265475
rect 382196 265401 382252 265410
rect 381600 252696 381662 252724
rect 381970 252844 382046 252872
rect 381970 252710 381998 252844
rect 382306 252724 382334 266997
rect 382582 266981 382634 266987
rect 382582 266923 382634 266929
rect 382678 266981 382730 266987
rect 382678 266923 382730 266929
rect 382594 266765 382622 266923
rect 382582 266759 382634 266765
rect 382582 266701 382634 266707
rect 382306 252696 382368 252724
rect 382690 252710 382718 266923
rect 383170 266173 383198 267219
rect 383554 266793 383774 266821
rect 383446 266537 383498 266543
rect 383554 266525 383582 266793
rect 383746 266765 383774 266793
rect 383638 266759 383690 266765
rect 383638 266701 383690 266707
rect 383734 266759 383786 266765
rect 383734 266701 383786 266707
rect 383498 266497 383582 266525
rect 383446 266479 383498 266485
rect 383350 266463 383402 266469
rect 383350 266405 383402 266411
rect 383362 266173 383390 266405
rect 383542 266389 383594 266395
rect 383542 266331 383594 266337
rect 383158 266167 383210 266173
rect 383158 266109 383210 266115
rect 383350 266167 383402 266173
rect 383350 266109 383402 266115
rect 383446 266019 383498 266025
rect 383446 265961 383498 265967
rect 383062 265945 383114 265951
rect 383114 265905 383198 265933
rect 383062 265887 383114 265893
rect 383170 263583 383198 265905
rect 383458 265623 383486 265961
rect 383444 265614 383500 265623
rect 383444 265549 383500 265558
rect 383158 263577 383210 263583
rect 383158 263519 383210 263525
rect 383446 262763 383498 262769
rect 383446 262705 383498 262711
rect 383062 262393 383114 262399
rect 383062 262335 383114 262341
rect 383074 257275 383102 262335
rect 383074 257247 383294 257275
rect 383156 257178 383212 257187
rect 383156 257113 383212 257122
rect 383062 257065 383114 257071
rect 383062 257007 383114 257013
rect 383074 256479 383102 257007
rect 383170 256775 383198 257113
rect 383158 256769 383210 256775
rect 383158 256711 383210 256717
rect 383062 256473 383114 256479
rect 383062 256415 383114 256421
rect 383266 256017 383294 257247
rect 383074 255989 383294 256017
rect 383074 252710 383102 255989
rect 383458 255115 383486 262705
rect 383444 255106 383500 255115
rect 383444 255041 383500 255050
rect 383554 254944 383582 266331
rect 383650 259439 383678 266701
rect 383830 266463 383882 266469
rect 383830 266405 383882 266411
rect 383638 259433 383690 259439
rect 383638 259375 383690 259381
rect 383650 256553 383774 256572
rect 383638 256547 383786 256553
rect 383690 256544 383734 256547
rect 383638 256489 383690 256495
rect 383734 256489 383786 256495
rect 383458 254916 383582 254944
rect 383458 252710 383486 254916
rect 383842 252724 383870 266405
rect 384034 262769 384062 275488
rect 385762 266543 385790 275502
rect 386326 266759 386378 266765
rect 386326 266701 386378 266707
rect 385750 266537 385802 266543
rect 385750 266479 385802 266485
rect 384214 265797 384266 265803
rect 384214 265739 384266 265745
rect 384022 262763 384074 262769
rect 384022 262705 384074 262711
rect 384226 252872 384254 265739
rect 385652 265466 385708 265475
rect 385652 265401 385708 265410
rect 384500 263246 384556 263255
rect 384500 263181 384556 263190
rect 383808 252696 383870 252724
rect 384178 252844 384254 252872
rect 384178 252710 384206 252844
rect 384514 252724 384542 263181
rect 385270 259433 385322 259439
rect 385270 259375 385322 259381
rect 384886 259359 384938 259365
rect 384886 259301 384938 259307
rect 384514 252696 384576 252724
rect 384898 252710 384926 259301
rect 385282 252710 385310 259375
rect 385666 252710 385694 265401
rect 386038 264983 386090 264989
rect 386038 264925 386090 264931
rect 386050 252724 386078 264925
rect 386338 252872 386366 266701
rect 386710 266685 386762 266691
rect 386710 266627 386762 266633
rect 386338 252844 386414 252872
rect 386016 252696 386078 252724
rect 386386 252710 386414 252844
rect 386722 252724 386750 266627
rect 386914 265507 386942 275502
rect 387286 268609 387338 268615
rect 387286 268551 387338 268557
rect 386998 267869 387050 267875
rect 386998 267811 387050 267817
rect 387010 265951 387038 267811
rect 386998 265945 387050 265951
rect 386998 265887 387050 265893
rect 386902 265501 386954 265507
rect 386902 265443 386954 265449
rect 386806 263577 386858 263583
rect 386806 263519 386858 263525
rect 386818 259088 386846 263519
rect 386818 259060 387134 259088
rect 386722 252696 386784 252724
rect 387106 252710 387134 259060
rect 387298 254819 387326 268551
rect 387862 266907 387914 266913
rect 387862 266849 387914 266855
rect 387476 264726 387532 264735
rect 387476 264661 387532 264670
rect 387284 254810 387340 254819
rect 387284 254745 387340 254754
rect 387490 252710 387518 264661
rect 387874 252710 387902 266849
rect 388162 259735 388190 275502
rect 388726 268683 388778 268689
rect 388726 268625 388778 268631
rect 388534 266167 388586 266173
rect 388534 266109 388586 266115
rect 388246 260247 388298 260253
rect 388246 260189 388298 260195
rect 388150 259729 388202 259735
rect 388150 259671 388202 259677
rect 388258 252724 388286 260189
rect 388436 257326 388492 257335
rect 388436 257261 388492 257270
rect 388450 253001 388478 257261
rect 388438 252995 388490 253001
rect 388438 252937 388490 252943
rect 388546 252872 388574 266109
rect 388738 265304 388766 268625
rect 389014 268387 389066 268393
rect 389014 268329 389066 268335
rect 388918 268239 388970 268245
rect 388918 268181 388970 268187
rect 388738 265276 388862 265304
rect 388726 256991 388778 256997
rect 388726 256933 388778 256939
rect 388738 255073 388766 256933
rect 388834 255832 388862 265276
rect 388930 262251 388958 268181
rect 389026 266173 389054 268329
rect 389014 266167 389066 266173
rect 389014 266109 389066 266115
rect 389110 265205 389162 265211
rect 389110 265147 389162 265153
rect 388918 262245 388970 262251
rect 388918 262187 388970 262193
rect 389122 258644 389150 265147
rect 389314 261363 389342 275502
rect 389878 268905 389930 268911
rect 389878 268847 389930 268853
rect 389974 268905 390026 268911
rect 389974 268847 390026 268853
rect 389686 268535 389738 268541
rect 389686 268477 389738 268483
rect 389590 265427 389642 265433
rect 389590 265369 389642 265375
rect 389302 261357 389354 261363
rect 389302 261299 389354 261305
rect 389602 259365 389630 265369
rect 389590 259359 389642 259365
rect 389590 259301 389642 259307
rect 389122 258616 389342 258644
rect 388834 255804 388958 255832
rect 388726 255067 388778 255073
rect 388726 255009 388778 255015
rect 388546 252844 388622 252872
rect 388224 252696 388286 252724
rect 388594 252710 388622 252844
rect 388930 252724 388958 255804
rect 388930 252696 388992 252724
rect 389314 252710 389342 258616
rect 389698 252710 389726 268477
rect 389890 268393 389918 268847
rect 389878 268387 389930 268393
rect 389878 268329 389930 268335
rect 389780 265614 389836 265623
rect 389780 265549 389836 265558
rect 389794 265433 389822 265549
rect 389782 265427 389834 265433
rect 389782 265369 389834 265375
rect 389986 254967 390014 268847
rect 390562 268541 390590 275502
rect 391126 272235 391178 272241
rect 391126 272177 391178 272183
rect 390550 268535 390602 268541
rect 390550 268477 390602 268483
rect 390358 268461 390410 268467
rect 390358 268403 390410 268409
rect 390070 259359 390122 259365
rect 390070 259301 390122 259307
rect 389972 254958 390028 254967
rect 389972 254893 390028 254902
rect 390082 252710 390110 259301
rect 390370 253020 390398 268403
rect 390838 267351 390890 267357
rect 390658 267311 390838 267339
rect 390658 267283 390686 267311
rect 390838 267293 390890 267299
rect 390646 267277 390698 267283
rect 390646 267219 390698 267225
rect 390742 265279 390794 265285
rect 390742 265221 390794 265227
rect 390370 252992 390446 253020
rect 390418 252710 390446 252992
rect 390754 252872 390782 265221
rect 390754 252844 390830 252872
rect 390802 252710 390830 252844
rect 391138 252724 391166 272177
rect 391714 268911 391742 275502
rect 392662 272309 392714 272315
rect 392662 272251 392714 272257
rect 391702 268905 391754 268911
rect 391702 268847 391754 268853
rect 391798 268461 391850 268467
rect 391798 268403 391850 268409
rect 391810 262325 391838 268403
rect 392278 266167 392330 266173
rect 392278 266109 392330 266115
rect 391894 265205 391946 265211
rect 391894 265147 391946 265153
rect 391798 262319 391850 262325
rect 391798 262261 391850 262267
rect 391604 259102 391660 259111
rect 391604 259037 391660 259046
rect 391618 256775 391646 259037
rect 391606 256769 391658 256775
rect 391606 256711 391658 256717
rect 391510 255067 391562 255073
rect 391510 255009 391562 255015
rect 391138 252696 391200 252724
rect 391522 252710 391550 255009
rect 391906 252710 391934 265147
rect 392290 252710 392318 266109
rect 392674 252724 392702 272251
rect 392866 265729 392894 275502
rect 393910 268757 393962 268763
rect 393910 268699 393962 268705
rect 393334 268313 393386 268319
rect 393334 268255 393386 268261
rect 393046 267055 393098 267061
rect 393046 266997 393098 267003
rect 393058 266765 393086 266997
rect 393046 266759 393098 266765
rect 393046 266701 393098 266707
rect 392854 265723 392906 265729
rect 392854 265665 392906 265671
rect 393046 257065 393098 257071
rect 393046 257007 393098 257013
rect 393058 256479 393086 257007
rect 393046 256473 393098 256479
rect 393046 256415 393098 256421
rect 392998 252995 393050 253001
rect 392998 252937 393050 252943
rect 392640 252696 392702 252724
rect 393010 252710 393038 252937
rect 393346 252724 393374 268255
rect 393430 266537 393482 266543
rect 393430 266479 393482 266485
rect 393442 266395 393470 266479
rect 393430 266389 393482 266395
rect 393430 266331 393482 266337
rect 393922 259828 393950 268699
rect 394114 265877 394142 275502
rect 395062 268017 395114 268023
rect 395062 267959 395114 267965
rect 394582 267943 394634 267949
rect 394582 267885 394634 267891
rect 394102 265871 394154 265877
rect 394102 265813 394154 265819
rect 394594 265211 394622 267885
rect 394870 266315 394922 266321
rect 394870 266257 394922 266263
rect 394582 265205 394634 265211
rect 394582 265147 394634 265153
rect 393922 259800 394142 259828
rect 393718 257213 393770 257219
rect 393718 257155 393770 257161
rect 393346 252696 393408 252724
rect 393730 252710 393758 257155
rect 394114 252710 394142 259800
rect 394486 257287 394538 257293
rect 394486 257229 394538 257235
rect 394498 252710 394526 257229
rect 394882 252724 394910 266257
rect 395074 252872 395102 267959
rect 395266 259809 395294 275502
rect 396514 268245 396542 275502
rect 397666 268911 397694 275502
rect 397654 268905 397706 268911
rect 397654 268847 397706 268853
rect 398914 268583 398942 275502
rect 398900 268574 398956 268583
rect 398900 268509 398956 268518
rect 398806 268387 398858 268393
rect 398806 268329 398858 268335
rect 396502 268239 396554 268245
rect 396502 268181 396554 268187
rect 398132 268130 398188 268139
rect 398132 268065 398188 268074
rect 397750 267795 397802 267801
rect 397750 267737 397802 267743
rect 397558 267647 397610 267653
rect 397558 267589 397610 267595
rect 395542 267425 395594 267431
rect 395542 267367 395594 267373
rect 395254 259803 395306 259809
rect 395254 259745 395306 259751
rect 395074 252844 395246 252872
rect 394848 252696 394910 252724
rect 395218 252710 395246 252844
rect 395554 252724 395582 267367
rect 397462 267351 397514 267357
rect 397462 267293 397514 267299
rect 397474 266617 397502 267293
rect 397462 266611 397514 266617
rect 397462 266553 397514 266559
rect 396694 265945 396746 265951
rect 396694 265887 396746 265893
rect 396310 257139 396362 257145
rect 396310 257081 396362 257087
rect 395926 256843 395978 256849
rect 395926 256785 395978 256791
rect 395554 252696 395616 252724
rect 395938 252710 395966 256785
rect 396322 252710 396350 257081
rect 396706 252710 396734 265887
rect 397076 257178 397132 257187
rect 397076 257113 397132 257122
rect 397090 252724 397118 257113
rect 397570 253020 397598 267589
rect 397654 266611 397706 266617
rect 397654 266553 397706 266559
rect 397666 262399 397694 266553
rect 397654 262393 397706 262399
rect 397654 262335 397706 262341
rect 397056 252696 397118 252724
rect 397426 252992 397598 253020
rect 397426 252710 397454 252992
rect 397762 252724 397790 267737
rect 397762 252696 397824 252724
rect 398146 252710 398174 268065
rect 398818 267283 398846 268329
rect 399574 268165 399626 268171
rect 399574 268107 399626 268113
rect 399382 267721 399434 267727
rect 399382 267663 399434 267669
rect 398998 267499 399050 267505
rect 398998 267441 399050 267447
rect 398422 267277 398474 267283
rect 398422 267219 398474 267225
rect 398806 267277 398858 267283
rect 398806 267219 398858 267225
rect 398434 259680 398462 267219
rect 398806 267129 398858 267135
rect 398806 267071 398858 267077
rect 398818 266839 398846 267071
rect 399010 266987 399038 267441
rect 399094 267425 399146 267431
rect 399094 267367 399146 267373
rect 399106 267209 399134 267367
rect 399094 267203 399146 267209
rect 399094 267145 399146 267151
rect 399190 267129 399242 267135
rect 399190 267071 399242 267077
rect 398998 266981 399050 266987
rect 398998 266923 399050 266929
rect 398518 266833 398570 266839
rect 398518 266775 398570 266781
rect 398806 266833 398858 266839
rect 398806 266775 398858 266781
rect 398530 266025 398558 266775
rect 398806 266389 398858 266395
rect 398806 266331 398858 266337
rect 398518 266019 398570 266025
rect 398518 265961 398570 265967
rect 398818 265803 398846 266331
rect 399202 266247 399230 267071
rect 399190 266241 399242 266247
rect 399190 266183 399242 266189
rect 398806 265797 398858 265803
rect 398806 265739 398858 265745
rect 398902 265205 398954 265211
rect 398902 265147 398954 265153
rect 398434 259652 398558 259680
rect 398530 252710 398558 259652
rect 398914 252710 398942 265147
rect 399394 252872 399422 267663
rect 399298 252844 399422 252872
rect 399586 252872 399614 268107
rect 399862 268091 399914 268097
rect 399862 268033 399914 268039
rect 399874 252872 399902 268033
rect 399970 267357 399998 275502
rect 400726 268905 400778 268911
rect 400726 268847 400778 268853
rect 400342 268535 400394 268541
rect 400342 268477 400394 268483
rect 399958 267351 400010 267357
rect 399958 267293 400010 267299
rect 399586 252844 399662 252872
rect 399874 252844 399998 252872
rect 399298 252724 399326 252844
rect 399264 252696 399326 252724
rect 399634 252710 399662 252844
rect 399970 252724 399998 252844
rect 399970 252696 400032 252724
rect 400354 252710 400382 268477
rect 400738 252710 400766 268847
rect 401218 268583 401246 275502
rect 401494 268905 401546 268911
rect 401494 268847 401546 268853
rect 401204 268574 401260 268583
rect 401204 268509 401260 268518
rect 401110 257287 401162 257293
rect 401110 257229 401162 257235
rect 401122 252710 401150 257229
rect 401506 252724 401534 268847
rect 401878 267943 401930 267949
rect 401878 267885 401930 267891
rect 401890 253020 401918 267885
rect 402166 267425 402218 267431
rect 402166 267367 402218 267373
rect 401472 252696 401534 252724
rect 401842 252992 401918 253020
rect 401842 252710 401870 252992
rect 402178 252724 402206 267367
rect 402370 259735 402398 275502
rect 403124 273606 403180 273615
rect 403124 273541 403126 273550
rect 403178 273541 403180 273550
rect 403126 273509 403178 273515
rect 403618 268467 403646 275502
rect 403606 268461 403658 268467
rect 403606 268403 403658 268409
rect 402550 267795 402602 267801
rect 402550 267737 402602 267743
rect 402358 259729 402410 259735
rect 402358 259671 402410 259677
rect 402178 252696 402240 252724
rect 402562 252710 402590 267737
rect 402934 267721 402986 267727
rect 402934 267663 402986 267669
rect 402946 252710 402974 267663
rect 404086 267647 404138 267653
rect 404086 267589 404138 267595
rect 403318 267573 403370 267579
rect 403318 267515 403370 267521
rect 403330 252710 403358 267515
rect 403702 260247 403754 260253
rect 403702 260189 403754 260195
rect 403714 252724 403742 260189
rect 404098 252872 404126 267589
rect 404374 267573 404426 267579
rect 404374 267515 404426 267521
rect 403680 252696 403742 252724
rect 404050 252844 404126 252872
rect 404050 252710 404078 252844
rect 404386 252724 404414 267515
rect 404770 257293 404798 275502
rect 404854 267499 404906 267505
rect 404854 267441 404906 267447
rect 404758 257287 404810 257293
rect 404758 257229 404810 257235
rect 404866 254944 404894 267441
rect 405142 266241 405194 266247
rect 405142 266183 405194 266189
rect 404770 254916 404894 254944
rect 404386 252696 404448 252724
rect 404770 252710 404798 254916
rect 405154 252710 405182 266183
rect 405910 265279 405962 265285
rect 405910 265221 405962 265227
rect 405526 260025 405578 260031
rect 405526 259967 405578 259973
rect 405538 252710 405566 259967
rect 405922 252724 405950 265221
rect 406018 259957 406046 275502
rect 406582 268535 406634 268541
rect 406582 268477 406634 268483
rect 406006 259951 406058 259957
rect 406006 259893 406058 259899
rect 406294 259803 406346 259809
rect 406294 259745 406346 259751
rect 406306 252872 406334 259745
rect 405888 252696 405950 252724
rect 406258 252844 406334 252872
rect 406258 252710 406286 252844
rect 406594 252724 406622 268477
rect 407170 259587 407198 275502
rect 408322 268911 408350 275502
rect 408310 268905 408362 268911
rect 408310 268847 408362 268853
rect 409570 268731 409598 275502
rect 410722 273911 410750 275502
rect 410708 273902 410764 273911
rect 410708 273837 410764 273846
rect 410422 273567 410474 273573
rect 410422 273509 410474 273515
rect 410434 273319 410462 273509
rect 410420 273310 410476 273319
rect 410420 273245 410476 273254
rect 411970 272167 411998 275502
rect 411958 272161 412010 272167
rect 411958 272103 412010 272109
rect 409556 268722 409612 268731
rect 407734 268683 407786 268689
rect 407734 268625 407786 268631
rect 408982 268683 409034 268689
rect 409556 268657 409612 268666
rect 408982 268625 409034 268631
rect 407350 267277 407402 267283
rect 407350 267219 407402 267225
rect 407158 259581 407210 259587
rect 407158 259523 407210 259529
rect 406966 257287 407018 257293
rect 406966 257229 407018 257235
rect 406594 252696 406656 252724
rect 406978 252710 407006 257229
rect 407362 252710 407390 267219
rect 407746 252710 407774 268625
rect 408694 268609 408746 268615
rect 408694 268551 408746 268557
rect 408598 268387 408650 268393
rect 408598 268329 408650 268335
rect 408118 266315 408170 266321
rect 408118 266257 408170 266263
rect 408130 252724 408158 266257
rect 408610 252872 408638 268329
rect 408706 257293 408734 268551
rect 408994 268245 409022 268625
rect 408982 268239 409034 268245
rect 408982 268181 409034 268187
rect 408790 259877 408842 259883
rect 408790 259819 408842 259825
rect 408694 257287 408746 257293
rect 408694 257229 408746 257235
rect 408096 252696 408158 252724
rect 408466 252844 408638 252872
rect 408466 252710 408494 252844
rect 408802 252724 408830 259819
rect 413122 259735 413150 275502
rect 414370 262473 414398 275502
rect 415522 267949 415550 275502
rect 416674 268879 416702 275502
rect 417622 268979 417674 268985
rect 417622 268921 417674 268927
rect 416660 268870 416716 268879
rect 416660 268805 416716 268814
rect 417634 268689 417662 268921
rect 417622 268683 417674 268689
rect 417622 268625 417674 268631
rect 417826 268287 417854 275502
rect 419088 275488 419390 275516
rect 418870 269053 418922 269059
rect 418870 268995 418922 269001
rect 417812 268278 417868 268287
rect 417812 268213 417868 268222
rect 418882 268171 418910 268995
rect 418966 268979 419018 268985
rect 418966 268921 419018 268927
rect 418978 268393 419006 268921
rect 419362 268879 419390 275488
rect 419348 268870 419404 268879
rect 419348 268805 419404 268814
rect 418966 268387 419018 268393
rect 418966 268329 419018 268335
rect 418870 268165 418922 268171
rect 418870 268107 418922 268113
rect 415510 267943 415562 267949
rect 415510 267885 415562 267891
rect 418966 266907 419018 266913
rect 418966 266849 419018 266855
rect 418978 266691 419006 266849
rect 418966 266685 419018 266691
rect 418966 266627 419018 266633
rect 414358 262467 414410 262473
rect 414358 262409 414410 262415
rect 420226 260105 420254 275502
rect 421474 262547 421502 275502
rect 421654 269201 421706 269207
rect 421654 269143 421706 269149
rect 421666 264989 421694 269143
rect 422626 267431 422654 275502
rect 423572 269906 423628 269915
rect 423572 269841 423628 269850
rect 423190 269793 423242 269799
rect 423190 269735 423242 269741
rect 422614 267425 422666 267431
rect 422614 267367 422666 267373
rect 421654 264983 421706 264989
rect 421654 264925 421706 264931
rect 421462 262541 421514 262547
rect 421462 262483 421514 262489
rect 420214 260099 420266 260105
rect 420214 260041 420266 260047
rect 413110 259729 413162 259735
rect 413110 259671 413162 259677
rect 420980 259102 421036 259111
rect 420980 259037 421036 259046
rect 414740 258954 414796 258963
rect 414740 258889 414796 258898
rect 411764 258806 411820 258815
rect 411764 258741 411820 258750
rect 409556 257326 409612 257335
rect 409174 257287 409226 257293
rect 409556 257261 409612 257270
rect 409174 257229 409226 257235
rect 408980 256142 409036 256151
rect 408980 256077 409036 256086
rect 408994 255855 409022 256077
rect 408980 255846 409036 255855
rect 408980 255781 409036 255790
rect 408802 252696 408864 252724
rect 409186 252710 409214 257229
rect 409570 252710 409598 257261
rect 410708 255698 410764 255707
rect 410708 255633 410764 255642
rect 409940 255254 409996 255263
rect 409940 255189 409996 255198
rect 409954 252710 409982 255189
rect 410324 254958 410380 254967
rect 410324 254893 410380 254902
rect 410338 252724 410366 254893
rect 410722 253020 410750 255633
rect 410996 253478 411052 253487
rect 410996 253413 411052 253422
rect 410304 252696 410366 252724
rect 410674 252992 410750 253020
rect 410674 252710 410702 252992
rect 411010 252724 411038 253413
rect 411382 252847 411434 252853
rect 411382 252789 411434 252795
rect 411010 252696 411072 252724
rect 411394 252710 411422 252789
rect 411778 252710 411806 258741
rect 413204 258510 413260 258519
rect 413204 258445 413260 258454
rect 412532 258362 412588 258371
rect 412532 258297 412588 258306
rect 412150 254623 412202 254629
rect 412150 254565 412202 254571
rect 412162 252710 412190 254565
rect 412546 252724 412574 258297
rect 412916 257178 412972 257187
rect 412916 257113 412972 257122
rect 412930 252872 412958 257113
rect 412512 252696 412574 252724
rect 412882 252844 412958 252872
rect 412882 252710 412910 252844
rect 413218 252724 413246 258445
rect 414358 254697 414410 254703
rect 414358 254639 414410 254645
rect 413974 254549 414026 254555
rect 413974 254491 414026 254497
rect 413588 253182 413644 253191
rect 413588 253117 413644 253126
rect 413218 252696 413280 252724
rect 413602 252710 413630 253117
rect 413986 252710 414014 254491
rect 414370 252710 414398 254639
rect 414754 252724 414782 258889
rect 418774 258767 418826 258773
rect 418774 258709 418826 258715
rect 418870 258767 418922 258773
rect 418870 258709 418922 258715
rect 415124 258658 415180 258667
rect 415124 258593 415180 258602
rect 415138 252872 415166 258593
rect 418786 257145 418814 258709
rect 418882 258255 418910 258709
rect 418870 258249 418922 258255
rect 418870 258191 418922 258197
rect 418774 257139 418826 257145
rect 418774 257081 418826 257087
rect 419156 255550 419212 255559
rect 419156 255485 419212 255494
rect 418772 255106 418828 255115
rect 418772 255041 418828 255050
rect 417620 254810 417676 254819
rect 417620 254745 417676 254754
rect 416180 253774 416236 253783
rect 416180 253709 416236 253718
rect 415412 253034 415468 253043
rect 415412 252969 415468 252978
rect 415796 253034 415852 253043
rect 415796 252969 415852 252978
rect 414720 252696 414782 252724
rect 415090 252844 415166 252872
rect 415090 252710 415118 252844
rect 415426 252724 415454 252969
rect 415426 252696 415488 252724
rect 415810 252710 415838 252969
rect 416194 252710 416222 253709
rect 416950 253143 417002 253149
rect 416950 253085 417002 253091
rect 416566 252921 416618 252927
rect 416566 252863 416618 252869
rect 416578 252710 416606 252863
rect 416962 252724 416990 253085
rect 417286 252847 417338 252853
rect 417286 252789 417338 252795
rect 416928 252696 416990 252724
rect 417298 252710 417326 252789
rect 417634 252724 417662 254745
rect 418388 253922 418444 253931
rect 418388 253857 418444 253866
rect 418006 253217 418058 253223
rect 418006 253159 418058 253165
rect 417634 252696 417696 252724
rect 418018 252710 418046 253159
rect 418402 252710 418430 253857
rect 418786 252710 418814 255041
rect 419170 252724 419198 255485
rect 419828 255402 419884 255411
rect 419828 255337 419884 255346
rect 419540 253626 419596 253635
rect 419540 253561 419596 253570
rect 419554 252872 419582 253561
rect 419136 252696 419198 252724
rect 419506 252844 419582 252872
rect 419506 252710 419534 252844
rect 419842 252724 419870 255337
rect 420214 254031 420266 254037
rect 420214 253973 420266 253979
rect 419842 252696 419904 252724
rect 420226 252710 420254 253973
rect 420598 253883 420650 253889
rect 420598 253825 420650 253831
rect 420610 252710 420638 253825
rect 420994 252710 421022 259037
rect 423202 257071 423230 269735
rect 423478 269719 423530 269725
rect 423478 269661 423530 269667
rect 423382 269645 423434 269651
rect 423382 269587 423434 269593
rect 423286 268387 423338 268393
rect 423286 268329 423338 268335
rect 423298 265285 423326 268329
rect 423286 265279 423338 265285
rect 423286 265221 423338 265227
rect 423394 258181 423422 269587
rect 423382 258175 423434 258181
rect 423382 258117 423434 258123
rect 423190 257065 423242 257071
rect 423190 257007 423242 257013
rect 423490 256997 423518 269661
rect 423586 263583 423614 269841
rect 423778 269027 423806 275502
rect 424438 270385 424490 270391
rect 424438 270327 424490 270333
rect 424246 270163 424298 270169
rect 424246 270105 424298 270111
rect 423764 269018 423820 269027
rect 423764 268953 423820 268962
rect 423670 267351 423722 267357
rect 423670 267293 423722 267299
rect 423574 263577 423626 263583
rect 423574 263519 423626 263525
rect 423682 257293 423710 267293
rect 424258 261363 424286 270105
rect 424450 267431 424478 270327
rect 424822 270163 424874 270169
rect 424822 270105 424874 270111
rect 424438 267425 424490 267431
rect 424438 267367 424490 267373
rect 424834 265359 424862 270105
rect 425026 268435 425054 275502
rect 425782 269941 425834 269947
rect 425782 269883 425834 269889
rect 425686 268461 425738 268467
rect 425012 268426 425068 268435
rect 425686 268403 425738 268409
rect 425012 268361 425068 268370
rect 424918 268313 424970 268319
rect 424918 268255 424970 268261
rect 424822 265353 424874 265359
rect 424822 265295 424874 265301
rect 424246 261357 424298 261363
rect 424246 261299 424298 261305
rect 424930 260031 424958 268255
rect 425590 265057 425642 265063
rect 425590 264999 425642 265005
rect 424918 260025 424970 260031
rect 424918 259967 424970 259973
rect 425014 259285 425066 259291
rect 425014 259227 425066 259233
rect 423670 257287 423722 257293
rect 423670 257229 423722 257235
rect 423478 256991 423530 256997
rect 423478 256933 423530 256939
rect 424628 256438 424684 256447
rect 424628 256373 424684 256382
rect 424244 256290 424300 256299
rect 424244 256225 424300 256234
rect 424436 256290 424492 256299
rect 424436 256225 424492 256234
rect 422422 256177 422474 256183
rect 422422 256119 422474 256125
rect 421558 255955 421610 255961
rect 421558 255897 421610 255903
rect 421570 255855 421598 255897
rect 421556 255846 421612 255855
rect 421556 255781 421612 255790
rect 421748 255846 421804 255855
rect 421748 255781 421804 255790
rect 421366 254179 421418 254185
rect 421366 254121 421418 254127
rect 421378 252724 421406 254121
rect 421762 252872 421790 255781
rect 422038 254105 422090 254111
rect 422038 254047 422090 254053
rect 421344 252696 421406 252724
rect 421714 252844 421790 252872
rect 421714 252710 421742 252844
rect 422050 252724 422078 254047
rect 422050 252696 422112 252724
rect 422434 252710 422462 256119
rect 423478 255881 423530 255887
rect 423478 255823 423530 255829
rect 423490 255684 423518 255823
rect 423862 255807 423914 255813
rect 423862 255749 423914 255755
rect 423394 255665 423518 255684
rect 423382 255659 423518 255665
rect 423434 255656 423518 255659
rect 423382 255601 423434 255607
rect 423190 253957 423242 253963
rect 423190 253899 423242 253905
rect 422806 253735 422858 253741
rect 422806 253677 422858 253683
rect 422818 252710 422846 253677
rect 423202 252710 423230 253899
rect 423574 253069 423626 253075
rect 423574 253011 423626 253017
rect 423586 252724 423614 253011
rect 423874 252872 423902 255749
rect 423874 252844 423950 252872
rect 423552 252696 423614 252724
rect 423922 252710 423950 252844
rect 424258 252724 424286 256225
rect 424450 255961 424478 256225
rect 424438 255955 424490 255961
rect 424438 255897 424490 255903
rect 424258 252696 424320 252724
rect 424642 252710 424670 256373
rect 425026 252710 425054 259227
rect 425396 254514 425452 254523
rect 425396 254449 425452 254458
rect 425410 252710 425438 254449
rect 425602 253020 425630 264999
rect 425698 259809 425726 268403
rect 425686 259803 425738 259809
rect 425686 259745 425738 259751
rect 425794 256923 425822 269883
rect 425876 269758 425932 269767
rect 425876 269693 425932 269702
rect 425782 256917 425834 256923
rect 425782 256859 425834 256865
rect 425890 256849 425918 269693
rect 425974 269571 426026 269577
rect 425974 269513 426026 269519
rect 425986 257293 426014 269513
rect 426178 269027 426206 275502
rect 426934 270681 426986 270687
rect 426934 270623 426986 270629
rect 426356 270498 426412 270507
rect 426356 270433 426412 270442
rect 426262 270015 426314 270021
rect 426262 269957 426314 269963
rect 426274 269651 426302 269957
rect 426262 269645 426314 269651
rect 426262 269587 426314 269593
rect 426164 269018 426220 269027
rect 426164 268953 426220 268962
rect 426262 268683 426314 268689
rect 426262 268625 426314 268631
rect 426274 262769 426302 268625
rect 426262 262763 426314 262769
rect 426262 262705 426314 262711
rect 426370 260105 426398 270433
rect 426838 269571 426890 269577
rect 426838 269513 426890 269519
rect 426454 269349 426506 269355
rect 426454 269291 426506 269297
rect 426466 262547 426494 269291
rect 426550 268905 426602 268911
rect 426550 268847 426602 268853
rect 426562 268171 426590 268847
rect 426550 268165 426602 268171
rect 426550 268107 426602 268113
rect 426454 262541 426506 262547
rect 426454 262483 426506 262489
rect 426358 260099 426410 260105
rect 426358 260041 426410 260047
rect 426850 259999 426878 269513
rect 426836 259990 426892 259999
rect 426836 259925 426892 259934
rect 426946 257515 426974 270623
rect 427318 270089 427370 270095
rect 427318 270031 427370 270037
rect 427126 270015 427178 270021
rect 427126 269957 427178 269963
rect 427138 262663 427166 269957
rect 427222 269941 427274 269947
rect 427222 269883 427274 269889
rect 427234 262811 427262 269883
rect 427220 262802 427276 262811
rect 427220 262737 427276 262746
rect 427124 262654 427180 262663
rect 427124 262589 427180 262598
rect 426838 257509 426890 257515
rect 426068 257474 426124 257483
rect 426838 257451 426890 257457
rect 426934 257509 426986 257515
rect 426934 257451 426986 257457
rect 426068 257409 426124 257418
rect 425974 257287 426026 257293
rect 425974 257229 426026 257235
rect 425878 256843 425930 256849
rect 425878 256785 425930 256791
rect 425684 254514 425740 254523
rect 425684 254449 425740 254458
rect 425698 253487 425726 254449
rect 425684 253478 425740 253487
rect 425684 253413 425740 253422
rect 426082 253020 426110 257409
rect 426454 257361 426506 257367
rect 426454 257303 426506 257309
rect 425602 252992 425774 253020
rect 426082 252992 426158 253020
rect 425746 252710 425774 252992
rect 426130 252710 426158 252992
rect 426466 252724 426494 257303
rect 426466 252696 426528 252724
rect 426850 252710 426878 257451
rect 427222 257435 427274 257441
rect 427222 257377 427274 257383
rect 427234 252710 427262 257377
rect 427330 257219 427358 270031
rect 427426 260179 427454 275502
rect 427894 270681 427946 270687
rect 427894 270623 427946 270629
rect 427798 270089 427850 270095
rect 427798 270031 427850 270037
rect 427510 269423 427562 269429
rect 427510 269365 427562 269371
rect 427522 265729 427550 269365
rect 427702 269201 427754 269207
rect 427702 269143 427754 269149
rect 427714 266321 427742 269143
rect 427702 266315 427754 266321
rect 427702 266257 427754 266263
rect 427510 265723 427562 265729
rect 427510 265665 427562 265671
rect 427810 263065 427838 270031
rect 427798 263059 427850 263065
rect 427798 263001 427850 263007
rect 427414 260173 427466 260179
rect 427414 260115 427466 260121
rect 427906 259883 427934 270623
rect 427990 270459 428042 270465
rect 427990 270401 428042 270407
rect 427894 259877 427946 259883
rect 427894 259819 427946 259825
rect 428002 259680 428030 270401
rect 428468 270054 428524 270063
rect 428468 269989 428524 269998
rect 427906 259652 428030 259680
rect 427606 257583 427658 257589
rect 427606 257525 427658 257531
rect 427318 257213 427370 257219
rect 427318 257155 427370 257161
rect 427618 252710 427646 257525
rect 427906 257515 427934 259652
rect 427990 258175 428042 258181
rect 427990 258117 428042 258123
rect 428182 258175 428234 258181
rect 428182 258117 428234 258123
rect 427894 257509 427946 257515
rect 427894 257451 427946 257457
rect 428002 252724 428030 258117
rect 428194 256923 428222 258117
rect 428482 257663 428510 269989
rect 428578 262621 428606 275502
rect 429236 273458 429292 273467
rect 429058 273416 429236 273444
rect 429058 273319 429086 273416
rect 429236 273393 429292 273402
rect 429044 273310 429100 273319
rect 429044 273245 429100 273254
rect 429334 270459 429386 270465
rect 429334 270401 429386 270407
rect 429238 270237 429290 270243
rect 429238 270179 429290 270185
rect 428950 269645 429002 269651
rect 428950 269587 429002 269593
rect 428566 262615 428618 262621
rect 428566 262557 428618 262563
rect 428278 257657 428330 257663
rect 428278 257599 428330 257605
rect 428470 257657 428522 257663
rect 428470 257599 428522 257605
rect 428182 256917 428234 256923
rect 428182 256859 428234 256865
rect 428290 252872 428318 257599
rect 428962 256997 428990 269587
rect 429142 269349 429194 269355
rect 429142 269291 429194 269297
rect 429046 269127 429098 269133
rect 429046 269069 429098 269075
rect 429058 268985 429086 269069
rect 429046 268979 429098 268985
rect 429046 268921 429098 268927
rect 429046 268683 429098 268689
rect 429046 268625 429098 268631
rect 429058 268245 429086 268625
rect 429046 268239 429098 268245
rect 429046 268181 429098 268187
rect 429154 266067 429182 269291
rect 429140 266058 429196 266067
rect 429140 265993 429196 266002
rect 429250 265063 429278 270179
rect 429346 265655 429374 270401
rect 429622 269793 429674 269799
rect 429622 269735 429674 269741
rect 429526 269719 429578 269725
rect 429526 269661 429578 269667
rect 429430 269423 429482 269429
rect 429430 269365 429482 269371
rect 429334 265649 429386 265655
rect 429334 265591 429386 265597
rect 429442 265581 429470 269365
rect 429430 265575 429482 265581
rect 429430 265517 429482 265523
rect 429238 265057 429290 265063
rect 429238 264999 429290 265005
rect 429538 262991 429566 269661
rect 429526 262985 429578 262991
rect 429526 262927 429578 262933
rect 429634 262917 429662 269735
rect 429718 269645 429770 269651
rect 429718 269587 429770 269593
rect 429622 262911 429674 262917
rect 429622 262853 429674 262859
rect 429730 262515 429758 269587
rect 429826 267801 429854 275502
rect 430292 270646 430348 270655
rect 430292 270581 430348 270590
rect 430100 270350 430156 270359
rect 430100 270285 430156 270294
rect 429910 269867 429962 269873
rect 429910 269809 429962 269815
rect 429814 267795 429866 267801
rect 429814 267737 429866 267743
rect 429716 262506 429772 262515
rect 429716 262441 429772 262450
rect 429922 259976 429950 269809
rect 430006 268979 430058 268985
rect 430006 268921 430058 268927
rect 429442 259948 429950 259976
rect 429046 257731 429098 257737
rect 429046 257673 429098 257679
rect 428662 256991 428714 256997
rect 428662 256933 428714 256939
rect 428950 256991 429002 256997
rect 428950 256933 429002 256939
rect 428290 252844 428366 252872
rect 427968 252696 428030 252724
rect 428338 252710 428366 252844
rect 428674 252724 428702 256933
rect 428674 252696 428736 252724
rect 429058 252710 429086 257673
rect 429442 252710 429470 259948
rect 430018 259661 430046 268921
rect 430006 259655 430058 259661
rect 430006 259597 430058 259603
rect 429814 259211 429866 259217
rect 429814 259153 429866 259159
rect 429718 259137 429770 259143
rect 429718 259079 429770 259085
rect 429730 256923 429758 259079
rect 429718 256917 429770 256923
rect 429718 256859 429770 256865
rect 429826 252710 429854 259153
rect 430114 259143 430142 270285
rect 430198 268905 430250 268911
rect 430198 268847 430250 268853
rect 430102 259137 430154 259143
rect 430102 259079 430154 259085
rect 430210 258625 430238 268847
rect 430102 258619 430154 258625
rect 430102 258561 430154 258567
rect 430198 258619 430250 258625
rect 430198 258561 430250 258567
rect 430114 257737 430142 258561
rect 430102 257731 430154 257737
rect 430102 257673 430154 257679
rect 430306 257589 430334 270581
rect 430486 268091 430538 268097
rect 430486 268033 430538 268039
rect 430498 266247 430526 268033
rect 430486 266241 430538 266247
rect 430486 266183 430538 266189
rect 430390 263577 430442 263583
rect 430390 263519 430442 263525
rect 430294 257583 430346 257589
rect 430294 257525 430346 257531
rect 430402 252872 430430 263519
rect 430978 262959 431006 275502
rect 432118 270237 432170 270243
rect 432226 270211 432254 275502
rect 433078 270607 433130 270613
rect 433078 270549 433130 270555
rect 432694 270459 432746 270465
rect 432694 270401 432746 270407
rect 432310 270385 432362 270391
rect 432310 270327 432362 270333
rect 432118 270179 432170 270185
rect 432212 270202 432268 270211
rect 431158 269867 431210 269873
rect 431158 269809 431210 269815
rect 431170 269429 431198 269809
rect 431158 269423 431210 269429
rect 431158 269365 431210 269371
rect 432022 269423 432074 269429
rect 432022 269365 432074 269371
rect 431156 269314 431212 269323
rect 431156 269249 431212 269258
rect 430964 262950 431020 262959
rect 430964 262885 431020 262894
rect 430870 261357 430922 261363
rect 430870 261299 430922 261305
rect 430486 258989 430538 258995
rect 430486 258931 430538 258937
rect 430210 252844 430430 252872
rect 430498 252872 430526 258931
rect 430498 252844 430574 252872
rect 430210 252724 430238 252844
rect 430176 252696 430238 252724
rect 430546 252710 430574 252844
rect 430882 252724 430910 261299
rect 431170 260179 431198 269249
rect 431638 267425 431690 267431
rect 431638 267367 431690 267373
rect 431158 260173 431210 260179
rect 431158 260115 431210 260121
rect 431254 256917 431306 256923
rect 431254 256859 431306 256865
rect 430882 252696 430944 252724
rect 431266 252710 431294 256859
rect 431650 252710 431678 267367
rect 432034 266215 432062 269365
rect 432020 266206 432076 266215
rect 432020 266141 432076 266150
rect 432130 265771 432158 270179
rect 432212 270137 432268 270146
rect 432322 265919 432350 270327
rect 432406 270311 432458 270317
rect 432406 270253 432458 270259
rect 432308 265910 432364 265919
rect 432308 265845 432364 265854
rect 432116 265762 432172 265771
rect 432116 265697 432172 265706
rect 432418 259976 432446 270253
rect 432706 269873 432734 270401
rect 432788 270054 432844 270063
rect 432788 269989 432844 269998
rect 432694 269867 432746 269873
rect 432694 269809 432746 269815
rect 432502 264983 432554 264989
rect 432502 264925 432554 264931
rect 432034 259948 432446 259976
rect 432034 252710 432062 259948
rect 432514 252872 432542 264925
rect 432802 260031 432830 269989
rect 432790 260025 432842 260031
rect 432790 259967 432842 259973
rect 432694 258915 432746 258921
rect 432694 258857 432746 258863
rect 432418 252844 432542 252872
rect 432706 252872 432734 258857
rect 432706 252844 432782 252872
rect 432418 252724 432446 252844
rect 432384 252696 432446 252724
rect 432754 252710 432782 252844
rect 433090 252724 433118 270549
rect 433282 269767 433310 275502
rect 433268 269758 433324 269767
rect 433268 269693 433324 269702
rect 433460 269462 433516 269471
rect 433460 269397 433516 269406
rect 433474 258995 433502 269397
rect 434530 260401 434558 275502
rect 434902 269867 434954 269873
rect 434902 269809 434954 269815
rect 434614 269053 434666 269059
rect 434614 268995 434666 269001
rect 434518 260395 434570 260401
rect 434518 260337 434570 260343
rect 433846 259211 433898 259217
rect 433846 259153 433898 259159
rect 433462 258989 433514 258995
rect 433462 258931 433514 258937
rect 433462 258841 433514 258847
rect 433462 258783 433514 258789
rect 433090 252696 433152 252724
rect 433474 252710 433502 258783
rect 433858 252710 433886 259153
rect 434228 257622 434284 257631
rect 434228 257557 434284 257566
rect 434242 252710 434270 257557
rect 434626 252724 434654 268995
rect 434914 267843 434942 269809
rect 434900 267834 434956 267843
rect 434900 267769 434956 267778
rect 434902 262763 434954 262769
rect 434902 262705 434954 262711
rect 434914 252909 434942 262705
rect 435682 262695 435710 275502
rect 436822 269275 436874 269281
rect 436822 269217 436874 269223
rect 435956 269166 436012 269175
rect 435956 269101 436012 269110
rect 435670 262689 435722 262695
rect 435670 262631 435722 262637
rect 435970 259069 435998 269101
rect 436054 260099 436106 260105
rect 436054 260041 436106 260047
rect 435958 259063 436010 259069
rect 435958 259005 436010 259011
rect 435668 258214 435724 258223
rect 435668 258149 435724 258158
rect 435284 258066 435340 258075
rect 435284 258001 435340 258010
rect 434914 252881 434990 252909
rect 434592 252696 434654 252724
rect 434962 252710 434990 252881
rect 435298 252724 435326 258001
rect 435298 252696 435360 252724
rect 435682 252710 435710 258149
rect 436066 252710 436094 260041
rect 436438 257953 436490 257959
rect 436438 257895 436490 257901
rect 436450 252710 436478 257895
rect 436834 252724 436862 269217
rect 436930 267727 436958 275502
rect 437782 273493 437834 273499
rect 437780 273458 437782 273467
rect 437834 273458 437836 273467
rect 437780 273393 437836 273402
rect 437204 269610 437260 269619
rect 437204 269545 437260 269554
rect 436918 267721 436970 267727
rect 436918 267663 436970 267669
rect 437218 258033 437246 269545
rect 437876 268426 437932 268435
rect 437876 268361 437932 268370
rect 437890 268139 437918 268361
rect 437876 268130 437932 268139
rect 437876 268065 437932 268074
rect 438082 263107 438110 275502
rect 439330 270359 439358 275502
rect 439316 270350 439372 270359
rect 439316 270285 439372 270294
rect 440086 269497 440138 269503
rect 440086 269439 440138 269445
rect 439126 268757 439178 268763
rect 439318 268757 439370 268763
rect 439178 268705 439318 268708
rect 439126 268699 439370 268705
rect 439138 268680 439358 268699
rect 438646 265723 438698 265729
rect 438646 265665 438698 265671
rect 438068 263098 438124 263107
rect 438068 263033 438124 263042
rect 437494 262541 437546 262547
rect 437494 262483 437546 262489
rect 437110 258027 437162 258033
rect 437110 257969 437162 257975
rect 437206 258027 437258 258033
rect 437206 257969 437258 257975
rect 437012 254366 437068 254375
rect 437012 254301 437068 254310
rect 437026 253487 437054 254301
rect 437012 253478 437068 253487
rect 437012 253413 437068 253422
rect 437122 252872 437150 257969
rect 437122 252844 437198 252872
rect 436800 252696 436862 252724
rect 437170 252710 437198 252844
rect 437506 252724 437534 262483
rect 437878 256843 437930 256849
rect 437878 256785 437930 256791
rect 437506 252696 437568 252724
rect 437890 252710 437918 256785
rect 438262 256695 438314 256701
rect 438262 256637 438314 256643
rect 438274 252710 438302 256637
rect 438658 252710 438686 265665
rect 439702 258693 439754 258699
rect 439702 258635 439754 258641
rect 438838 258101 438890 258107
rect 438838 258043 438890 258049
rect 438850 252909 438878 258043
rect 438934 257287 438986 257293
rect 438934 257229 438986 257235
rect 438946 253020 438974 257229
rect 439028 255254 439084 255263
rect 439028 255189 439084 255198
rect 439042 254944 439070 255189
rect 439508 254958 439564 254967
rect 439042 254916 439508 254944
rect 439508 254893 439564 254902
rect 438946 252992 439406 253020
rect 438850 252881 439022 252909
rect 438994 252710 439022 252881
rect 439378 252710 439406 252992
rect 439714 252724 439742 258635
rect 439714 252696 439776 252724
rect 440098 252710 440126 269439
rect 440482 268435 440510 275502
rect 440566 270533 440618 270539
rect 440566 270475 440618 270481
rect 440468 268426 440524 268435
rect 440468 268361 440524 268370
rect 440578 259217 440606 270475
rect 440662 268165 440714 268171
rect 440662 268107 440714 268113
rect 440674 268023 440702 268107
rect 440662 268017 440714 268023
rect 440662 267959 440714 267965
rect 441634 263403 441662 275502
rect 442882 270507 442910 275502
rect 443540 273754 443596 273763
rect 443540 273689 443596 273698
rect 443554 273499 443582 273689
rect 443542 273493 443594 273499
rect 443542 273435 443594 273441
rect 444034 270655 444062 275502
rect 444020 270646 444076 270655
rect 444020 270581 444076 270590
rect 442868 270498 442924 270507
rect 442868 270433 442924 270442
rect 443446 265057 443498 265063
rect 443446 264999 443498 265005
rect 441620 263394 441676 263403
rect 441620 263329 441676 263338
rect 443254 260173 443306 260179
rect 443254 260115 443306 260121
rect 443158 260025 443210 260031
rect 443158 259967 443210 259973
rect 440566 259211 440618 259217
rect 440566 259153 440618 259159
rect 443170 258773 443198 259967
rect 443266 258847 443294 260115
rect 443254 258841 443306 258847
rect 443254 258783 443306 258789
rect 443062 258767 443114 258773
rect 443062 258709 443114 258715
rect 443158 258767 443210 258773
rect 443158 258709 443210 258715
rect 441526 258249 441578 258255
rect 441526 258191 441578 258197
rect 441238 258175 441290 258181
rect 441238 258117 441290 258123
rect 440854 257139 440906 257145
rect 440854 257081 440906 257087
rect 440470 257065 440522 257071
rect 440470 257007 440522 257013
rect 440278 253217 440330 253223
rect 440278 253159 440330 253165
rect 440290 253043 440318 253159
rect 440276 253034 440332 253043
rect 440276 252969 440332 252978
rect 440482 252710 440510 257007
rect 440758 254993 440810 254999
rect 440758 254935 440810 254941
rect 440662 254771 440714 254777
rect 440662 254713 440714 254719
rect 440674 254523 440702 254713
rect 440660 254514 440716 254523
rect 440660 254449 440716 254458
rect 440770 254375 440798 254935
rect 440756 254366 440812 254375
rect 440756 254301 440812 254310
rect 440866 252710 440894 257081
rect 441250 252724 441278 258117
rect 441538 252872 441566 258191
rect 442678 257213 442730 257219
rect 442678 257155 442730 257161
rect 441910 256991 441962 256997
rect 441910 256933 441962 256939
rect 441538 252844 441614 252872
rect 441216 252696 441278 252724
rect 441586 252710 441614 252844
rect 441922 252724 441950 256933
rect 442294 256621 442346 256627
rect 442294 256563 442346 256569
rect 441922 252696 441984 252724
rect 442306 252710 442334 256563
rect 442690 252710 442718 257155
rect 443074 252710 443102 258709
rect 443458 252724 443486 264999
rect 445282 260327 445310 275502
rect 446434 268985 446462 275502
rect 446422 268979 446474 268985
rect 446422 268921 446474 268927
rect 445270 260321 445322 260327
rect 445270 260263 445322 260269
rect 447682 260253 447710 275502
rect 448834 267695 448862 275502
rect 449986 270655 450014 275502
rect 449972 270646 450028 270655
rect 449972 270581 450028 270590
rect 451138 270507 451166 275502
rect 451124 270498 451180 270507
rect 451124 270433 451180 270442
rect 448820 267686 448876 267695
rect 448820 267621 448876 267630
rect 452386 260475 452414 275502
rect 452662 269275 452714 269281
rect 452662 269217 452714 269223
rect 452374 260469 452426 260475
rect 452374 260411 452426 260417
rect 447670 260247 447722 260253
rect 447670 260189 447722 260195
rect 445654 259211 445706 259217
rect 445654 259153 445706 259159
rect 445270 258545 445322 258551
rect 445270 258487 445322 258493
rect 444502 258471 444554 258477
rect 444502 258413 444554 258419
rect 443734 258323 443786 258329
rect 443734 258265 443786 258271
rect 443542 255733 443594 255739
rect 443638 255733 443690 255739
rect 443594 255681 443638 255684
rect 443542 255675 443690 255681
rect 443554 255656 443678 255675
rect 443638 254919 443690 254925
rect 443638 254861 443690 254867
rect 443542 254845 443594 254851
rect 443542 254787 443594 254793
rect 443554 254523 443582 254787
rect 443540 254514 443596 254523
rect 443540 254449 443596 254458
rect 443650 254375 443678 254861
rect 443636 254366 443692 254375
rect 443636 254301 443692 254310
rect 443746 252872 443774 258265
rect 444118 257509 444170 257515
rect 444118 257451 444170 257457
rect 443746 252844 443822 252872
rect 443424 252696 443486 252724
rect 443794 252710 443822 252844
rect 444130 252724 444158 257451
rect 444310 254327 444362 254333
rect 444310 254269 444362 254275
rect 444322 254079 444350 254269
rect 444308 254070 444364 254079
rect 444308 254005 444364 254014
rect 444130 252696 444192 252724
rect 444514 252710 444542 258413
rect 444886 257435 444938 257441
rect 444886 257377 444938 257383
rect 444898 252710 444926 257377
rect 444980 253330 445036 253339
rect 444980 253265 445036 253274
rect 444994 252927 445022 253265
rect 444982 252921 445034 252927
rect 444982 252863 445034 252869
rect 445282 252710 445310 258487
rect 445366 254401 445418 254407
rect 445366 254343 445418 254349
rect 445378 253487 445406 254343
rect 445364 253478 445420 253487
rect 445364 253413 445420 253422
rect 445364 253034 445420 253043
rect 445364 252969 445366 252978
rect 445418 252969 445420 252978
rect 445366 252937 445418 252943
rect 445666 252724 445694 259153
rect 447862 259137 447914 259143
rect 447862 259079 447914 259085
rect 447958 259137 448010 259143
rect 447958 259079 448010 259085
rect 451894 259137 451946 259143
rect 451894 259079 451946 259085
rect 447094 258619 447146 258625
rect 447094 258561 447146 258567
rect 446710 258397 446762 258403
rect 446710 258339 446762 258345
rect 445942 257731 445994 257737
rect 445942 257673 445994 257679
rect 445954 252872 445982 257673
rect 446326 257657 446378 257663
rect 446326 257599 446378 257605
rect 446228 253034 446284 253043
rect 446228 252969 446284 252978
rect 446242 252927 446270 252969
rect 446230 252921 446282 252927
rect 445954 252844 446030 252872
rect 446230 252863 446282 252869
rect 445632 252696 445694 252724
rect 446002 252710 446030 252844
rect 446338 252724 446366 257599
rect 446422 254475 446474 254481
rect 446422 254417 446474 254423
rect 446434 254375 446462 254417
rect 446420 254366 446476 254375
rect 446420 254301 446476 254310
rect 446422 254253 446474 254259
rect 446420 254218 446422 254227
rect 446474 254218 446476 254227
rect 446420 254153 446476 254162
rect 446422 253143 446474 253149
rect 446422 253085 446474 253091
rect 446434 253043 446462 253085
rect 446420 253034 446476 253043
rect 446420 252969 446476 252978
rect 446338 252696 446400 252724
rect 446722 252710 446750 258339
rect 447106 252710 447134 258561
rect 447476 257770 447532 257779
rect 447476 257705 447532 257714
rect 447490 252710 447518 257705
rect 447874 252724 447902 259079
rect 447970 258995 447998 259079
rect 449398 259063 449450 259069
rect 449398 259005 449450 259011
rect 447958 258989 448010 258995
rect 447958 258931 448010 258937
rect 448148 257918 448204 257927
rect 448148 257853 448204 257862
rect 448162 253020 448190 257853
rect 448918 257805 448970 257811
rect 448918 257747 448970 257753
rect 448534 257583 448586 257589
rect 448534 257525 448586 257531
rect 448162 252992 448238 253020
rect 447840 252696 447902 252724
rect 448210 252710 448238 252992
rect 448546 252724 448574 257525
rect 448546 252696 448608 252724
rect 448930 252710 448958 257747
rect 449410 252872 449438 259005
rect 451126 258767 451178 258773
rect 451126 258709 451178 258715
rect 450358 258027 450410 258033
rect 450358 257969 450410 257975
rect 449590 257879 449642 257885
rect 449590 257821 449642 257827
rect 449602 254056 449630 257821
rect 450070 256473 450122 256479
rect 450070 256415 450122 256421
rect 449602 254028 449726 254056
rect 449314 252844 449438 252872
rect 449314 252710 449342 252844
rect 449698 252710 449726 254028
rect 450082 252724 450110 256415
rect 450370 252872 450398 257969
rect 450742 256399 450794 256405
rect 450742 256341 450794 256347
rect 450370 252844 450446 252872
rect 450048 252696 450110 252724
rect 450418 252710 450446 252844
rect 450754 252724 450782 256341
rect 450754 252696 450816 252724
rect 451138 252710 451166 258709
rect 451510 256547 451562 256553
rect 451510 256489 451562 256495
rect 451522 252710 451550 256489
rect 451906 252710 451934 259079
rect 452278 256769 452330 256775
rect 452278 256711 452330 256717
rect 452290 252724 452318 256711
rect 452674 253020 452702 269217
rect 453538 262843 453566 275502
rect 454690 267653 454718 275502
rect 454678 267647 454730 267653
rect 454678 267589 454730 267595
rect 455938 264883 455966 275502
rect 456802 275488 457104 275516
rect 457954 275488 458352 275516
rect 455924 264874 455980 264883
rect 455924 264809 455980 264818
rect 453526 262837 453578 262843
rect 453526 262779 453578 262785
rect 452950 258989 453002 258995
rect 452950 258931 453002 258937
rect 452256 252696 452318 252724
rect 452626 252992 452702 253020
rect 452626 252710 452654 252992
rect 452962 252724 452990 258931
rect 456802 257811 456830 275488
rect 455446 257805 455498 257811
rect 455446 257747 455498 257753
rect 456790 257805 456842 257811
rect 456790 257747 456842 257753
rect 452962 252696 453024 252724
rect 288598 239675 288650 239681
rect 288598 239617 288650 239623
rect 288406 239231 288458 239237
rect 288406 239173 288458 239179
rect 288310 237899 288362 237905
rect 288310 237841 288362 237847
rect 287926 237751 287978 237757
rect 287926 237693 287978 237699
rect 287830 236567 287882 236573
rect 287830 236509 287882 236515
rect 287542 236419 287594 236425
rect 287542 236361 287594 236367
rect 287446 236271 287498 236277
rect 287446 236213 287498 236219
rect 287158 236197 287210 236203
rect 287158 236139 287210 236145
rect 286966 231091 287018 231097
rect 286966 231033 287018 231039
rect 288706 229025 288734 239834
rect 289042 239700 289070 239834
rect 288994 239672 289070 239700
rect 288994 239575 289022 239672
rect 289426 239607 289454 239834
rect 289414 239601 289466 239607
rect 288980 239566 289036 239575
rect 289762 239575 289790 239834
rect 289414 239543 289466 239549
rect 289748 239566 289804 239575
rect 288980 239501 289036 239510
rect 289748 239501 289804 239510
rect 289556 239418 289612 239427
rect 289556 239353 289612 239362
rect 289570 238793 289598 239353
rect 289558 238787 289610 238793
rect 289558 238729 289610 238735
rect 290146 236055 290174 239834
rect 290530 239681 290558 239834
rect 290518 239675 290570 239681
rect 290518 239617 290570 239623
rect 290914 239575 290942 239834
rect 291250 239700 291278 239834
rect 291634 239700 291662 239834
rect 291250 239672 291422 239700
rect 291394 239575 291422 239672
rect 291586 239672 291662 239700
rect 291586 239575 291614 239672
rect 291970 239575 291998 239834
rect 292354 239575 292382 239834
rect 292738 239575 292766 239834
rect 293122 239575 293150 239834
rect 293458 239700 293486 239834
rect 293842 239700 293870 239834
rect 293410 239672 293486 239700
rect 293794 239672 293870 239700
rect 290900 239566 290956 239575
rect 290900 239501 290956 239510
rect 291188 239566 291244 239575
rect 291188 239501 291190 239510
rect 291242 239501 291244 239510
rect 291380 239566 291436 239575
rect 291380 239501 291436 239510
rect 291572 239566 291628 239575
rect 291572 239501 291628 239510
rect 291956 239566 292012 239575
rect 291956 239501 292012 239510
rect 292340 239566 292396 239575
rect 292340 239501 292396 239510
rect 292724 239566 292780 239575
rect 292724 239501 292780 239510
rect 293108 239566 293164 239575
rect 293108 239501 293164 239510
rect 291190 239469 291242 239475
rect 293410 239427 293438 239672
rect 293108 239418 293164 239427
rect 293108 239353 293164 239362
rect 293396 239418 293452 239427
rect 293396 239353 293452 239362
rect 293122 239311 293150 239353
rect 293110 239305 293162 239311
rect 293110 239247 293162 239253
rect 293794 239131 293822 239672
rect 293780 239122 293836 239131
rect 293780 239057 293836 239066
rect 290134 236049 290186 236055
rect 290134 235991 290186 235997
rect 294178 235981 294206 239834
rect 294562 236023 294590 239834
rect 294946 239575 294974 239834
rect 294932 239566 294988 239575
rect 294932 239501 294988 239510
rect 295330 236171 295358 239834
rect 295666 239700 295694 239834
rect 296050 239700 296078 239834
rect 295618 239672 295694 239700
rect 296002 239672 296078 239700
rect 295316 236162 295372 236171
rect 295316 236097 295372 236106
rect 294548 236014 294604 236023
rect 294166 235975 294218 235981
rect 294548 235949 294604 235958
rect 294166 235917 294218 235923
rect 295618 235875 295646 239672
rect 296002 238983 296030 239672
rect 295988 238974 296044 238983
rect 295988 238909 296044 238918
rect 295604 235866 295660 235875
rect 295604 235801 295660 235810
rect 296386 235579 296414 239834
rect 296564 236458 296620 236467
rect 296564 236393 296620 236402
rect 296578 236351 296606 236393
rect 296566 236345 296618 236351
rect 296566 236287 296618 236293
rect 296770 235727 296798 239834
rect 296756 235718 296812 235727
rect 296756 235653 296812 235662
rect 296372 235570 296428 235579
rect 296372 235505 296428 235514
rect 297154 235135 297182 239834
rect 297538 235875 297566 239834
rect 297874 239700 297902 239834
rect 297826 239672 297902 239700
rect 297826 239279 297854 239672
rect 298258 239552 298286 239834
rect 298210 239524 298286 239552
rect 297812 239270 297868 239279
rect 297812 239205 297868 239214
rect 298004 238974 298060 238983
rect 298004 238909 298060 238918
rect 298018 238687 298046 238909
rect 298004 238678 298060 238687
rect 298004 238613 298060 238622
rect 298210 236129 298238 239524
rect 298198 236123 298250 236129
rect 298198 236065 298250 236071
rect 297524 235866 297580 235875
rect 297524 235801 297580 235810
rect 298594 235431 298622 239834
rect 298978 236467 299006 239834
rect 298964 236458 299020 236467
rect 298964 236393 299020 236402
rect 299362 236319 299390 239834
rect 299746 236615 299774 239834
rect 300082 239552 300110 239834
rect 300466 239552 300494 239834
rect 300082 239524 300158 239552
rect 300466 239524 300542 239552
rect 300130 236763 300158 239524
rect 300514 237207 300542 239524
rect 300500 237198 300556 237207
rect 300500 237133 300556 237142
rect 300802 236911 300830 239834
rect 301186 237503 301214 239834
rect 301570 237947 301598 239834
rect 301556 237938 301612 237947
rect 301556 237873 301612 237882
rect 301172 237494 301228 237503
rect 301172 237429 301228 237438
rect 301954 237059 301982 239834
rect 302290 239552 302318 239834
rect 302242 239524 302318 239552
rect 302674 239552 302702 239834
rect 302674 239524 302750 239552
rect 301940 237050 301996 237059
rect 301940 236985 301996 236994
rect 300788 236902 300844 236911
rect 300788 236837 300844 236846
rect 300116 236754 300172 236763
rect 300116 236689 300172 236698
rect 299732 236606 299788 236615
rect 299732 236541 299788 236550
rect 299348 236310 299404 236319
rect 299348 236245 299404 236254
rect 302242 235759 302270 239524
rect 302230 235753 302282 235759
rect 302230 235695 302282 235701
rect 298580 235422 298636 235431
rect 298580 235357 298636 235366
rect 297140 235126 297196 235135
rect 297140 235061 297196 235070
rect 302722 234247 302750 239524
rect 302708 234238 302764 234247
rect 302708 234173 302764 234182
rect 303010 233507 303038 239834
rect 302996 233498 303052 233507
rect 302996 233433 303052 233442
rect 288694 229019 288746 229025
rect 288694 228961 288746 228967
rect 286486 228797 286538 228803
rect 286486 228739 286538 228745
rect 285622 228723 285674 228729
rect 285622 228665 285674 228671
rect 284278 228353 284330 228359
rect 284278 228295 284330 228301
rect 283798 228131 283850 228137
rect 283798 228073 283850 228079
rect 242038 227761 242090 227767
rect 241954 227721 242038 227749
rect 221878 227613 221930 227619
rect 221878 227555 221930 227561
rect 221782 227539 221834 227545
rect 221782 227481 221834 227487
rect 221794 227416 221822 227481
rect 221890 227416 221918 227555
rect 221794 227388 221918 227416
rect 215746 223836 215822 223864
rect 215794 223554 215822 223836
rect 241954 223554 241982 227721
rect 242038 227703 242090 227709
rect 293398 227687 293450 227693
rect 293398 227629 293450 227635
rect 242038 227613 242090 227619
rect 242038 227555 242090 227561
rect 242050 227397 242078 227555
rect 242038 227391 242090 227397
rect 242038 227333 242090 227339
rect 293410 223864 293438 227629
rect 303394 227143 303422 239834
rect 303778 227439 303806 239834
rect 303764 227430 303820 227439
rect 303764 227365 303820 227374
rect 303380 227134 303436 227143
rect 303380 227069 303436 227078
rect 304162 226287 304190 239834
rect 304498 239552 304526 239834
rect 304882 239552 304910 239834
rect 304498 239524 304574 239552
rect 304882 239524 304958 239552
rect 304546 226995 304574 239524
rect 304532 226986 304588 226995
rect 304532 226921 304588 226930
rect 304150 226281 304202 226287
rect 304150 226223 304202 226229
rect 304930 226139 304958 239524
rect 305108 238234 305164 238243
rect 305108 238169 305164 238178
rect 305122 238053 305150 238169
rect 305110 238047 305162 238053
rect 305110 237989 305162 237995
rect 305218 227291 305246 239834
rect 305204 227282 305260 227291
rect 305204 227217 305260 227226
rect 305602 226435 305630 239834
rect 305590 226429 305642 226435
rect 305590 226371 305642 226377
rect 304918 226133 304970 226139
rect 305986 226107 306014 239834
rect 306370 226213 306398 239834
rect 306706 239552 306734 239834
rect 307090 239552 307118 239834
rect 306706 239524 306782 239552
rect 307090 239524 307166 239552
rect 306754 226699 306782 239524
rect 306740 226690 306796 226699
rect 306740 226625 306796 226634
rect 307138 226583 307166 239524
rect 307426 226847 307454 239834
rect 307412 226838 307468 226847
rect 307412 226773 307468 226782
rect 307126 226577 307178 226583
rect 307126 226519 307178 226525
rect 307810 226361 307838 239834
rect 307798 226355 307850 226361
rect 307798 226297 307850 226303
rect 308194 226255 308222 239834
rect 308578 233539 308606 239834
rect 308914 239552 308942 239834
rect 309298 239552 309326 239834
rect 308914 239524 308990 239552
rect 309298 239524 309374 239552
rect 308962 233687 308990 239524
rect 309346 235389 309374 239524
rect 309334 235383 309386 235389
rect 309334 235325 309386 235331
rect 309634 234691 309662 239834
rect 310018 234871 310046 239834
rect 310006 234865 310058 234871
rect 310402 234839 310430 239834
rect 310006 234807 310058 234813
rect 310388 234830 310444 234839
rect 310388 234765 310444 234774
rect 309620 234682 309676 234691
rect 309620 234617 309676 234626
rect 310786 234353 310814 239834
rect 311122 239552 311150 239834
rect 311506 239552 311534 239834
rect 311122 239524 311198 239552
rect 311506 239524 311582 239552
rect 311170 235093 311198 239524
rect 311554 235463 311582 239524
rect 311542 235457 311594 235463
rect 311542 235399 311594 235405
rect 311158 235087 311210 235093
rect 311158 235029 311210 235035
rect 311842 234501 311870 239834
rect 311830 234495 311882 234501
rect 311830 234437 311882 234443
rect 312226 234427 312254 239834
rect 312610 235135 312638 239834
rect 312994 235537 313022 239834
rect 313330 239552 313358 239834
rect 313714 239552 313742 239834
rect 313330 239524 313406 239552
rect 313714 239524 313790 239552
rect 312982 235531 313034 235537
rect 312982 235473 313034 235479
rect 313378 235283 313406 239524
rect 313364 235274 313420 235283
rect 313364 235209 313420 235218
rect 312596 235126 312652 235135
rect 312596 235061 312652 235070
rect 312214 234421 312266 234427
rect 312214 234363 312266 234369
rect 310774 234347 310826 234353
rect 310774 234289 310826 234295
rect 313762 234131 313790 239524
rect 314050 235167 314078 239834
rect 314038 235161 314090 235167
rect 314038 235103 314090 235109
rect 313750 234125 313802 234131
rect 313750 234067 313802 234073
rect 314434 234057 314462 239834
rect 314818 235727 314846 239834
rect 314804 235718 314860 235727
rect 314804 235653 314860 235662
rect 314422 234051 314474 234057
rect 314422 233993 314474 233999
rect 308950 233681 309002 233687
rect 308950 233623 309002 233629
rect 308566 233533 308618 233539
rect 308566 233475 308618 233481
rect 315202 227027 315230 239834
rect 315538 239552 315566 239834
rect 315922 239552 315950 239834
rect 315538 239524 315614 239552
rect 315922 239524 315998 239552
rect 315586 235431 315614 239524
rect 315572 235422 315628 235431
rect 315572 235357 315628 235366
rect 315970 227175 315998 239524
rect 316258 235579 316286 239834
rect 316244 235570 316300 235579
rect 316244 235505 316300 235514
rect 315958 227169 316010 227175
rect 315958 227111 316010 227117
rect 316642 227101 316670 239834
rect 317026 235241 317054 239834
rect 317014 235235 317066 235241
rect 317014 235177 317066 235183
rect 317410 234723 317438 239834
rect 317746 239552 317774 239834
rect 318130 239552 318158 239834
rect 317746 239524 317822 239552
rect 318130 239524 318206 239552
rect 317398 234717 317450 234723
rect 317398 234659 317450 234665
rect 316630 227095 316682 227101
rect 316630 227037 316682 227043
rect 315190 227021 315242 227027
rect 315190 226963 315242 226969
rect 317794 226731 317822 239524
rect 318178 234797 318206 239524
rect 318166 234791 318218 234797
rect 318166 234733 318218 234739
rect 317782 226725 317834 226731
rect 317782 226667 317834 226673
rect 318466 226657 318494 239834
rect 318850 235019 318878 239834
rect 318838 235013 318890 235019
rect 318838 234955 318890 234961
rect 318838 229019 318890 229025
rect 318838 228961 318890 228967
rect 318454 226651 318506 226657
rect 318454 226593 318506 226599
rect 308180 226246 308236 226255
rect 306358 226207 306410 226213
rect 308180 226181 308236 226190
rect 306358 226149 306410 226155
rect 304918 226075 304970 226081
rect 305972 226098 306028 226107
rect 305972 226033 306028 226042
rect 293410 223836 293486 223864
rect 293458 223554 293486 223836
rect 318850 223554 318878 228961
rect 319234 226509 319262 239834
rect 319618 233909 319646 239834
rect 319954 239552 319982 239834
rect 320338 239552 320366 239834
rect 319954 239524 320030 239552
rect 320338 239524 320414 239552
rect 319606 233903 319658 233909
rect 319606 233845 319658 233851
rect 320002 233835 320030 239524
rect 320386 234279 320414 239524
rect 320374 234273 320426 234279
rect 320374 234215 320426 234221
rect 319990 233829 320042 233835
rect 319990 233771 320042 233777
rect 320674 233761 320702 239834
rect 321058 234945 321086 239834
rect 321046 234939 321098 234945
rect 321046 234881 321098 234887
rect 320662 233755 320714 233761
rect 320662 233697 320714 233703
rect 321442 233613 321470 239834
rect 321430 233607 321482 233613
rect 321430 233549 321482 233555
rect 321826 232725 321854 239834
rect 322162 239552 322190 239834
rect 322546 239700 322574 239834
rect 322498 239672 322574 239700
rect 322162 239524 322238 239552
rect 322210 233983 322238 239524
rect 322198 233977 322250 233983
rect 322198 233919 322250 233925
rect 321814 232719 321866 232725
rect 321814 232661 321866 232667
rect 322498 231911 322526 239672
rect 322882 233465 322910 239834
rect 322870 233459 322922 233465
rect 322870 233401 322922 233407
rect 323266 232059 323294 239834
rect 323650 234205 323678 239834
rect 323638 234199 323690 234205
rect 323638 234141 323690 234147
rect 324034 232133 324062 239834
rect 324370 239552 324398 239834
rect 324754 239552 324782 239834
rect 324370 239524 324446 239552
rect 324754 239524 324830 239552
rect 324418 236055 324446 239524
rect 324406 236049 324458 236055
rect 324406 235991 324458 235997
rect 324802 232207 324830 239524
rect 325090 235981 325118 239834
rect 325474 239089 325502 239834
rect 325462 239083 325514 239089
rect 325462 239025 325514 239031
rect 325558 237899 325610 237905
rect 325558 237841 325610 237847
rect 325570 237799 325598 237841
rect 325556 237790 325612 237799
rect 325556 237725 325612 237734
rect 325078 235975 325130 235981
rect 325078 235917 325130 235923
rect 324790 232201 324842 232207
rect 324790 232143 324842 232149
rect 324022 232127 324074 232133
rect 324022 232069 324074 232075
rect 323254 232053 323306 232059
rect 323254 231995 323306 232001
rect 322486 231905 322538 231911
rect 322486 231847 322538 231853
rect 319222 226503 319274 226509
rect 319222 226445 319274 226451
rect 325858 224215 325886 239834
rect 325942 237899 325994 237905
rect 325942 237841 325994 237847
rect 325954 237799 325982 237841
rect 325940 237790 325996 237799
rect 325940 237725 325996 237734
rect 326242 232577 326270 239834
rect 326578 239552 326606 239834
rect 326962 239552 326990 239834
rect 326578 239524 326654 239552
rect 326962 239524 327038 239552
rect 326230 232571 326282 232577
rect 326230 232513 326282 232519
rect 326626 226879 326654 239524
rect 326902 233681 326954 233687
rect 326902 233623 326954 233629
rect 326806 233533 326858 233539
rect 326806 233475 326858 233481
rect 326818 227249 326846 233475
rect 326806 227243 326858 227249
rect 326806 227185 326858 227191
rect 326614 226873 326666 226879
rect 326614 226815 326666 226821
rect 326914 226403 326942 233623
rect 327010 232651 327038 239524
rect 327298 236129 327326 239834
rect 327286 236123 327338 236129
rect 327286 236065 327338 236071
rect 327190 234125 327242 234131
rect 327190 234067 327242 234073
rect 327094 234051 327146 234057
rect 327094 233993 327146 233999
rect 327106 233761 327134 233993
rect 327094 233755 327146 233761
rect 327094 233697 327146 233703
rect 327202 233687 327230 234067
rect 327190 233681 327242 233687
rect 327190 233623 327242 233629
rect 326998 232645 327050 232651
rect 326998 232587 327050 232593
rect 327682 232503 327710 239834
rect 327670 232497 327722 232503
rect 327670 232439 327722 232445
rect 326900 226394 326956 226403
rect 326900 226329 326956 226338
rect 325846 224209 325898 224215
rect 325846 224151 325898 224157
rect 328066 224067 328094 239834
rect 328450 235315 328478 239834
rect 328786 239552 328814 239834
rect 329170 239552 329198 239834
rect 328786 239524 328862 239552
rect 329170 239524 329246 239552
rect 328438 235309 328490 235315
rect 328438 235251 328490 235257
rect 328726 234125 328778 234131
rect 328726 234067 328778 234073
rect 328738 233687 328766 234067
rect 328834 233687 328862 239524
rect 328726 233681 328778 233687
rect 328726 233623 328778 233629
rect 328822 233681 328874 233687
rect 328822 233623 328874 233629
rect 329218 227471 329246 239524
rect 329506 234501 329534 239834
rect 329890 234649 329918 239834
rect 329878 234643 329930 234649
rect 329878 234585 329930 234591
rect 329494 234495 329546 234501
rect 329494 234437 329546 234443
rect 329206 227465 329258 227471
rect 329206 227407 329258 227413
rect 328054 224061 328106 224067
rect 328054 224003 328106 224009
rect 330274 223845 330302 239834
rect 330454 233681 330506 233687
rect 330454 233623 330506 233629
rect 330466 223919 330494 233623
rect 330658 232471 330686 239834
rect 330994 239552 331022 239834
rect 331378 239552 331406 239834
rect 330994 239524 331070 239552
rect 331378 239524 331454 239552
rect 331042 232767 331070 239524
rect 331426 237609 331454 239524
rect 331414 237603 331466 237609
rect 331414 237545 331466 237551
rect 331028 232758 331084 232767
rect 331028 232693 331084 232702
rect 330644 232462 330700 232471
rect 330644 232397 330700 232406
rect 331714 232323 331742 239834
rect 332098 237461 332126 239834
rect 332086 237455 332138 237461
rect 332086 237397 332138 237403
rect 332482 237387 332510 239834
rect 332470 237381 332522 237387
rect 332470 237323 332522 237329
rect 332866 232915 332894 239834
rect 333202 239552 333230 239834
rect 333586 239552 333614 239834
rect 333202 239524 333278 239552
rect 333586 239524 333662 239552
rect 333250 237165 333278 239524
rect 333238 237159 333290 237165
rect 333238 237101 333290 237107
rect 332852 232906 332908 232915
rect 332852 232841 332908 232850
rect 331700 232314 331756 232323
rect 331700 232249 331756 232258
rect 333634 231837 333662 239524
rect 333622 231831 333674 231837
rect 333622 231773 333674 231779
rect 333922 226953 333950 239834
rect 334306 235759 334334 239834
rect 334690 237535 334718 239834
rect 334678 237529 334730 237535
rect 334678 237471 334730 237477
rect 334294 235753 334346 235759
rect 334294 235695 334346 235701
rect 335074 231985 335102 239834
rect 335410 239552 335438 239834
rect 335794 239552 335822 239834
rect 335410 239524 335486 239552
rect 335794 239524 335870 239552
rect 335458 237313 335486 239524
rect 335446 237307 335498 237313
rect 335446 237249 335498 237255
rect 335842 232281 335870 239524
rect 336130 237239 336158 239834
rect 336118 237233 336170 237239
rect 336118 237175 336170 237181
rect 336514 232947 336542 239834
rect 336502 232941 336554 232947
rect 336502 232883 336554 232889
rect 335830 232275 335882 232281
rect 335830 232217 335882 232223
rect 335062 231979 335114 231985
rect 335062 231921 335114 231927
rect 336898 231615 336926 239834
rect 337282 238645 337310 239834
rect 337618 239552 337646 239834
rect 338002 239552 338030 239834
rect 337618 239524 337694 239552
rect 337174 238639 337226 238645
rect 337174 238581 337226 238587
rect 337270 238639 337322 238645
rect 337270 238581 337322 238587
rect 337186 238127 337214 238581
rect 337174 238121 337226 238127
rect 337174 238063 337226 238069
rect 337666 232355 337694 239524
rect 337954 239524 338030 239552
rect 337654 232349 337706 232355
rect 337654 232291 337706 232297
rect 336886 231609 336938 231615
rect 336886 231551 336938 231557
rect 337954 231435 337982 239524
rect 338338 236740 338366 239834
rect 338518 237603 338570 237609
rect 338518 237545 338570 237551
rect 338050 236712 338366 236740
rect 337940 231426 337996 231435
rect 337940 231361 337996 231370
rect 338050 231319 338078 236712
rect 338242 236573 338462 236592
rect 338242 236567 338474 236573
rect 338242 236564 338422 236567
rect 338242 236425 338270 236564
rect 338422 236509 338474 236515
rect 338230 236419 338282 236425
rect 338230 236361 338282 236367
rect 338326 236419 338378 236425
rect 338326 236361 338378 236367
rect 338338 236277 338366 236361
rect 338326 236271 338378 236277
rect 338326 236213 338378 236219
rect 338230 236049 338282 236055
rect 338230 235991 338282 235997
rect 338326 236049 338378 236055
rect 338530 236023 338558 237545
rect 338326 235991 338378 235997
rect 338516 236014 338572 236023
rect 338242 235611 338270 235991
rect 338230 235605 338282 235611
rect 338230 235547 338282 235553
rect 338338 235537 338366 235991
rect 338516 235949 338572 235958
rect 338722 235704 338750 239834
rect 339106 238275 339134 239834
rect 339490 238719 339518 239834
rect 339826 239552 339854 239834
rect 340210 239552 340238 239834
rect 339826 239524 339902 239552
rect 339478 238713 339530 238719
rect 339478 238655 339530 238661
rect 339874 238497 339902 239524
rect 340162 239524 340238 239552
rect 340162 238867 340190 239524
rect 340150 238861 340202 238867
rect 340150 238803 340202 238809
rect 340546 238571 340574 239834
rect 340534 238565 340586 238571
rect 340534 238507 340586 238513
rect 339862 238491 339914 238497
rect 339862 238433 339914 238439
rect 340930 238423 340958 239834
rect 340918 238417 340970 238423
rect 340918 238359 340970 238365
rect 341014 238417 341066 238423
rect 341014 238359 341066 238365
rect 339094 238269 339146 238275
rect 339094 238211 339146 238217
rect 341026 236795 341054 238359
rect 341110 238121 341162 238127
rect 341110 238063 341162 238069
rect 341122 236795 341150 238063
rect 341014 236789 341066 236795
rect 341014 236731 341066 236737
rect 341110 236789 341162 236795
rect 341110 236731 341162 236737
rect 338722 235676 338846 235704
rect 338710 235605 338762 235611
rect 338710 235547 338762 235553
rect 338326 235531 338378 235537
rect 338326 235473 338378 235479
rect 338614 235457 338666 235463
rect 338614 235399 338666 235405
rect 338134 235309 338186 235315
rect 338518 235309 338570 235315
rect 338186 235257 338462 235260
rect 338134 235251 338462 235257
rect 338518 235251 338570 235257
rect 338146 235232 338462 235251
rect 338434 235167 338462 235232
rect 338326 235161 338378 235167
rect 338326 235103 338378 235109
rect 338422 235161 338474 235167
rect 338422 235103 338474 235109
rect 338338 234871 338366 235103
rect 338230 234865 338282 234871
rect 338230 234807 338282 234813
rect 338326 234865 338378 234871
rect 338530 234816 338558 235251
rect 338326 234807 338378 234813
rect 338242 234668 338270 234807
rect 338434 234788 338558 234816
rect 338434 234668 338462 234788
rect 338242 234640 338462 234668
rect 338626 234205 338654 235399
rect 338518 234199 338570 234205
rect 338518 234141 338570 234147
rect 338614 234199 338666 234205
rect 338614 234141 338666 234147
rect 338326 234051 338378 234057
rect 338326 233993 338378 233999
rect 338338 233539 338366 233993
rect 338422 233977 338474 233983
rect 338422 233919 338474 233925
rect 338434 233761 338462 233919
rect 338422 233755 338474 233761
rect 338422 233697 338474 233703
rect 338530 233539 338558 234141
rect 338722 233983 338750 235547
rect 338818 235463 338846 235676
rect 338998 235605 339050 235611
rect 338998 235547 339050 235553
rect 338806 235457 338858 235463
rect 338806 235399 338858 235405
rect 339010 234501 339038 235547
rect 341314 234987 341342 239834
rect 341590 239083 341642 239089
rect 341590 239025 341642 239031
rect 341300 234978 341356 234987
rect 341300 234913 341356 234922
rect 338998 234495 339050 234501
rect 338998 234437 339050 234443
rect 338710 233977 338762 233983
rect 338710 233919 338762 233925
rect 338326 233533 338378 233539
rect 338326 233475 338378 233481
rect 338518 233533 338570 233539
rect 338518 233475 338570 233481
rect 341602 232429 341630 239025
rect 341698 238983 341726 239834
rect 342034 239552 342062 239834
rect 342418 239552 342446 239834
rect 342034 239524 342110 239552
rect 342418 239524 342494 239552
rect 341684 238974 341740 238983
rect 341684 238909 341740 238918
rect 341590 232423 341642 232429
rect 341590 232365 341642 232371
rect 338038 231313 338090 231319
rect 338038 231255 338090 231261
rect 342082 230843 342110 239524
rect 342466 238687 342494 239524
rect 342754 239108 342782 239834
rect 342754 239080 342878 239108
rect 342742 239009 342794 239015
rect 342742 238951 342794 238957
rect 342754 238867 342782 238951
rect 342742 238861 342794 238867
rect 342742 238803 342794 238809
rect 342452 238678 342508 238687
rect 342452 238613 342508 238622
rect 342740 235866 342796 235875
rect 342740 235801 342796 235810
rect 342754 234501 342782 235801
rect 342742 234495 342794 234501
rect 342742 234437 342794 234443
rect 342850 230991 342878 239080
rect 343138 232619 343166 239834
rect 343124 232610 343180 232619
rect 343124 232545 343180 232554
rect 342836 230982 342892 230991
rect 342836 230917 342892 230926
rect 342068 230834 342124 230843
rect 342068 230769 342124 230778
rect 333910 226947 333962 226953
rect 333910 226889 333962 226895
rect 343522 224331 343550 239834
rect 343906 237799 343934 239834
rect 344242 239552 344270 239834
rect 344626 239552 344654 239834
rect 344242 239524 344318 239552
rect 344626 239524 344702 239552
rect 344290 239015 344318 239524
rect 344278 239009 344330 239015
rect 344278 238951 344330 238957
rect 344674 238127 344702 239524
rect 344962 238275 344990 239834
rect 345346 238867 345374 239834
rect 345334 238861 345386 238867
rect 345334 238803 345386 238809
rect 345730 238497 345758 239834
rect 345814 239083 345866 239089
rect 345814 239025 345866 239031
rect 345718 238491 345770 238497
rect 345718 238433 345770 238439
rect 344950 238269 345002 238275
rect 344950 238211 345002 238217
rect 345620 238234 345676 238243
rect 345620 238169 345622 238178
rect 345674 238169 345676 238178
rect 345622 238137 345674 238143
rect 344662 238121 344714 238127
rect 344662 238063 344714 238069
rect 345526 238047 345578 238053
rect 345826 238035 345854 239025
rect 346114 238571 346142 239834
rect 346450 239552 346478 239834
rect 346834 239552 346862 239834
rect 346450 239524 346526 239552
rect 346834 239524 346910 239552
rect 346498 238719 346526 239524
rect 346882 238867 346910 239524
rect 346870 238861 346922 238867
rect 346870 238803 346922 238809
rect 346486 238713 346538 238719
rect 346486 238655 346538 238661
rect 346102 238565 346154 238571
rect 346102 238507 346154 238513
rect 345908 238234 345964 238243
rect 345908 238169 345964 238178
rect 345578 238007 345854 238035
rect 345526 237989 345578 237995
rect 343892 237790 343948 237799
rect 343892 237725 343948 237734
rect 345622 236271 345674 236277
rect 345622 236213 345674 236219
rect 344470 235161 344522 235167
rect 344470 235103 344522 235109
rect 344482 234649 344510 235103
rect 344470 234643 344522 234649
rect 344470 234585 344522 234591
rect 344278 234569 344330 234575
rect 344278 234511 344330 234517
rect 343796 227726 343852 227735
rect 343796 227661 343852 227670
rect 343508 224322 343564 224331
rect 343508 224257 343564 224266
rect 338326 224209 338378 224215
rect 338326 224151 338378 224157
rect 330454 223913 330506 223919
rect 330454 223855 330506 223861
rect 338338 223845 338366 224151
rect 343810 223864 343838 227661
rect 344290 227323 344318 234511
rect 345634 231023 345662 236213
rect 345622 231017 345674 231023
rect 345622 230959 345674 230965
rect 345922 230875 345950 238169
rect 347170 238095 347198 239834
rect 347554 238243 347582 239834
rect 347540 238234 347596 238243
rect 347540 238169 347596 238178
rect 347156 238086 347212 238095
rect 347156 238021 347212 238030
rect 346774 235605 346826 235611
rect 346774 235547 346826 235553
rect 346786 234131 346814 235547
rect 346678 234125 346730 234131
rect 346678 234067 346730 234073
rect 346774 234125 346826 234131
rect 346774 234067 346826 234073
rect 345910 230869 345962 230875
rect 345910 230811 345962 230817
rect 346486 229019 346538 229025
rect 346486 228961 346538 228967
rect 346102 228427 346154 228433
rect 346102 228369 346154 228375
rect 344948 228318 345004 228327
rect 344948 228253 345004 228262
rect 344278 227317 344330 227323
rect 344278 227259 344330 227265
rect 330262 223839 330314 223845
rect 330262 223781 330314 223787
rect 338326 223839 338378 223845
rect 343810 223836 343886 223864
rect 338326 223781 338378 223787
rect 343858 223554 343886 223836
rect 344962 223554 344990 228253
rect 345332 228170 345388 228179
rect 345332 228105 345388 228114
rect 345346 223554 345374 228105
rect 345716 227578 345772 227587
rect 345716 227513 345772 227522
rect 345730 223554 345758 227513
rect 346114 223864 346142 228369
rect 346498 223864 346526 228961
rect 346690 227397 346718 234067
rect 347938 233669 347966 239834
rect 348322 233669 348350 239834
rect 348658 239552 348686 239834
rect 349042 239552 349070 239834
rect 348658 239524 348734 239552
rect 349042 239524 349118 239552
rect 348502 233681 348554 233687
rect 347938 233641 348062 233669
rect 348322 233641 348446 233669
rect 347926 229611 347978 229617
rect 347926 229553 347978 229559
rect 347158 229389 347210 229395
rect 347158 229331 347210 229337
rect 346774 228353 346826 228359
rect 346774 228295 346826 228301
rect 346678 227391 346730 227397
rect 346678 227333 346730 227339
rect 346066 223836 346142 223864
rect 346450 223836 346526 223864
rect 346066 223554 346094 223836
rect 346450 223554 346478 223836
rect 346786 223554 346814 228295
rect 347170 223554 347198 229331
rect 347542 229315 347594 229321
rect 347542 229257 347594 229263
rect 347554 223554 347582 229257
rect 347938 223554 347966 229553
rect 348034 224627 348062 233641
rect 348310 229685 348362 229691
rect 348310 229627 348362 229633
rect 348214 227465 348266 227471
rect 348214 227407 348266 227413
rect 348226 226805 348254 227407
rect 348214 226799 348266 226805
rect 348214 226741 348266 226747
rect 348020 224618 348076 224627
rect 348020 224553 348076 224562
rect 348322 223864 348350 229627
rect 348418 226551 348446 233641
rect 348502 233623 348554 233629
rect 348514 227471 348542 233623
rect 348598 233459 348650 233465
rect 348598 233401 348650 233407
rect 348502 227465 348554 227471
rect 348502 227407 348554 227413
rect 348404 226542 348460 226551
rect 348404 226477 348460 226486
rect 348610 224067 348638 233401
rect 348706 232873 348734 239524
rect 348886 236049 348938 236055
rect 348886 235991 348938 235997
rect 348788 234830 348844 234839
rect 348788 234765 348844 234774
rect 348694 232867 348746 232873
rect 348694 232809 348746 232815
rect 348694 229759 348746 229765
rect 348694 229701 348746 229707
rect 348598 224061 348650 224067
rect 348598 224003 348650 224009
rect 348706 223864 348734 229701
rect 348802 225959 348830 234765
rect 348788 225950 348844 225959
rect 348788 225885 348844 225894
rect 348898 224733 348926 235991
rect 349090 233021 349118 239524
rect 349378 238941 349406 239834
rect 349366 238935 349418 238941
rect 349366 238877 349418 238883
rect 349174 233977 349226 233983
rect 349174 233919 349226 233925
rect 349078 233015 349130 233021
rect 349078 232957 349130 232963
rect 348982 229833 349034 229839
rect 348982 229775 349034 229781
rect 348886 224727 348938 224733
rect 348886 224669 348938 224675
rect 348274 223836 348350 223864
rect 348658 223836 348734 223864
rect 348274 223554 348302 223836
rect 348658 223554 348686 223836
rect 348994 223554 349022 229775
rect 349186 223887 349214 233919
rect 349762 231245 349790 239834
rect 350146 237683 350174 239834
rect 350134 237677 350186 237683
rect 350134 237619 350186 237625
rect 349750 231239 349802 231245
rect 349750 231181 349802 231187
rect 350134 229981 350186 229987
rect 350134 229923 350186 229929
rect 349750 229907 349802 229913
rect 349750 229849 349802 229855
rect 349366 228649 349418 228655
rect 349366 228591 349418 228597
rect 349172 223878 349228 223887
rect 349172 223813 349228 223822
rect 349378 223554 349406 228591
rect 349762 223554 349790 229849
rect 350146 223554 350174 229923
rect 350530 229543 350558 239834
rect 350866 239552 350894 239834
rect 351250 239552 351278 239834
rect 350866 239524 350942 239552
rect 351250 239524 351326 239552
rect 350710 238935 350762 238941
rect 350710 238877 350762 238883
rect 350722 237979 350750 238877
rect 350710 237973 350762 237979
rect 350710 237915 350762 237921
rect 350806 237973 350858 237979
rect 350806 237915 350858 237921
rect 350818 237757 350846 237915
rect 350914 237757 350942 239524
rect 350806 237751 350858 237757
rect 350806 237693 350858 237699
rect 350902 237751 350954 237757
rect 350902 237693 350954 237699
rect 351298 231393 351326 239524
rect 351586 237609 351614 239834
rect 351574 237603 351626 237609
rect 351574 237545 351626 237551
rect 351970 236888 351998 239834
rect 351970 236860 352094 236888
rect 351958 236715 352010 236721
rect 351958 236657 352010 236663
rect 351970 236351 351998 236657
rect 351958 236345 352010 236351
rect 351958 236287 352010 236293
rect 351764 234682 351820 234691
rect 351764 234617 351820 234626
rect 351670 234347 351722 234353
rect 351670 234289 351722 234295
rect 351478 234051 351530 234057
rect 351478 233993 351530 233999
rect 351382 233607 351434 233613
rect 351382 233549 351434 233555
rect 351286 231387 351338 231393
rect 351286 231329 351338 231335
rect 350518 229537 350570 229543
rect 350518 229479 350570 229485
rect 350326 228945 350378 228951
rect 350326 228887 350378 228893
rect 350338 228285 350366 228887
rect 350518 228871 350570 228877
rect 350518 228813 350570 228819
rect 350326 228279 350378 228285
rect 350326 228221 350378 228227
rect 350530 223864 350558 228813
rect 351190 227835 351242 227841
rect 351190 227777 351242 227783
rect 350902 227761 350954 227767
rect 350902 227703 350954 227709
rect 350914 223864 350942 227703
rect 350482 223836 350558 223864
rect 350866 223836 350942 223864
rect 350482 223554 350510 223836
rect 350866 223554 350894 223836
rect 351202 223554 351230 227777
rect 351394 224363 351422 233549
rect 351382 224357 351434 224363
rect 351382 224299 351434 224305
rect 351490 224215 351518 233993
rect 351574 227909 351626 227915
rect 351574 227851 351626 227857
rect 351478 224209 351530 224215
rect 351478 224151 351530 224157
rect 351586 223554 351614 227851
rect 351682 225621 351710 234289
rect 351778 225811 351806 234617
rect 351958 230055 352010 230061
rect 351958 229997 352010 230003
rect 351764 225802 351820 225811
rect 351764 225737 351820 225746
rect 351670 225615 351722 225621
rect 351670 225557 351722 225563
rect 351970 223554 351998 229997
rect 352066 227989 352094 236860
rect 352150 235383 352202 235389
rect 352150 235325 352202 235331
rect 352054 227983 352106 227989
rect 352054 227925 352106 227931
rect 352162 225769 352190 235325
rect 352354 234057 352382 239834
rect 352738 234131 352766 239834
rect 353074 239552 353102 239834
rect 353458 239552 353486 239834
rect 353074 239524 353150 239552
rect 353458 239524 353534 239552
rect 352630 234125 352682 234131
rect 352630 234067 352682 234073
rect 352726 234125 352778 234131
rect 352726 234067 352778 234073
rect 352342 234051 352394 234057
rect 352342 233993 352394 233999
rect 352642 233687 352670 234067
rect 352630 233681 352682 233687
rect 352630 233623 352682 233629
rect 353122 233613 353150 239524
rect 353206 238935 353258 238941
rect 353206 238877 353258 238883
rect 353110 233607 353162 233613
rect 353110 233549 353162 233555
rect 353218 230949 353246 238877
rect 353506 234353 353534 239524
rect 353684 237346 353740 237355
rect 353684 237281 353740 237290
rect 353590 236123 353642 236129
rect 353590 236065 353642 236071
rect 353602 235537 353630 236065
rect 353590 235531 353642 235537
rect 353590 235473 353642 235479
rect 353494 234347 353546 234353
rect 353494 234289 353546 234295
rect 353398 231461 353450 231467
rect 353398 231403 353450 231409
rect 353206 230943 353258 230949
rect 353206 230885 353258 230891
rect 352342 230129 352394 230135
rect 352342 230071 352394 230077
rect 352150 225763 352202 225769
rect 352150 225705 352202 225711
rect 352354 223554 352382 230071
rect 353012 229058 353068 229067
rect 353012 228993 353068 229002
rect 352630 228575 352682 228581
rect 352630 228517 352682 228523
rect 352642 223864 352670 228517
rect 353026 223864 353054 228993
rect 352642 223836 352718 223864
rect 353026 223836 353102 223864
rect 352690 223554 352718 223836
rect 353074 223554 353102 223836
rect 353410 223554 353438 231403
rect 353698 228933 353726 237281
rect 353794 236129 353822 239834
rect 353782 236123 353834 236129
rect 353782 236065 353834 236071
rect 354178 229543 354206 239834
rect 354562 239108 354590 239834
rect 354562 239080 354686 239108
rect 354454 238935 354506 238941
rect 354454 238877 354506 238883
rect 354550 238935 354602 238941
rect 354550 238877 354602 238883
rect 354466 238793 354494 238877
rect 354358 238787 354410 238793
rect 354358 238729 354410 238735
rect 354454 238787 354506 238793
rect 354454 238729 354506 238735
rect 354370 237036 354398 238729
rect 354562 237207 354590 238877
rect 354548 237198 354604 237207
rect 354548 237133 354604 237142
rect 354370 237008 354590 237036
rect 354454 233903 354506 233909
rect 354454 233845 354506 233851
rect 354262 233829 354314 233835
rect 354262 233771 354314 233777
rect 354070 229537 354122 229543
rect 354068 229502 354070 229511
rect 354166 229537 354218 229543
rect 354122 229502 354124 229511
rect 354166 229479 354218 229485
rect 354068 229437 354124 229446
rect 354164 229206 354220 229215
rect 354164 229141 354220 229150
rect 353698 228905 353822 228933
rect 353794 223554 353822 228905
rect 354178 223554 354206 229141
rect 354274 224511 354302 233771
rect 354262 224505 354314 224511
rect 354262 224447 354314 224453
rect 354466 224437 354494 233845
rect 354454 224431 354506 224437
rect 354454 224373 354506 224379
rect 354562 223554 354590 237008
rect 354658 236055 354686 239080
rect 354742 239009 354794 239015
rect 354742 238951 354794 238957
rect 354838 239009 354890 239015
rect 354838 238951 354890 238957
rect 354754 236795 354782 238951
rect 354850 236911 354878 238951
rect 354836 236902 354892 236911
rect 354836 236837 354892 236846
rect 354742 236789 354794 236795
rect 354742 236731 354794 236737
rect 354646 236049 354698 236055
rect 354646 235991 354698 235997
rect 354838 235309 354890 235315
rect 354838 235251 354890 235257
rect 354742 234421 354794 234427
rect 354742 234363 354794 234369
rect 354754 225473 354782 234363
rect 354742 225467 354794 225473
rect 354742 225409 354794 225415
rect 354850 225399 354878 235251
rect 354946 235241 354974 239834
rect 355282 239552 355310 239834
rect 355138 239524 355310 239552
rect 355666 239552 355694 239834
rect 355666 239524 355742 239552
rect 354934 235235 354986 235241
rect 354934 235177 354986 235183
rect 355030 235087 355082 235093
rect 355030 235029 355082 235035
rect 354934 228057 354986 228063
rect 354934 227999 354986 228005
rect 354838 225393 354890 225399
rect 354838 225335 354890 225341
rect 354946 223864 354974 227999
rect 355042 225991 355070 235029
rect 355138 234839 355166 239524
rect 355510 236715 355562 236721
rect 355510 236657 355562 236663
rect 355222 236197 355274 236203
rect 355222 236139 355274 236145
rect 355124 234830 355180 234839
rect 355124 234765 355180 234774
rect 355126 234199 355178 234205
rect 355126 234141 355178 234147
rect 355030 225985 355082 225991
rect 355030 225927 355082 225933
rect 355138 225325 355166 234141
rect 355126 225319 355178 225325
rect 355126 225261 355178 225267
rect 354898 223836 354974 223864
rect 355234 223864 355262 236139
rect 355522 225196 355550 236657
rect 355714 235315 355742 239524
rect 356002 236444 356030 239834
rect 356278 237085 356330 237091
rect 356278 237027 356330 237033
rect 356002 236416 356222 236444
rect 355702 235309 355754 235315
rect 355702 235251 355754 235257
rect 356086 234791 356138 234797
rect 356086 234733 356138 234739
rect 355894 234717 355946 234723
rect 355894 234659 355946 234665
rect 355906 234353 355934 234659
rect 355894 234347 355946 234353
rect 355894 234289 355946 234295
rect 356098 233983 356126 234733
rect 356086 233977 356138 233983
rect 356086 233919 356138 233925
rect 356194 231139 356222 236416
rect 356290 235260 356318 237027
rect 356386 235389 356414 239834
rect 356374 235383 356426 235389
rect 356374 235325 356426 235331
rect 356290 235232 356414 235260
rect 356180 231130 356236 231139
rect 356180 231065 356236 231074
rect 355990 231017 356042 231023
rect 355990 230959 356042 230965
rect 355522 225168 355646 225196
rect 355234 223836 355310 223864
rect 354898 223554 354926 223836
rect 355282 223554 355310 223836
rect 355618 223554 355646 225168
rect 356002 223554 356030 230959
rect 356278 229241 356330 229247
rect 356278 229183 356330 229189
rect 356290 228581 356318 229183
rect 356278 228575 356330 228581
rect 356278 228517 356330 228523
rect 356386 223554 356414 235232
rect 356770 234987 356798 239834
rect 357044 237050 357100 237059
rect 357044 236985 357100 236994
rect 357058 236351 357086 236985
rect 357046 236345 357098 236351
rect 357046 236287 357098 236293
rect 357044 236014 357100 236023
rect 357044 235949 357100 235958
rect 357058 235611 357086 235949
rect 357046 235605 357098 235611
rect 357046 235547 357098 235553
rect 357154 235019 357182 239834
rect 357490 239552 357518 239834
rect 357874 239552 357902 239834
rect 357490 239524 357566 239552
rect 357874 239524 357950 239552
rect 357430 236493 357482 236499
rect 357430 236435 357482 236441
rect 356854 235013 356906 235019
rect 356756 234978 356812 234987
rect 356854 234955 356906 234961
rect 357142 235013 357194 235019
rect 357142 234955 357194 234961
rect 356756 234913 356812 234922
rect 356866 233465 356894 234955
rect 356854 233459 356906 233465
rect 356854 233401 356906 233407
rect 356758 231017 356810 231023
rect 356758 230959 356810 230965
rect 356770 223554 356798 230959
rect 357442 228156 357470 236435
rect 357538 234691 357566 239524
rect 357922 235093 357950 239524
rect 358102 236863 358154 236869
rect 358102 236805 358154 236811
rect 357910 235087 357962 235093
rect 357910 235029 357962 235035
rect 357718 234939 357770 234945
rect 357718 234881 357770 234887
rect 357524 234682 357580 234691
rect 357524 234617 357580 234626
rect 357730 233835 357758 234881
rect 357718 233829 357770 233835
rect 357718 233771 357770 233777
rect 357814 230351 357866 230357
rect 357814 230293 357866 230299
rect 357826 229025 357854 230293
rect 357814 229019 357866 229025
rect 357814 228961 357866 228967
rect 357250 228128 357470 228156
rect 357814 228131 357866 228137
rect 357250 223864 357278 228128
rect 357814 228073 357866 228079
rect 357526 227613 357578 227619
rect 357526 227555 357578 227561
rect 357538 223864 357566 227555
rect 357106 223836 357278 223864
rect 357490 223836 357566 223864
rect 357106 223554 357134 223836
rect 357490 223554 357518 223836
rect 357826 223554 357854 228073
rect 358114 227601 358142 236805
rect 358210 236171 358238 239834
rect 358486 238639 358538 238645
rect 358486 238581 358538 238587
rect 358498 237091 358526 238581
rect 358486 237085 358538 237091
rect 358486 237027 358538 237033
rect 358196 236162 358252 236171
rect 358196 236097 358252 236106
rect 358292 235718 358348 235727
rect 358292 235653 358348 235662
rect 358198 229167 358250 229173
rect 358198 229109 358250 229115
rect 358210 228748 358238 229109
rect 358306 229044 358334 235653
rect 358594 234797 358622 239834
rect 358868 235126 358924 235135
rect 358868 235061 358924 235070
rect 358582 234791 358634 234797
rect 358582 234733 358634 234739
rect 358390 229537 358442 229543
rect 358390 229479 358442 229485
rect 358486 229537 358538 229543
rect 358486 229479 358538 229485
rect 358772 229502 358828 229511
rect 358402 229192 358430 229479
rect 358498 229321 358526 229479
rect 358772 229437 358828 229446
rect 358486 229315 358538 229321
rect 358486 229257 358538 229263
rect 358582 229315 358634 229321
rect 358582 229257 358634 229263
rect 358594 229192 358622 229257
rect 358402 229164 358622 229192
rect 358786 229173 358814 229437
rect 358774 229167 358826 229173
rect 358774 229109 358826 229115
rect 358306 229016 358814 229044
rect 358210 228720 358718 228748
rect 358484 228466 358540 228475
rect 358484 228401 358540 228410
rect 358390 228353 358442 228359
rect 358390 228295 358442 228301
rect 358402 227883 358430 228295
rect 358498 227989 358526 228401
rect 358582 228131 358634 228137
rect 358582 228073 358634 228079
rect 358486 227983 358538 227989
rect 358486 227925 358538 227931
rect 358388 227874 358444 227883
rect 358388 227809 358444 227818
rect 358018 227573 358142 227601
rect 358018 227527 358046 227573
rect 358018 227499 358238 227527
rect 358210 223554 358238 227499
rect 358594 223554 358622 228073
rect 358690 227989 358718 228720
rect 358678 227983 358730 227989
rect 358678 227925 358730 227931
rect 358786 225917 358814 229016
rect 358774 225911 358826 225917
rect 358774 225853 358826 225859
rect 358882 225515 358910 235061
rect 358978 233655 359006 239834
rect 359158 238787 359210 238793
rect 359158 238729 359210 238735
rect 359170 236763 359198 238729
rect 359156 236754 359212 236763
rect 359156 236689 359212 236698
rect 359254 236567 359306 236573
rect 359254 236509 359306 236515
rect 358964 233646 359020 233655
rect 358964 233581 359020 233590
rect 359156 227874 359212 227883
rect 359156 227809 359212 227818
rect 359170 227693 359198 227809
rect 358966 227687 359018 227693
rect 358966 227629 359018 227635
rect 359158 227687 359210 227693
rect 359158 227629 359210 227635
rect 358868 225506 358924 225515
rect 358868 225441 358924 225450
rect 358978 223554 359006 227629
rect 359266 223864 359294 236509
rect 359362 234945 359390 239834
rect 359698 239552 359726 239834
rect 360082 239552 360110 239834
rect 359698 239524 359774 239552
rect 360082 239524 360158 239552
rect 359638 236419 359690 236425
rect 359638 236361 359690 236367
rect 359444 235274 359500 235283
rect 359444 235209 359500 235218
rect 359350 234939 359402 234945
rect 359350 234881 359402 234887
rect 359458 225663 359486 235209
rect 359542 233755 359594 233761
rect 359542 233697 359594 233703
rect 359444 225654 359500 225663
rect 359444 225589 359500 225598
rect 359554 223887 359582 233697
rect 359540 223878 359596 223887
rect 359266 223836 359342 223864
rect 359314 223554 359342 223836
rect 359650 223864 359678 236361
rect 359746 233951 359774 239524
rect 360130 236425 360158 239524
rect 360118 236419 360170 236425
rect 360118 236361 360170 236367
rect 360418 236277 360446 239834
rect 360502 238639 360554 238645
rect 360502 238581 360554 238587
rect 360514 236615 360542 238581
rect 360598 236641 360650 236647
rect 360500 236606 360556 236615
rect 360598 236583 360650 236589
rect 360500 236541 360556 236550
rect 360310 236271 360362 236277
rect 360310 236213 360362 236219
rect 360406 236271 360458 236277
rect 360406 236213 360458 236219
rect 360322 235875 360350 236213
rect 360308 235866 360364 235875
rect 360308 235801 360364 235810
rect 360116 235718 360172 235727
rect 360116 235653 360172 235662
rect 360500 235718 360556 235727
rect 360500 235653 360556 235662
rect 360130 235537 360158 235653
rect 360118 235531 360170 235537
rect 360118 235473 360170 235479
rect 360118 235383 360170 235389
rect 360406 235383 360458 235389
rect 360170 235343 360350 235371
rect 360118 235325 360170 235331
rect 359830 234865 359882 234871
rect 359830 234807 359882 234813
rect 359732 233942 359788 233951
rect 359732 233877 359788 233886
rect 359842 226065 359870 234807
rect 359926 234273 359978 234279
rect 359926 234215 359978 234221
rect 359830 226059 359882 226065
rect 359830 226001 359882 226007
rect 359938 224881 359966 234215
rect 360322 230505 360350 235343
rect 360406 235325 360458 235331
rect 360310 230499 360362 230505
rect 360310 230441 360362 230447
rect 360020 230390 360076 230399
rect 360020 230325 360076 230334
rect 360034 228285 360062 230325
rect 360022 228279 360074 228285
rect 360022 228221 360074 228227
rect 360022 227539 360074 227545
rect 360022 227481 360074 227487
rect 359926 224875 359978 224881
rect 359926 224817 359978 224823
rect 359650 223836 359726 223864
rect 359540 223813 359596 223822
rect 359698 223554 359726 223836
rect 360034 223554 360062 227481
rect 360418 223554 360446 235325
rect 360514 224035 360542 235653
rect 360610 227545 360638 236583
rect 360692 235866 360748 235875
rect 360692 235801 360748 235810
rect 360706 235389 360734 235801
rect 360694 235383 360746 235389
rect 360694 235325 360746 235331
rect 360802 235167 360830 239834
rect 360694 235161 360746 235167
rect 360694 235103 360746 235109
rect 360790 235161 360842 235167
rect 360790 235103 360842 235109
rect 360598 227539 360650 227545
rect 360598 227481 360650 227487
rect 360706 225547 360734 235103
rect 361186 234871 361214 239834
rect 361462 237973 361514 237979
rect 361462 237915 361514 237921
rect 361174 234865 361226 234871
rect 361174 234807 361226 234813
rect 360982 234421 361034 234427
rect 360982 234363 361034 234369
rect 360994 233835 361022 234363
rect 360982 233829 361034 233835
rect 360982 233771 361034 233777
rect 361174 231683 361226 231689
rect 361174 231625 361226 231631
rect 360982 228649 361034 228655
rect 360982 228591 361034 228597
rect 361078 228649 361130 228655
rect 361078 228591 361130 228597
rect 360790 228205 360842 228211
rect 360790 228147 360842 228153
rect 360886 228205 360938 228211
rect 360886 228147 360938 228153
rect 360694 225541 360746 225547
rect 360694 225483 360746 225489
rect 360500 224026 360556 224035
rect 360500 223961 360556 223970
rect 360802 223554 360830 228147
rect 360898 228063 360926 228147
rect 360994 228063 361022 228591
rect 361090 228475 361118 228591
rect 361076 228466 361132 228475
rect 361076 228401 361132 228410
rect 360886 228057 360938 228063
rect 360886 227999 360938 228005
rect 360982 228057 361034 228063
rect 360982 227999 361034 228005
rect 361186 223554 361214 231625
rect 361474 223864 361502 237915
rect 361570 234279 361598 239834
rect 361906 239552 361934 239834
rect 362290 239552 362318 239834
rect 361906 239524 361982 239552
rect 362290 239524 362366 239552
rect 361954 234427 361982 239524
rect 362134 238417 362186 238423
rect 362134 238359 362186 238365
rect 361942 234421 361994 234427
rect 361942 234363 361994 234369
rect 361558 234273 361610 234279
rect 361558 234215 361610 234221
rect 362146 233965 362174 238359
rect 362228 235570 362284 235579
rect 362228 235505 362284 235514
rect 362242 234076 362270 235505
rect 362338 234205 362366 239524
rect 362420 235422 362476 235431
rect 362420 235357 362476 235366
rect 362326 234199 362378 234205
rect 362326 234141 362378 234147
rect 362242 234048 362366 234076
rect 362146 233937 362270 233965
rect 361846 228501 361898 228507
rect 361846 228443 361898 228449
rect 361858 223864 361886 228443
rect 361474 223836 361550 223864
rect 361858 223836 361934 223864
rect 361522 223554 361550 223836
rect 361906 223554 361934 223836
rect 362242 223554 362270 233937
rect 362338 225695 362366 234048
rect 362434 225843 362462 235357
rect 362626 235283 362654 239834
rect 362612 235274 362668 235283
rect 362612 235209 362668 235218
rect 362806 234125 362858 234131
rect 362806 234067 362858 234073
rect 362818 233539 362846 234067
rect 362710 233533 362762 233539
rect 362710 233475 362762 233481
rect 362806 233533 362858 233539
rect 362806 233475 362858 233481
rect 362614 231535 362666 231541
rect 362614 231477 362666 231483
rect 362422 225837 362474 225843
rect 362422 225779 362474 225785
rect 362326 225689 362378 225695
rect 362326 225631 362378 225637
rect 362626 223554 362654 231477
rect 362722 223887 362750 233475
rect 363010 231467 363038 239834
rect 363394 234099 363422 239834
rect 363478 234347 363530 234353
rect 363478 234289 363530 234295
rect 363380 234090 363436 234099
rect 363380 234025 363436 234034
rect 363382 232793 363434 232799
rect 363382 232735 363434 232741
rect 362998 231461 363050 231467
rect 362998 231403 363050 231409
rect 362998 231165 363050 231171
rect 362998 231107 363050 231113
rect 362708 223878 362764 223887
rect 362708 223813 362764 223822
rect 363010 223554 363038 231107
rect 363394 223554 363422 232735
rect 363490 225029 363518 234289
rect 363574 233977 363626 233983
rect 363574 233919 363626 233925
rect 363586 225177 363614 233919
rect 363670 231757 363722 231763
rect 363670 231699 363722 231705
rect 363574 225171 363626 225177
rect 363574 225113 363626 225119
rect 363478 225023 363530 225029
rect 363478 224965 363530 224971
rect 363682 223864 363710 231699
rect 363778 231541 363806 239834
rect 364114 239552 364142 239834
rect 364498 239552 364526 239834
rect 364114 239524 364190 239552
rect 364498 239524 364574 239552
rect 364162 235135 364190 239524
rect 364148 235126 364204 235135
rect 364148 235061 364204 235070
rect 364546 233909 364574 239524
rect 364726 237011 364778 237017
rect 364726 236953 364778 236959
rect 364534 233903 364586 233909
rect 364534 233845 364586 233851
rect 363766 231535 363818 231541
rect 363766 231477 363818 231483
rect 364054 231091 364106 231097
rect 364054 231033 364106 231039
rect 363862 224135 363914 224141
rect 363862 224077 363914 224083
rect 363874 223919 363902 224077
rect 363862 223913 363914 223919
rect 363682 223836 363758 223864
rect 363862 223855 363914 223861
rect 364066 223864 364094 231033
rect 364438 230869 364490 230875
rect 364438 230811 364490 230817
rect 364342 224135 364394 224141
rect 364342 224077 364394 224083
rect 364354 223919 364382 224077
rect 364342 223913 364394 223919
rect 364244 223878 364300 223887
rect 364066 223836 364142 223864
rect 363730 223554 363758 223836
rect 364114 223554 364142 223836
rect 364342 223855 364394 223861
rect 364244 223813 364246 223822
rect 364298 223813 364300 223822
rect 364246 223781 364298 223787
rect 364450 223554 364478 230811
rect 364738 225196 364766 236953
rect 364834 232799 364862 239834
rect 365218 233835 365246 239834
rect 365602 239256 365630 239834
rect 365410 239228 365630 239256
rect 365302 236937 365354 236943
rect 365302 236879 365354 236885
rect 365110 233829 365162 233835
rect 365110 233771 365162 233777
rect 365206 233829 365258 233835
rect 365206 233771 365258 233777
rect 365122 233632 365150 233771
rect 365122 233604 365246 233632
rect 365218 233465 365246 233604
rect 365110 233459 365162 233465
rect 365110 233401 365162 233407
rect 365206 233459 365258 233465
rect 365206 233401 365258 233407
rect 364822 232793 364874 232799
rect 364822 232735 364874 232741
rect 365122 225251 365150 233401
rect 365314 228563 365342 236879
rect 365410 235431 365438 239228
rect 365494 239083 365546 239089
rect 365494 239025 365546 239031
rect 365506 238035 365534 239025
rect 365686 238047 365738 238053
rect 365506 238007 365686 238035
rect 365686 237989 365738 237995
rect 365396 235422 365452 235431
rect 365396 235357 365452 235366
rect 365986 234353 366014 239834
rect 366322 239552 366350 239834
rect 366706 239681 366734 239834
rect 366694 239675 366746 239681
rect 366694 239617 366746 239623
rect 366322 239524 366398 239552
rect 366370 237979 366398 239524
rect 366358 237973 366410 237979
rect 366358 237915 366410 237921
rect 367042 235579 367070 239834
rect 367028 235570 367084 235579
rect 367028 235505 367084 235514
rect 365974 234347 366026 234353
rect 365974 234289 366026 234295
rect 366646 233755 366698 233761
rect 366646 233697 366698 233703
rect 366658 233632 366686 233697
rect 367126 233681 367178 233687
rect 366658 233604 366782 233632
rect 367126 233623 367178 233629
rect 366454 233459 366506 233465
rect 366454 233401 366506 233407
rect 365494 230943 365546 230949
rect 365494 230885 365546 230891
rect 365218 228535 365342 228563
rect 365110 225245 365162 225251
rect 364738 225168 364862 225196
rect 365110 225187 365162 225193
rect 364630 224283 364682 224289
rect 364630 224225 364682 224231
rect 364642 224067 364670 224225
rect 364630 224061 364682 224067
rect 364630 224003 364682 224009
rect 364834 223554 364862 225168
rect 365218 223554 365246 228535
rect 365506 225196 365534 230885
rect 366466 228877 366494 233401
rect 366646 229241 366698 229247
rect 366646 229183 366698 229189
rect 366454 228871 366506 228877
rect 366454 228813 366506 228819
rect 366262 228797 366314 228803
rect 366262 228739 366314 228745
rect 365878 228723 365930 228729
rect 365878 228665 365930 228671
rect 365506 225168 365630 225196
rect 365602 223554 365630 225168
rect 365890 223864 365918 228665
rect 366274 223864 366302 228739
rect 365890 223836 365966 223864
rect 366274 223836 366350 223864
rect 365938 223554 365966 223836
rect 366322 223554 366350 223836
rect 366658 223554 366686 229183
rect 366754 225103 366782 233604
rect 367030 228575 367082 228581
rect 367030 228517 367082 228523
rect 366742 225097 366794 225103
rect 366742 225039 366794 225045
rect 367042 223554 367070 228517
rect 367138 224183 367166 233623
rect 367426 231560 367454 239834
rect 367606 233533 367658 233539
rect 367606 233475 367658 233481
rect 367426 231532 367550 231560
rect 367414 230351 367466 230357
rect 367414 230293 367466 230299
rect 367124 224174 367180 224183
rect 367124 224109 367180 224118
rect 367426 223554 367454 230293
rect 367522 230209 367550 231532
rect 367618 230357 367646 233475
rect 367606 230351 367658 230357
rect 367606 230293 367658 230299
rect 367510 230203 367562 230209
rect 367510 230145 367562 230151
rect 367810 229215 367838 239834
rect 367990 234347 368042 234353
rect 367990 234289 368042 234295
rect 367894 229315 367946 229321
rect 367894 229257 367946 229263
rect 367796 229206 367852 229215
rect 367796 229141 367852 229150
rect 367906 229025 367934 229257
rect 367798 229019 367850 229025
rect 367798 228961 367850 228967
rect 367894 229019 367946 229025
rect 367894 228961 367946 228967
rect 367810 223554 367838 228961
rect 368002 228803 368030 234289
rect 368084 229650 368140 229659
rect 368194 229617 368222 239834
rect 368530 239552 368558 239834
rect 368914 239552 368942 239834
rect 368530 239524 368606 239552
rect 368914 239524 368990 239552
rect 368578 236023 368606 239524
rect 368564 236014 368620 236023
rect 368564 235949 368620 235958
rect 368662 234347 368714 234353
rect 368662 234289 368714 234295
rect 368674 234205 368702 234289
rect 368662 234199 368714 234205
rect 368662 234141 368714 234147
rect 368662 233829 368714 233835
rect 368662 233771 368714 233777
rect 368674 233539 368702 233771
rect 368662 233533 368714 233539
rect 368662 233475 368714 233481
rect 368566 233385 368618 233391
rect 368662 233385 368714 233391
rect 368618 233345 368662 233373
rect 368566 233327 368618 233333
rect 368662 233327 368714 233333
rect 368854 230277 368906 230283
rect 368854 230219 368906 230225
rect 368084 229585 368086 229594
rect 368138 229585 368140 229594
rect 368182 229611 368234 229617
rect 368086 229553 368138 229559
rect 368182 229553 368234 229559
rect 368182 229167 368234 229173
rect 368182 229109 368234 229115
rect 367990 228797 368042 228803
rect 367990 228739 368042 228745
rect 368194 228359 368222 229109
rect 368470 228945 368522 228951
rect 368470 228887 368522 228893
rect 368374 228649 368426 228655
rect 368374 228591 368426 228597
rect 368086 228353 368138 228359
rect 368086 228295 368138 228301
rect 368182 228353 368234 228359
rect 368182 228295 368234 228301
rect 368098 223864 368126 228295
rect 368386 224955 368414 228591
rect 368374 224949 368426 224955
rect 368374 224891 368426 224897
rect 368482 224493 368510 228887
rect 368290 224465 368510 224493
rect 368290 223864 368318 224465
rect 368098 223836 368174 223864
rect 368290 223836 368558 223864
rect 368146 223554 368174 223836
rect 368530 223554 368558 223836
rect 368866 223554 368894 230219
rect 368962 228581 368990 239524
rect 369250 229363 369278 239834
rect 369526 230425 369578 230431
rect 369526 230367 369578 230373
rect 369430 230203 369482 230209
rect 369430 230145 369482 230151
rect 369236 229354 369292 229363
rect 369236 229289 369292 229298
rect 369442 229247 369470 230145
rect 369430 229241 369482 229247
rect 369430 229183 369482 229189
rect 368950 228575 369002 228581
rect 368950 228517 369002 228523
rect 369238 227983 369290 227989
rect 369238 227925 369290 227931
rect 369250 223554 369278 227925
rect 369538 225196 369566 230367
rect 369634 230209 369662 239834
rect 370018 235727 370046 239834
rect 370004 235718 370060 235727
rect 370004 235653 370060 235662
rect 370402 230357 370430 239834
rect 370738 239552 370766 239834
rect 370690 239524 370766 239552
rect 371122 239552 371150 239834
rect 371458 239700 371486 239834
rect 371362 239672 371486 239700
rect 371122 239524 371198 239552
rect 370294 230351 370346 230357
rect 370294 230293 370346 230299
rect 370390 230351 370442 230357
rect 370390 230293 370442 230299
rect 369622 230203 369674 230209
rect 369622 230145 369674 230151
rect 370198 229463 370250 229469
rect 370198 229405 370250 229411
rect 370210 228951 370238 229405
rect 370306 229173 370334 230293
rect 370390 229463 370442 229469
rect 370390 229405 370442 229411
rect 370294 229167 370346 229173
rect 370294 229109 370346 229115
rect 370198 228945 370250 228951
rect 370198 228887 370250 228893
rect 370006 228723 370058 228729
rect 370006 228665 370058 228671
rect 369538 225168 369662 225196
rect 369634 223554 369662 225168
rect 370018 223554 370046 228665
rect 370402 223864 370430 229405
rect 370690 229067 370718 239524
rect 371170 233687 371198 239524
rect 371362 235875 371390 239672
rect 371348 235866 371404 235875
rect 371348 235801 371404 235810
rect 371158 233681 371210 233687
rect 371158 233623 371210 233629
rect 371062 230425 371114 230431
rect 371842 230376 371870 239834
rect 371926 233681 371978 233687
rect 371926 233623 371978 233629
rect 371062 230367 371114 230373
rect 370774 230277 370826 230283
rect 370774 230219 370826 230225
rect 370676 229058 370732 229067
rect 370676 228993 370732 229002
rect 370786 223864 370814 230219
rect 370354 223836 370430 223864
rect 370738 223836 370814 223864
rect 370354 223554 370382 223836
rect 370738 223554 370766 223836
rect 371074 223554 371102 230367
rect 371458 230348 371870 230376
rect 371458 223554 371486 230348
rect 371938 225196 371966 233623
rect 372226 230547 372254 239834
rect 372310 233681 372362 233687
rect 372310 233623 372362 233629
rect 372322 233317 372350 233623
rect 372310 233311 372362 233317
rect 372310 233253 372362 233259
rect 372212 230538 372268 230547
rect 372212 230473 372268 230482
rect 372610 230431 372638 239834
rect 372946 239552 372974 239834
rect 373330 239552 373358 239834
rect 372946 239524 373022 239552
rect 372994 235093 373022 239524
rect 373282 239524 373358 239552
rect 372790 235087 372842 235093
rect 372790 235029 372842 235035
rect 372982 235087 373034 235093
rect 372982 235029 373034 235035
rect 372694 231387 372746 231393
rect 372694 231329 372746 231335
rect 372598 230425 372650 230431
rect 372598 230367 372650 230373
rect 372214 230351 372266 230357
rect 372214 230293 372266 230299
rect 371842 225168 371966 225196
rect 371842 223554 371870 225168
rect 372226 223554 372254 230293
rect 372502 230203 372554 230209
rect 372502 230145 372554 230151
rect 372514 223864 372542 230145
rect 372706 229099 372734 231329
rect 372694 229093 372746 229099
rect 372694 229035 372746 229041
rect 372802 228507 372830 235029
rect 373282 230283 373310 239524
rect 373666 230283 373694 239834
rect 373942 239675 373994 239681
rect 373942 239617 373994 239623
rect 373750 231239 373802 231245
rect 373750 231181 373802 231187
rect 373270 230277 373322 230283
rect 373270 230219 373322 230225
rect 373654 230277 373706 230283
rect 373654 230219 373706 230225
rect 373762 230209 373790 231181
rect 373750 230203 373802 230209
rect 373750 230145 373802 230151
rect 373364 229650 373420 229659
rect 373270 229611 373322 229617
rect 373364 229585 373366 229594
rect 373270 229553 373322 229559
rect 373418 229585 373420 229594
rect 373366 229553 373418 229559
rect 372886 228575 372938 228581
rect 372886 228517 372938 228523
rect 372790 228501 372842 228507
rect 372790 228443 372842 228449
rect 372898 223864 372926 228517
rect 372514 223836 372590 223864
rect 372898 223836 372974 223864
rect 372562 223554 372590 223836
rect 372946 223554 372974 223836
rect 373282 223554 373310 229553
rect 373654 229241 373706 229247
rect 373654 229183 373706 229189
rect 373666 223554 373694 229183
rect 373954 224160 373982 239617
rect 374050 229469 374078 239834
rect 374434 235907 374462 239834
rect 374326 235901 374378 235907
rect 374326 235843 374378 235849
rect 374422 235901 374474 235907
rect 374422 235843 374474 235849
rect 374338 233909 374366 235843
rect 374326 233903 374378 233909
rect 374326 233845 374378 233851
rect 374710 233533 374762 233539
rect 374710 233475 374762 233481
rect 374326 232793 374378 232799
rect 374326 232735 374378 232741
rect 374038 229463 374090 229469
rect 374038 229405 374090 229411
rect 374338 228475 374366 232735
rect 374422 228797 374474 228803
rect 374422 228739 374474 228745
rect 374324 228466 374380 228475
rect 374324 228401 374380 228410
rect 373954 224132 374078 224160
rect 374050 223554 374078 224132
rect 374434 223554 374462 228739
rect 374722 223864 374750 233475
rect 374818 228729 374846 239834
rect 375154 239552 375182 239834
rect 375538 239552 375566 239834
rect 375154 239524 375230 239552
rect 375538 239524 375614 239552
rect 374998 235975 375050 235981
rect 374998 235917 375050 235923
rect 375094 235975 375146 235981
rect 375094 235917 375146 235923
rect 375010 234205 375038 235917
rect 375106 235685 375134 235917
rect 375094 235679 375146 235685
rect 375094 235621 375146 235627
rect 374998 234199 375050 234205
rect 374998 234141 375050 234147
rect 375094 233977 375146 233983
rect 375094 233919 375146 233925
rect 374806 228723 374858 228729
rect 374806 228665 374858 228671
rect 374998 224875 375050 224881
rect 374998 224817 375050 224823
rect 375010 224585 375038 224817
rect 374998 224579 375050 224585
rect 374998 224521 375050 224527
rect 375106 223864 375134 233919
rect 375202 229469 375230 239524
rect 375286 235679 375338 235685
rect 375286 235621 375338 235627
rect 375298 235537 375326 235621
rect 375286 235531 375338 235537
rect 375286 235473 375338 235479
rect 375382 235013 375434 235019
rect 375382 234955 375434 234961
rect 375190 229463 375242 229469
rect 375190 229405 375242 229411
rect 375394 228581 375422 234955
rect 375586 234945 375614 239524
rect 375574 234939 375626 234945
rect 375574 234881 375626 234887
rect 375874 234668 375902 239834
rect 376258 235167 376286 239834
rect 376246 235161 376298 235167
rect 376246 235103 376298 235109
rect 375874 234640 376094 234668
rect 375958 234569 376010 234575
rect 375958 234511 376010 234517
rect 375970 234131 375998 234511
rect 375958 234125 376010 234131
rect 375958 234067 376010 234073
rect 375478 231535 375530 231541
rect 375478 231477 375530 231483
rect 375382 228575 375434 228581
rect 375382 228517 375434 228523
rect 374722 223836 374798 223864
rect 375106 223836 375182 223864
rect 374770 223554 374798 223836
rect 375154 223554 375182 223836
rect 375490 223554 375518 231477
rect 375862 231461 375914 231467
rect 375862 231403 375914 231409
rect 375874 223554 375902 231403
rect 376066 228803 376094 234640
rect 376246 234347 376298 234353
rect 376246 234289 376298 234295
rect 376054 228797 376106 228803
rect 376054 228739 376106 228745
rect 376258 223554 376286 234289
rect 376534 234273 376586 234279
rect 376534 234215 376586 234221
rect 376546 228600 376574 234215
rect 376642 233928 376670 239834
rect 377026 235463 377054 239834
rect 377362 239552 377390 239834
rect 377746 239552 377774 239834
rect 377362 239524 377438 239552
rect 377746 239524 377822 239552
rect 377302 236419 377354 236425
rect 377302 236361 377354 236367
rect 377110 236271 377162 236277
rect 377110 236213 377162 236219
rect 377014 235457 377066 235463
rect 377014 235399 377066 235405
rect 376822 235235 376874 235241
rect 376822 235177 376874 235183
rect 376642 233900 376766 233928
rect 376738 229247 376766 233900
rect 376726 229241 376778 229247
rect 376726 229183 376778 229189
rect 376546 228572 376670 228600
rect 376642 223554 376670 228572
rect 376834 223864 376862 235177
rect 376918 233755 376970 233761
rect 376918 233697 376970 233703
rect 376930 233465 376958 233697
rect 377122 233465 377150 236213
rect 377206 235901 377258 235907
rect 377206 235843 377258 235849
rect 377218 234279 377246 235843
rect 377206 234273 377258 234279
rect 377206 234215 377258 234221
rect 376918 233459 376970 233465
rect 376918 233401 376970 233407
rect 377110 233459 377162 233465
rect 377110 233401 377162 233407
rect 377314 223864 377342 236361
rect 377410 231583 377438 239524
rect 377686 235013 377738 235019
rect 377686 234955 377738 234961
rect 377396 231574 377452 231583
rect 377396 231509 377452 231518
rect 376834 223836 377006 223864
rect 377314 223836 377390 223864
rect 376978 223554 377006 223836
rect 377362 223554 377390 223836
rect 377698 223554 377726 234955
rect 377794 234723 377822 239524
rect 378082 234964 378110 239834
rect 378466 235019 378494 239834
rect 378850 236000 378878 239834
rect 378850 235972 378974 236000
rect 378838 235827 378890 235833
rect 378838 235769 378890 235775
rect 378454 235013 378506 235019
rect 378082 234936 378206 234964
rect 378454 234955 378506 234961
rect 378070 234791 378122 234797
rect 378070 234733 378122 234739
rect 377782 234717 377834 234723
rect 377782 234659 377834 234665
rect 378082 223554 378110 234733
rect 378178 229955 378206 234936
rect 378742 234865 378794 234871
rect 378742 234807 378794 234813
rect 378646 234643 378698 234649
rect 378646 234585 378698 234591
rect 378658 233983 378686 234585
rect 378646 233977 378698 233983
rect 378646 233919 378698 233925
rect 378754 233539 378782 234807
rect 378850 234649 378878 235769
rect 378838 234643 378890 234649
rect 378838 234585 378890 234591
rect 378742 233533 378794 233539
rect 378742 233475 378794 233481
rect 378164 229946 378220 229955
rect 378164 229881 378220 229890
rect 378946 228771 378974 235972
rect 379234 235241 379262 239834
rect 379570 239552 379598 239834
rect 379954 239552 379982 239834
rect 379570 239524 379646 239552
rect 379954 239524 380030 239552
rect 379510 235383 379562 235389
rect 379510 235325 379562 235331
rect 379222 235235 379274 235241
rect 379222 235177 379274 235183
rect 379126 230499 379178 230505
rect 379126 230441 379178 230447
rect 378932 228762 378988 228771
rect 378932 228697 378988 228706
rect 378838 228575 378890 228581
rect 378838 228517 378890 228523
rect 378454 228501 378506 228507
rect 378454 228443 378506 228449
rect 378466 223554 378494 228443
rect 378646 227983 378698 227989
rect 378646 227925 378698 227931
rect 378658 227619 378686 227925
rect 378646 227613 378698 227619
rect 378646 227555 378698 227561
rect 378550 224061 378602 224067
rect 378550 224003 378602 224009
rect 378562 223845 378590 224003
rect 378550 223839 378602 223845
rect 378550 223781 378602 223787
rect 378850 223554 378878 228517
rect 379138 223864 379166 230441
rect 379318 223987 379370 223993
rect 379318 223929 379370 223935
rect 379138 223836 379214 223864
rect 379330 223845 379358 223929
rect 379412 223878 379468 223887
rect 379186 223554 379214 223836
rect 379318 223839 379370 223845
rect 379522 223864 379550 235325
rect 379618 230103 379646 239524
rect 380002 235389 380030 239524
rect 379990 235383 380042 235389
rect 379990 235325 380042 235331
rect 379894 235309 379946 235315
rect 379894 235251 379946 235257
rect 379604 230094 379660 230103
rect 379604 230029 379660 230038
rect 379522 223836 379598 223864
rect 379412 223813 379414 223822
rect 379318 223781 379370 223787
rect 379466 223813 379468 223822
rect 379414 223781 379466 223787
rect 379570 223554 379598 223836
rect 379906 223554 379934 235251
rect 380290 233211 380318 239834
rect 380674 234797 380702 239834
rect 380662 234791 380714 234797
rect 380662 234733 380714 234739
rect 380276 233202 380332 233211
rect 380276 233137 380332 233146
rect 381058 229340 381086 239834
rect 381442 234945 381470 239834
rect 381526 239675 381578 239681
rect 381526 239617 381578 239623
rect 381538 239533 381566 239617
rect 381778 239552 381806 239834
rect 382162 239552 382190 239834
rect 381526 239527 381578 239533
rect 381778 239524 381854 239552
rect 382162 239524 382238 239552
rect 381526 239469 381578 239475
rect 381430 234939 381482 234945
rect 381430 234881 381482 234887
rect 381826 229807 381854 239524
rect 382210 235315 382238 239524
rect 382198 235309 382250 235315
rect 382198 235251 382250 235257
rect 382498 230376 382526 239834
rect 382882 235463 382910 239834
rect 382870 235457 382922 235463
rect 382870 235399 382922 235405
rect 383266 231731 383294 239834
rect 383348 237050 383404 237059
rect 383348 236985 383404 236994
rect 383252 231722 383308 231731
rect 383252 231657 383308 231666
rect 382498 230348 382622 230376
rect 382486 230203 382538 230209
rect 382486 230145 382538 230151
rect 381812 229798 381868 229807
rect 381812 229733 381868 229742
rect 381058 229312 381182 229340
rect 381046 229167 381098 229173
rect 381046 229109 381098 229115
rect 380278 229019 380330 229025
rect 380278 228961 380330 228967
rect 380566 229019 380618 229025
rect 380566 228961 380618 228967
rect 380290 223554 380318 228961
rect 380578 228803 380606 228961
rect 380662 228871 380714 228877
rect 380662 228813 380714 228819
rect 380566 228797 380618 228803
rect 380566 228739 380618 228745
rect 380674 223554 380702 228813
rect 381058 223554 381086 229109
rect 381154 227735 381182 229312
rect 381718 229093 381770 229099
rect 381718 229035 381770 229041
rect 381140 227726 381196 227735
rect 381140 227661 381196 227670
rect 381334 224949 381386 224955
rect 381334 224891 381386 224897
rect 381346 223864 381374 224891
rect 381730 223864 381758 229035
rect 382102 228353 382154 228359
rect 382102 228295 382154 228301
rect 381346 223836 381422 223864
rect 381730 223836 381806 223864
rect 381394 223554 381422 223836
rect 381778 223554 381806 223836
rect 382114 223554 382142 228295
rect 382498 223554 382526 230145
rect 382594 228623 382622 230348
rect 382870 230277 382922 230283
rect 382870 230219 382922 230225
rect 382774 229463 382826 229469
rect 382774 229405 382826 229411
rect 382786 229247 382814 229405
rect 382774 229241 382826 229247
rect 382774 229183 382826 229189
rect 382882 229173 382910 230219
rect 382870 229167 382922 229173
rect 382870 229109 382922 229115
rect 382580 228614 382636 228623
rect 382580 228549 382636 228558
rect 382870 228575 382922 228581
rect 382870 228517 382922 228523
rect 382882 223554 382910 228517
rect 383362 225196 383390 236985
rect 383650 233063 383678 239834
rect 383986 239552 384014 239834
rect 383938 239524 384014 239552
rect 384370 239552 384398 239834
rect 384370 239524 384446 239552
rect 383636 233054 383692 233063
rect 383636 232989 383692 232998
rect 383638 230573 383690 230579
rect 383638 230515 383690 230521
rect 383266 225168 383390 225196
rect 383266 223554 383294 225168
rect 383650 223864 383678 230515
rect 383938 230251 383966 239524
rect 384418 233359 384446 239524
rect 384404 233350 384460 233359
rect 384404 233285 384460 233294
rect 383924 230242 383980 230251
rect 383924 230177 383980 230186
rect 384706 229511 384734 239834
rect 385090 234543 385118 239834
rect 385172 237346 385228 237355
rect 385172 237281 385228 237290
rect 385076 234534 385132 234543
rect 385076 234469 385132 234478
rect 384790 231239 384842 231245
rect 384790 231181 384842 231187
rect 384692 229502 384748 229511
rect 384692 229437 384748 229446
rect 384310 228871 384362 228877
rect 384310 228813 384362 228819
rect 384022 227539 384074 227545
rect 384022 227481 384074 227487
rect 384034 223864 384062 227481
rect 383602 223836 383678 223864
rect 383986 223836 384062 223864
rect 383602 223554 383630 223836
rect 383986 223554 384014 223836
rect 384322 223554 384350 228813
rect 384802 225196 384830 231181
rect 385186 225196 385214 237281
rect 385474 229659 385502 239834
rect 385556 239566 385612 239575
rect 385556 239501 385612 239510
rect 385460 229650 385516 229659
rect 385460 229585 385516 229594
rect 385570 225196 385598 239501
rect 385858 234395 385886 239834
rect 386194 239552 386222 239834
rect 386578 239552 386606 239834
rect 386146 239524 386222 239552
rect 386530 239524 386606 239552
rect 385844 234386 385900 234395
rect 385844 234321 385900 234330
rect 386146 233095 386174 239524
rect 386530 233169 386558 239524
rect 386914 233761 386942 239834
rect 387298 238349 387326 239834
rect 387286 238343 387338 238349
rect 387286 238285 387338 238291
rect 387682 233835 387710 239834
rect 387956 236754 388012 236763
rect 387956 236689 388012 236698
rect 387670 233829 387722 233835
rect 387670 233771 387722 233777
rect 386902 233755 386954 233761
rect 386902 233697 386954 233703
rect 386518 233163 386570 233169
rect 386518 233105 386570 233111
rect 386134 233089 386186 233095
rect 386134 233031 386186 233037
rect 386518 231535 386570 231541
rect 386518 231477 386570 231483
rect 384706 225168 384830 225196
rect 385090 225168 385214 225196
rect 385474 225168 385598 225196
rect 384706 223554 384734 225168
rect 385090 223554 385118 225168
rect 385474 223554 385502 225168
rect 386228 225062 386284 225071
rect 386228 224997 386284 225006
rect 385844 224914 385900 224923
rect 385844 224849 385900 224858
rect 385858 223716 385886 224849
rect 386242 223827 386270 224997
rect 385810 223688 385886 223716
rect 386194 223799 386270 223827
rect 385810 223554 385838 223688
rect 386194 223554 386222 223799
rect 386530 223554 386558 231477
rect 387670 230721 387722 230727
rect 387670 230663 387722 230669
rect 387286 230277 387338 230283
rect 387286 230219 387338 230225
rect 386902 227613 386954 227619
rect 386902 227555 386954 227561
rect 386914 223554 386942 227555
rect 387298 223554 387326 230219
rect 387682 223554 387710 230663
rect 387970 223864 387998 236689
rect 388066 234353 388094 239834
rect 388402 239552 388430 239834
rect 388786 239700 388814 239834
rect 388354 239524 388430 239552
rect 388738 239672 388814 239700
rect 388918 239675 388970 239681
rect 388354 238835 388382 239524
rect 388340 238826 388396 238835
rect 388340 238761 388396 238770
rect 388054 234347 388106 234353
rect 388054 234289 388106 234295
rect 388342 233903 388394 233909
rect 388342 233845 388394 233851
rect 387970 223836 388046 223864
rect 388018 223554 388046 223836
rect 388354 223827 388382 233845
rect 388738 233243 388766 239672
rect 388918 239617 388970 239623
rect 388930 239311 388958 239617
rect 388918 239305 388970 239311
rect 388918 239247 388970 239253
rect 389122 235833 389150 239834
rect 389506 236911 389534 239834
rect 389890 239131 389918 239834
rect 389876 239122 389932 239131
rect 389876 239057 389932 239066
rect 390166 238417 390218 238423
rect 390166 238359 390218 238365
rect 390178 238053 390206 238359
rect 390166 238047 390218 238053
rect 390166 237989 390218 237995
rect 389492 236902 389548 236911
rect 389492 236837 389548 236846
rect 389206 236567 389258 236573
rect 389206 236509 389258 236515
rect 389110 235827 389162 235833
rect 389110 235769 389162 235775
rect 388726 233237 388778 233243
rect 388726 233179 388778 233185
rect 389218 229192 389246 236509
rect 390166 236197 390218 236203
rect 390166 236139 390218 236145
rect 390178 235611 390206 236139
rect 390166 235605 390218 235611
rect 390166 235547 390218 235553
rect 389684 232166 389740 232175
rect 389684 232101 389740 232110
rect 389698 231287 389726 232101
rect 389684 231278 389740 231287
rect 389684 231213 389740 231222
rect 389878 230943 389930 230949
rect 389878 230885 389930 230891
rect 389494 230795 389546 230801
rect 389494 230737 389546 230743
rect 389122 229164 389246 229192
rect 388726 228723 388778 228729
rect 388726 228665 388778 228671
rect 388738 224775 388766 228665
rect 388724 224766 388780 224775
rect 388724 224701 388780 224710
rect 388724 223878 388780 223887
rect 388354 223799 388430 223827
rect 388724 223813 388780 223822
rect 388402 223554 388430 223799
rect 388738 223554 388766 223813
rect 389122 223554 389150 229164
rect 389506 223554 389534 230737
rect 389890 223554 389918 230885
rect 390274 229488 390302 239834
rect 390610 239552 390638 239834
rect 390994 239552 391022 239834
rect 390610 239524 390686 239552
rect 390994 239524 391070 239552
rect 390658 238983 390686 239524
rect 390644 238974 390700 238983
rect 390644 238909 390700 238918
rect 390550 234643 390602 234649
rect 390550 234585 390602 234591
rect 390274 229460 390398 229488
rect 390262 228427 390314 228433
rect 390262 228369 390314 228375
rect 390274 223716 390302 228369
rect 390370 223887 390398 229460
rect 390356 223878 390412 223887
rect 390562 223864 390590 234585
rect 390934 231091 390986 231097
rect 390934 231033 390986 231039
rect 390562 223836 390638 223864
rect 390356 223813 390412 223822
rect 390226 223688 390302 223716
rect 390226 223554 390254 223688
rect 390610 223554 390638 223836
rect 390946 223554 390974 231033
rect 391042 225219 391070 239524
rect 391330 239163 391358 239834
rect 391318 239157 391370 239163
rect 391318 239099 391370 239105
rect 391714 239089 391742 239834
rect 391702 239083 391754 239089
rect 391702 239025 391754 239031
rect 392098 238835 392126 239834
rect 392084 238826 392140 238835
rect 392084 238761 392140 238770
rect 392482 238539 392510 239834
rect 392818 239552 392846 239834
rect 392770 239524 392846 239552
rect 393202 239552 393230 239834
rect 393202 239524 393278 239552
rect 392662 239083 392714 239089
rect 392662 239025 392714 239031
rect 392674 238539 392702 239025
rect 392468 238530 392524 238539
rect 392468 238465 392524 238474
rect 392660 238530 392716 238539
rect 392660 238465 392716 238474
rect 391510 235975 391562 235981
rect 391510 235917 391562 235923
rect 391126 232497 391178 232503
rect 391126 232439 391178 232445
rect 391138 231171 391166 232439
rect 391414 232423 391466 232429
rect 391414 232365 391466 232371
rect 391426 232300 391454 232365
rect 391234 232272 391454 232300
rect 391234 232207 391262 232272
rect 391222 232201 391274 232207
rect 391222 232143 391274 232149
rect 391414 231461 391466 231467
rect 391234 231421 391414 231449
rect 391234 231319 391262 231421
rect 391414 231403 391466 231409
rect 391222 231313 391274 231319
rect 391222 231255 391274 231261
rect 391126 231165 391178 231171
rect 391126 231107 391178 231113
rect 391522 229451 391550 235917
rect 392470 233681 392522 233687
rect 392470 233623 392522 233629
rect 391606 231387 391658 231393
rect 391606 231329 391658 231335
rect 391330 229423 391550 229451
rect 391028 225210 391084 225219
rect 391028 225145 391084 225154
rect 391330 223554 391358 229423
rect 391618 227545 391646 231329
rect 392086 230869 392138 230875
rect 392086 230811 392138 230817
rect 391702 230647 391754 230653
rect 391702 230589 391754 230595
rect 391606 227539 391658 227545
rect 391606 227481 391658 227487
rect 391714 224775 391742 230589
rect 391700 224766 391756 224775
rect 391700 224701 391756 224710
rect 391894 224283 391946 224289
rect 391894 224225 391946 224231
rect 391906 224183 391934 224225
rect 391892 224174 391948 224183
rect 391892 224109 391948 224118
rect 391700 223878 391756 223887
rect 391700 223813 391756 223822
rect 391714 223554 391742 223813
rect 392098 223554 392126 230811
rect 392482 223864 392510 233623
rect 392770 224183 392798 239524
rect 392854 238343 392906 238349
rect 392854 238285 392906 238291
rect 392756 224174 392812 224183
rect 392756 224109 392812 224118
rect 392866 223864 392894 238285
rect 393046 231165 393098 231171
rect 393046 231107 393098 231113
rect 393058 228179 393086 231107
rect 393044 228170 393100 228179
rect 393044 228105 393100 228114
rect 393140 228022 393196 228031
rect 393140 227957 393196 227966
rect 392434 223836 392510 223864
rect 392818 223836 392894 223864
rect 392434 223554 392462 223836
rect 392818 223554 392846 223836
rect 393154 223554 393182 227957
rect 393250 225367 393278 239524
rect 393538 234427 393566 239834
rect 393922 238053 393950 239834
rect 393910 238047 393962 238053
rect 393910 237989 393962 237995
rect 393430 234421 393482 234427
rect 393430 234363 393482 234369
rect 393526 234421 393578 234427
rect 393526 234363 393578 234369
rect 393442 233835 393470 234363
rect 393430 233829 393482 233835
rect 393430 233771 393482 233777
rect 393526 230351 393578 230357
rect 393526 230293 393578 230299
rect 393236 225358 393292 225367
rect 393236 225293 393292 225302
rect 393538 223554 393566 230293
rect 394306 229488 394334 239834
rect 394582 234199 394634 234205
rect 394582 234141 394634 234147
rect 394306 229460 394430 229488
rect 394294 228871 394346 228877
rect 394294 228813 394346 228819
rect 393910 228797 393962 228803
rect 393910 228739 393962 228745
rect 393922 223554 393950 228739
rect 394198 228723 394250 228729
rect 394198 228665 394250 228671
rect 394210 228507 394238 228665
rect 394198 228501 394250 228507
rect 394198 228443 394250 228449
rect 394306 223554 394334 228813
rect 394402 224479 394430 229460
rect 394594 224807 394622 234141
rect 394690 231689 394718 239834
rect 395026 239552 395054 239834
rect 394978 239524 395054 239552
rect 395410 239552 395438 239834
rect 395410 239524 395486 239552
rect 394774 233903 394826 233909
rect 394774 233845 394826 233851
rect 394678 231683 394730 231689
rect 394678 231625 394730 231631
rect 394582 224801 394634 224807
rect 394582 224743 394634 224749
rect 394388 224470 394444 224479
rect 394388 224405 394444 224414
rect 394786 223864 394814 233845
rect 394978 224775 395006 239524
rect 395158 234125 395210 234131
rect 395158 234067 395210 234073
rect 395062 228353 395114 228359
rect 395062 228295 395114 228301
rect 394964 224766 395020 224775
rect 394964 224701 395020 224710
rect 395074 223864 395102 228295
rect 395170 224955 395198 234067
rect 395254 233977 395306 233983
rect 395254 233919 395306 233925
rect 395158 224949 395210 224955
rect 395158 224891 395210 224897
rect 395266 224881 395294 233919
rect 395350 230425 395402 230431
rect 395350 230367 395402 230373
rect 395254 224875 395306 224881
rect 395254 224817 395306 224823
rect 394642 223836 394814 223864
rect 395026 223836 395102 223864
rect 394642 223554 394670 223836
rect 395026 223554 395054 223836
rect 395362 223554 395390 230367
rect 395458 228179 395486 239524
rect 395746 235907 395774 239834
rect 396130 239681 396158 239834
rect 396118 239675 396170 239681
rect 396118 239617 396170 239623
rect 396514 238391 396542 239834
rect 396500 238382 396556 238391
rect 396500 238317 396556 238326
rect 396308 237642 396364 237651
rect 396308 237577 396364 237586
rect 396500 237642 396556 237651
rect 396500 237577 396556 237586
rect 396322 236615 396350 237577
rect 396308 236606 396364 236615
rect 396308 236541 396364 236550
rect 396514 236351 396542 237577
rect 396502 236345 396554 236351
rect 396502 236287 396554 236293
rect 395734 235901 395786 235907
rect 395734 235843 395786 235849
rect 395734 234643 395786 234649
rect 395734 234585 395786 234591
rect 395444 228170 395500 228179
rect 395444 228105 395500 228114
rect 395746 223554 395774 234585
rect 396502 234569 396554 234575
rect 396502 234511 396554 234517
rect 396118 233755 396170 233761
rect 396118 233697 396170 233703
rect 395830 224653 395882 224659
rect 395830 224595 395882 224601
rect 395842 224141 395870 224595
rect 396022 224209 396074 224215
rect 396022 224151 396074 224157
rect 395830 224135 395882 224141
rect 395830 224077 395882 224083
rect 395926 224135 395978 224141
rect 395926 224077 395978 224083
rect 395938 224035 395966 224077
rect 395924 224026 395980 224035
rect 395924 223961 395980 223970
rect 396034 223919 396062 224151
rect 396022 223913 396074 223919
rect 396022 223855 396074 223861
rect 396130 223554 396158 233697
rect 396514 223554 396542 234511
rect 396898 234131 396926 239834
rect 397234 239552 397262 239834
rect 397618 239552 397646 239834
rect 397234 239524 397310 239552
rect 397618 239524 397694 239552
rect 397282 236943 397310 239524
rect 397462 239083 397514 239089
rect 397462 239025 397514 239031
rect 397270 236937 397322 236943
rect 397270 236879 397322 236885
rect 397366 234273 397418 234279
rect 397366 234215 397418 234221
rect 397270 234199 397322 234205
rect 397270 234141 397322 234147
rect 396886 234125 396938 234131
rect 396886 234067 396938 234073
rect 397078 233385 397130 233391
rect 397078 233327 397130 233333
rect 397090 223864 397118 233327
rect 397282 223864 397310 234141
rect 397378 231879 397406 234215
rect 397364 231870 397420 231879
rect 397364 231805 397420 231814
rect 397474 228951 397502 239025
rect 397558 234199 397610 234205
rect 397558 234141 397610 234147
rect 397462 228945 397514 228951
rect 397462 228887 397514 228893
rect 396898 223836 397118 223864
rect 397234 223836 397310 223864
rect 396898 223716 396926 223836
rect 396850 223688 396926 223716
rect 396850 223554 396878 223688
rect 397234 223554 397262 223836
rect 397570 223554 397598 234141
rect 397666 228951 397694 239524
rect 397846 236493 397898 236499
rect 397846 236435 397898 236441
rect 397750 236271 397802 236277
rect 397750 236213 397802 236219
rect 397762 233465 397790 236213
rect 397750 233459 397802 233465
rect 397750 233401 397802 233407
rect 397654 228945 397706 228951
rect 397654 228887 397706 228893
rect 397858 227416 397886 236435
rect 397954 231763 397982 239834
rect 398134 237011 398186 237017
rect 398134 236953 398186 236959
rect 398146 234501 398174 236953
rect 398134 234495 398186 234501
rect 398134 234437 398186 234443
rect 397942 231757 397994 231763
rect 397942 231699 397994 231705
rect 398132 230686 398188 230695
rect 398132 230621 398188 230630
rect 398146 228729 398174 230621
rect 398338 229469 398366 239834
rect 398516 239270 398572 239279
rect 398516 239205 398572 239214
rect 398422 235975 398474 235981
rect 398422 235917 398474 235923
rect 398434 233539 398462 235917
rect 398422 233533 398474 233539
rect 398422 233475 398474 233481
rect 398530 230283 398558 239205
rect 398722 236592 398750 239834
rect 398902 237899 398954 237905
rect 398902 237841 398954 237847
rect 398804 237346 398860 237355
rect 398804 237281 398860 237290
rect 398818 237059 398846 237281
rect 398804 237050 398860 237059
rect 398804 236985 398860 236994
rect 398806 236863 398858 236869
rect 398806 236805 398858 236811
rect 398626 236564 398750 236592
rect 398626 233040 398654 236564
rect 398710 236419 398762 236425
rect 398710 236361 398762 236367
rect 398722 233613 398750 236361
rect 398818 235685 398846 236805
rect 398914 236721 398942 237841
rect 398902 236715 398954 236721
rect 398902 236657 398954 236663
rect 398998 236641 399050 236647
rect 398998 236583 399050 236589
rect 398902 236345 398954 236351
rect 398902 236287 398954 236293
rect 398806 235679 398858 235685
rect 398806 235621 398858 235627
rect 398914 234057 398942 236287
rect 398902 234051 398954 234057
rect 398902 233993 398954 233999
rect 398902 233829 398954 233835
rect 398902 233771 398954 233777
rect 398710 233607 398762 233613
rect 398710 233549 398762 233555
rect 398626 233012 398846 233040
rect 398818 232947 398846 233012
rect 398710 232941 398762 232947
rect 398710 232883 398762 232889
rect 398806 232941 398858 232947
rect 398806 232883 398858 232889
rect 398722 232799 398750 232883
rect 398710 232793 398762 232799
rect 398710 232735 398762 232741
rect 398806 232127 398858 232133
rect 398806 232069 398858 232075
rect 398818 231911 398846 232069
rect 398806 231905 398858 231911
rect 398806 231847 398858 231853
rect 398518 230277 398570 230283
rect 398518 230219 398570 230225
rect 398710 230203 398762 230209
rect 398710 230145 398762 230151
rect 398326 229463 398378 229469
rect 398326 229405 398378 229411
rect 398134 228723 398186 228729
rect 398134 228665 398186 228671
rect 398326 228723 398378 228729
rect 398326 228665 398378 228671
rect 397858 227388 397982 227416
rect 397954 223554 397982 227388
rect 398338 223554 398366 228665
rect 398722 223554 398750 230145
rect 398914 227883 398942 233771
rect 399010 233507 399038 236583
rect 398996 233498 399052 233507
rect 398996 233433 399052 233442
rect 399106 230283 399134 239834
rect 399442 239552 399470 239834
rect 399826 239552 399854 239834
rect 399442 239524 399518 239552
rect 399826 239524 399902 239552
rect 399490 237831 399518 239524
rect 399478 237825 399530 237831
rect 399478 237767 399530 237773
rect 399188 237050 399244 237059
rect 399188 236985 399244 236994
rect 399380 237050 399436 237059
rect 399380 236985 399436 236994
rect 399202 236573 399230 236985
rect 399190 236567 399242 236573
rect 399190 236509 399242 236515
rect 399286 235827 399338 235833
rect 399286 235769 399338 235775
rect 399190 235753 399242 235759
rect 399190 235695 399242 235701
rect 399202 235611 399230 235695
rect 399190 235605 399242 235611
rect 399190 235547 399242 235553
rect 399190 234495 399242 234501
rect 399190 234437 399242 234443
rect 399094 230277 399146 230283
rect 399094 230219 399146 230225
rect 399094 228353 399146 228359
rect 399094 228295 399146 228301
rect 398900 227874 398956 227883
rect 398900 227809 398956 227818
rect 399106 227619 399134 228295
rect 398902 227613 398954 227619
rect 398902 227555 398954 227561
rect 399094 227613 399146 227619
rect 399094 227555 399146 227561
rect 398914 224035 398942 227555
rect 398900 224026 398956 224035
rect 398900 223961 398956 223970
rect 399202 223864 399230 234437
rect 399298 234279 399326 235769
rect 399286 234273 399338 234279
rect 399286 234215 399338 234221
rect 399394 228433 399422 236985
rect 399478 236197 399530 236203
rect 399478 236139 399530 236145
rect 399490 235611 399518 236139
rect 399478 235605 399530 235611
rect 399478 235547 399530 235553
rect 399478 234273 399530 234279
rect 399478 234215 399530 234221
rect 399668 234238 399724 234247
rect 399382 228427 399434 228433
rect 399382 228369 399434 228375
rect 399490 223864 399518 234215
rect 399668 234173 399724 234182
rect 399682 223887 399710 234173
rect 399874 233835 399902 239524
rect 399958 236493 400010 236499
rect 399958 236435 400010 236441
rect 400054 236493 400106 236499
rect 400054 236435 400106 236441
rect 399970 236203 399998 236435
rect 399958 236197 400010 236203
rect 399958 236139 400010 236145
rect 400066 236129 400094 236435
rect 400054 236123 400106 236129
rect 400054 236065 400106 236071
rect 400162 235852 400190 239834
rect 400546 236999 400574 239834
rect 400450 236971 400574 236999
rect 400342 236567 400394 236573
rect 400342 236509 400394 236515
rect 400246 236197 400298 236203
rect 400246 236139 400298 236145
rect 400258 235981 400286 236139
rect 400354 236055 400382 236509
rect 400342 236049 400394 236055
rect 400342 235991 400394 235997
rect 400246 235975 400298 235981
rect 400246 235917 400298 235923
rect 400066 235824 400190 235852
rect 399862 233829 399914 233835
rect 399862 233771 399914 233777
rect 399766 233237 399818 233243
rect 399766 233179 399818 233185
rect 399058 223836 399230 223864
rect 399442 223836 399518 223864
rect 399668 223878 399724 223887
rect 399058 223554 399086 223836
rect 399442 223554 399470 223836
rect 399668 223813 399724 223822
rect 399778 223554 399806 233179
rect 400066 232651 400094 235824
rect 400246 234421 400298 234427
rect 400246 234363 400298 234369
rect 400342 234421 400394 234427
rect 400342 234363 400394 234369
rect 400258 234247 400286 234363
rect 400244 234238 400300 234247
rect 400244 234173 400300 234182
rect 400354 234076 400382 234363
rect 400150 234051 400202 234057
rect 400150 233993 400202 233999
rect 400258 234048 400382 234076
rect 399958 232645 400010 232651
rect 399958 232587 400010 232593
rect 400054 232645 400106 232651
rect 400054 232587 400106 232593
rect 399970 231911 399998 232587
rect 399958 231905 400010 231911
rect 399958 231847 400010 231853
rect 400162 223554 400190 233993
rect 400258 230209 400286 234048
rect 400450 230209 400478 236971
rect 400534 235975 400586 235981
rect 400534 235917 400586 235923
rect 400546 233909 400574 235917
rect 400930 234076 400958 239834
rect 400930 234048 401054 234076
rect 400630 233977 400682 233983
rect 400630 233919 400682 233925
rect 400534 233903 400586 233909
rect 400534 233845 400586 233851
rect 400246 230203 400298 230209
rect 400246 230145 400298 230151
rect 400438 230203 400490 230209
rect 400438 230145 400490 230151
rect 400642 226676 400670 233919
rect 400918 233903 400970 233909
rect 400918 233845 400970 233851
rect 400546 226648 400670 226676
rect 400244 225062 400300 225071
rect 400244 224997 400300 225006
rect 400258 223887 400286 224997
rect 400244 223878 400300 223887
rect 400244 223813 400300 223822
rect 400546 223554 400574 226648
rect 400930 223554 400958 233845
rect 401026 233095 401054 234048
rect 401314 233687 401342 239834
rect 401650 239552 401678 239834
rect 402034 239552 402062 239834
rect 401650 239524 401726 239552
rect 401398 239453 401450 239459
rect 401398 239395 401450 239401
rect 401206 233681 401258 233687
rect 401206 233623 401258 233629
rect 401302 233681 401354 233687
rect 401302 233623 401354 233629
rect 401218 233507 401246 233623
rect 401204 233498 401260 233507
rect 401204 233433 401260 233442
rect 401014 233089 401066 233095
rect 401014 233031 401066 233037
rect 401410 224012 401438 239395
rect 401698 236055 401726 239524
rect 401878 239527 401930 239533
rect 402034 239524 402110 239552
rect 401878 239469 401930 239475
rect 401890 239311 401918 239469
rect 401878 239305 401930 239311
rect 401878 239247 401930 239253
rect 401686 236049 401738 236055
rect 401686 235991 401738 235997
rect 401876 233794 401932 233803
rect 401876 233729 401878 233738
rect 401930 233729 401932 233738
rect 401974 233755 402026 233761
rect 401878 233697 401930 233703
rect 401974 233697 402026 233703
rect 401686 233607 401738 233613
rect 401686 233549 401738 233555
rect 401218 223984 401438 224012
rect 401218 223864 401246 223984
rect 401218 223836 401294 223864
rect 401266 223554 401294 223836
rect 401698 223827 401726 233549
rect 401650 223799 401726 223827
rect 401650 223554 401678 223799
rect 401986 223554 402014 233697
rect 402082 233539 402110 239524
rect 402070 233533 402122 233539
rect 402070 233475 402122 233481
rect 402370 233169 402398 239834
rect 402646 238195 402698 238201
rect 402646 238137 402698 238143
rect 402658 233317 402686 238137
rect 402754 236037 402782 239834
rect 403138 238201 403166 239834
rect 403126 238195 403178 238201
rect 403126 238137 403178 238143
rect 403222 238195 403274 238201
rect 403222 238137 403274 238143
rect 403234 237503 403262 238137
rect 403220 237494 403276 237503
rect 403220 237429 403276 237438
rect 402754 236009 403166 236037
rect 402934 233533 402986 233539
rect 402986 233493 403070 233521
rect 402934 233475 402986 233481
rect 403042 233317 403070 233493
rect 402646 233311 402698 233317
rect 402646 233253 402698 233259
rect 402934 233311 402986 233317
rect 402934 233253 402986 233259
rect 403030 233311 403082 233317
rect 403030 233253 403082 233259
rect 402358 233163 402410 233169
rect 402358 233105 402410 233111
rect 402742 230425 402794 230431
rect 402260 230390 402316 230399
rect 402742 230367 402794 230373
rect 402260 230325 402262 230334
rect 402314 230325 402316 230334
rect 402358 230351 402410 230357
rect 402262 230293 402314 230299
rect 402358 230293 402410 230299
rect 402370 223554 402398 230293
rect 402754 223554 402782 230367
rect 402946 228359 402974 233253
rect 403030 228575 403082 228581
rect 403030 228517 403082 228523
rect 402934 228353 402986 228359
rect 402934 228295 402986 228301
rect 403042 225071 403070 228517
rect 403028 225062 403084 225071
rect 403028 224997 403084 225006
rect 403138 223554 403166 236009
rect 403522 234224 403550 239834
rect 403858 239552 403886 239834
rect 404242 239552 404270 239834
rect 403858 239524 403934 239552
rect 403906 236055 403934 239524
rect 404194 239524 404270 239552
rect 403798 236049 403850 236055
rect 403798 235991 403850 235997
rect 403894 236049 403946 236055
rect 403894 235991 403946 235997
rect 403522 234196 403646 234224
rect 403316 233646 403372 233655
rect 403372 233604 403550 233632
rect 403316 233581 403372 233590
rect 403522 233465 403550 233604
rect 403510 233459 403562 233465
rect 403510 233401 403562 233407
rect 403222 233311 403274 233317
rect 403222 233253 403274 233259
rect 403234 228859 403262 233253
rect 403618 231523 403646 234196
rect 403810 233780 403838 235991
rect 403810 233752 403934 233780
rect 403906 231856 403934 233752
rect 404086 233681 404138 233687
rect 404086 233623 404138 233629
rect 403906 231828 404030 231856
rect 404002 231763 404030 231828
rect 403894 231757 403946 231763
rect 403894 231699 403946 231705
rect 403990 231757 404042 231763
rect 403990 231699 404042 231705
rect 403522 231495 403646 231523
rect 403318 230721 403370 230727
rect 403318 230663 403370 230669
rect 403330 230339 403358 230663
rect 403522 230431 403550 231495
rect 403606 231461 403658 231467
rect 403606 231403 403658 231409
rect 403702 231461 403754 231467
rect 403702 231403 403754 231409
rect 403618 230968 403646 231403
rect 403714 231097 403742 231403
rect 403906 231097 403934 231699
rect 403702 231091 403754 231097
rect 403702 231033 403754 231039
rect 403894 231091 403946 231097
rect 403894 231033 403946 231039
rect 403618 230940 404030 230968
rect 403702 230869 403754 230875
rect 403702 230811 403754 230817
rect 403606 230795 403658 230801
rect 403606 230737 403658 230743
rect 403618 230653 403646 230737
rect 403606 230647 403658 230653
rect 403606 230589 403658 230595
rect 403714 230505 403742 230811
rect 403894 230721 403946 230727
rect 403894 230663 403946 230669
rect 403702 230499 403754 230505
rect 403702 230441 403754 230447
rect 403510 230425 403562 230431
rect 403510 230367 403562 230373
rect 403906 230339 403934 230663
rect 403330 230311 403934 230339
rect 404002 228877 404030 230940
rect 403990 228871 404042 228877
rect 403234 228831 403454 228859
rect 403222 228797 403274 228803
rect 403222 228739 403274 228745
rect 403234 228581 403262 228739
rect 403222 228575 403274 228581
rect 403222 228517 403274 228523
rect 403318 228501 403370 228507
rect 403318 228443 403370 228449
rect 403330 228179 403358 228443
rect 403316 228170 403372 228179
rect 403316 228105 403372 228114
rect 403222 227539 403274 227545
rect 403222 227481 403274 227487
rect 403234 223993 403262 227481
rect 403222 223987 403274 223993
rect 403222 223929 403274 223935
rect 403426 223864 403454 228831
rect 403990 228813 404042 228819
rect 404098 223864 404126 233623
rect 404194 230357 404222 239524
rect 404468 236902 404524 236911
rect 404468 236837 404524 236846
rect 404482 236129 404510 236837
rect 404578 236129 404606 239834
rect 404470 236123 404522 236129
rect 404470 236065 404522 236071
rect 404566 236123 404618 236129
rect 404566 236065 404618 236071
rect 404662 234199 404714 234205
rect 404662 234141 404714 234147
rect 404468 233942 404524 233951
rect 404468 233877 404524 233886
rect 404482 233391 404510 233877
rect 404674 233835 404702 234141
rect 404566 233829 404618 233835
rect 404566 233771 404618 233777
rect 404662 233829 404714 233835
rect 404662 233771 404714 233777
rect 404470 233385 404522 233391
rect 404470 233327 404522 233333
rect 404278 231609 404330 231615
rect 404278 231551 404330 231557
rect 404290 230357 404318 231551
rect 404372 230390 404428 230399
rect 404182 230351 404234 230357
rect 404182 230293 404234 230299
rect 404278 230351 404330 230357
rect 404372 230325 404428 230334
rect 404278 230293 404330 230299
rect 404386 230209 404414 230325
rect 404182 230203 404234 230209
rect 404182 230145 404234 230151
rect 404374 230203 404426 230209
rect 404374 230145 404426 230151
rect 403426 223836 403502 223864
rect 403474 223554 403502 223836
rect 403858 223836 404126 223864
rect 403858 223554 403886 223836
rect 404194 223554 404222 230145
rect 404578 223554 404606 233771
rect 404962 233761 404990 239834
rect 405346 239385 405374 239834
rect 405334 239379 405386 239385
rect 405334 239321 405386 239327
rect 405236 236162 405292 236171
rect 405236 236097 405292 236106
rect 405428 236162 405484 236171
rect 405428 236097 405484 236106
rect 405046 234569 405098 234575
rect 405046 234511 405098 234517
rect 405058 233761 405086 234511
rect 405142 234125 405194 234131
rect 405142 234067 405194 234073
rect 404950 233755 405002 233761
rect 404950 233697 405002 233703
rect 405046 233755 405098 233761
rect 405046 233697 405098 233703
rect 404950 230277 405002 230283
rect 404950 230219 405002 230225
rect 404962 223554 404990 230219
rect 405154 223993 405182 234067
rect 405250 233687 405278 236097
rect 405442 235907 405470 236097
rect 405430 235901 405482 235907
rect 405430 235843 405482 235849
rect 405238 233681 405290 233687
rect 405238 233623 405290 233629
rect 405730 233613 405758 239834
rect 406066 239552 406094 239834
rect 406450 239552 406478 239834
rect 406066 239524 406238 239552
rect 405910 238343 405962 238349
rect 405910 238285 405962 238291
rect 406102 238343 406154 238349
rect 406102 238285 406154 238291
rect 405922 234205 405950 238285
rect 406114 237947 406142 238285
rect 406100 237938 406156 237947
rect 406006 237899 406058 237905
rect 406100 237873 406156 237882
rect 406006 237841 406058 237847
rect 405910 234199 405962 234205
rect 405910 234141 405962 234147
rect 405718 233607 405770 233613
rect 405718 233549 405770 233555
rect 405238 231757 405290 231763
rect 405238 231699 405290 231705
rect 405250 230209 405278 231699
rect 405238 230203 405290 230209
rect 405238 230145 405290 230151
rect 405334 229463 405386 229469
rect 405334 229405 405386 229411
rect 405142 223987 405194 223993
rect 405142 223929 405194 223935
rect 405346 223554 405374 229405
rect 405622 228945 405674 228951
rect 405622 228887 405674 228893
rect 405430 224209 405482 224215
rect 405430 224151 405482 224157
rect 405442 223919 405470 224151
rect 405634 224012 405662 228887
rect 406018 228341 406046 237841
rect 406102 235827 406154 235833
rect 406102 235769 406154 235775
rect 406114 234247 406142 235769
rect 406100 234238 406156 234247
rect 406100 234173 406156 234182
rect 406210 231763 406238 239524
rect 406402 239524 406478 239552
rect 406582 239527 406634 239533
rect 406402 239459 406430 239524
rect 406582 239469 406634 239475
rect 406390 239453 406442 239459
rect 406390 239395 406442 239401
rect 406594 239311 406622 239469
rect 406582 239305 406634 239311
rect 406582 239247 406634 239253
rect 406294 239231 406346 239237
rect 406294 239173 406346 239179
rect 406306 234247 406334 239173
rect 406676 236606 406732 236615
rect 406676 236541 406732 236550
rect 406292 234238 406348 234247
rect 406292 234173 406348 234182
rect 406690 233169 406718 236541
rect 406678 233163 406730 233169
rect 406678 233105 406730 233111
rect 406580 231870 406636 231879
rect 406580 231805 406636 231814
rect 406198 231757 406250 231763
rect 406198 231699 406250 231705
rect 406594 231287 406622 231805
rect 406786 231689 406814 239834
rect 406868 236606 406924 236615
rect 406868 236541 406924 236550
rect 406774 231683 406826 231689
rect 406774 231625 406826 231631
rect 406388 231278 406444 231287
rect 406388 231213 406444 231222
rect 406580 231278 406636 231287
rect 406580 231213 406636 231222
rect 406402 229469 406430 231213
rect 406882 229784 406910 236541
rect 407062 234273 407114 234279
rect 407062 234215 407114 234221
rect 407074 233095 407102 234215
rect 407170 233909 407198 239834
rect 407554 239311 407582 239834
rect 407542 239305 407594 239311
rect 407542 239247 407594 239253
rect 407830 238417 407882 238423
rect 407830 238359 407882 238365
rect 407158 233903 407210 233909
rect 407158 233845 407210 233851
rect 407254 233903 407306 233909
rect 407254 233845 407306 233851
rect 407266 233803 407294 233845
rect 407252 233794 407308 233803
rect 407252 233729 407308 233738
rect 407542 233163 407594 233169
rect 407542 233105 407594 233111
rect 407062 233089 407114 233095
rect 407062 233031 407114 233037
rect 407158 233089 407210 233095
rect 407158 233031 407210 233037
rect 406964 231870 407020 231879
rect 406964 231805 407020 231814
rect 406978 231615 407006 231805
rect 406966 231609 407018 231615
rect 406966 231551 407018 231557
rect 406786 229756 406910 229784
rect 406390 229463 406442 229469
rect 406390 229405 406442 229411
rect 406018 228313 406430 228341
rect 405718 224653 405770 224659
rect 405718 224595 405770 224601
rect 405730 224215 405758 224595
rect 405718 224209 405770 224215
rect 405718 224151 405770 224157
rect 405634 223984 405758 224012
rect 405430 223913 405482 223919
rect 405430 223855 405482 223861
rect 405730 223716 405758 223984
rect 406102 223987 406154 223993
rect 406102 223929 406154 223935
rect 406114 223827 406142 223929
rect 405682 223688 405758 223716
rect 406066 223799 406142 223827
rect 405682 223554 405710 223688
rect 406066 223554 406094 223799
rect 406402 223554 406430 228313
rect 406786 223554 406814 229756
rect 407170 223554 407198 233031
rect 407554 223554 407582 233105
rect 407842 223864 407870 238359
rect 407938 233983 407966 239834
rect 408274 239552 408302 239834
rect 408658 239552 408686 239834
rect 408274 239524 408350 239552
rect 408022 238417 408074 238423
rect 408022 238359 408074 238365
rect 408034 234427 408062 238359
rect 408212 237494 408268 237503
rect 408212 237429 408268 237438
rect 408022 234421 408074 234427
rect 408022 234363 408074 234369
rect 408118 234421 408170 234427
rect 408118 234363 408170 234369
rect 407926 233977 407978 233983
rect 407926 233919 407978 233925
rect 408130 227619 408158 234363
rect 408118 227613 408170 227619
rect 408118 227555 408170 227561
rect 408226 223864 408254 237429
rect 408322 234575 408350 239524
rect 408610 239524 408686 239552
rect 408884 239566 408940 239575
rect 408502 239231 408554 239237
rect 408502 239173 408554 239179
rect 408310 234569 408362 234575
rect 408310 234511 408362 234517
rect 408406 234347 408458 234353
rect 408406 234289 408458 234295
rect 408418 233951 408446 234289
rect 408404 233942 408460 233951
rect 408404 233877 408460 233886
rect 408514 225196 408542 239173
rect 408610 234057 408638 239524
rect 408884 239501 408886 239510
rect 408938 239501 408940 239510
rect 408886 239469 408938 239475
rect 408884 239418 408940 239427
rect 408884 239353 408940 239362
rect 408898 239311 408926 239353
rect 408886 239305 408938 239311
rect 408886 239247 408938 239253
rect 408994 237905 409022 239834
rect 409270 239601 409322 239607
rect 409270 239543 409322 239549
rect 408982 237899 409034 237905
rect 408982 237841 409034 237847
rect 408788 236902 408844 236911
rect 408788 236837 408844 236846
rect 408802 236740 408830 236837
rect 408994 236823 409214 236851
rect 408802 236712 408926 236740
rect 408898 235981 408926 236712
rect 408790 235975 408842 235981
rect 408790 235917 408842 235923
rect 408886 235975 408938 235981
rect 408886 235917 408938 235923
rect 408802 235889 408830 235917
rect 408994 235889 409022 236823
rect 409186 236721 409214 236823
rect 409078 236715 409130 236721
rect 409078 236657 409130 236663
rect 409174 236715 409226 236721
rect 409174 236657 409226 236663
rect 408802 235861 409022 235889
rect 408694 234643 408746 234649
rect 408694 234585 408746 234591
rect 408598 234051 408650 234057
rect 408598 233993 408650 233999
rect 408706 233507 408734 234585
rect 408790 234495 408842 234501
rect 408790 234437 408842 234443
rect 408982 234495 409034 234501
rect 408982 234437 409034 234443
rect 408802 234372 408830 234437
rect 408802 234344 408926 234372
rect 408898 234131 408926 234344
rect 408886 234125 408938 234131
rect 408886 234067 408938 234073
rect 408994 233507 409022 234437
rect 408692 233498 408748 233507
rect 408692 233433 408748 233442
rect 408980 233498 409036 233507
rect 408980 233433 409036 233442
rect 408886 231905 408938 231911
rect 408886 231847 408938 231853
rect 408898 228179 408926 231847
rect 409090 230968 409118 236657
rect 408994 230940 409118 230968
rect 409174 230943 409226 230949
rect 408884 228170 408940 228179
rect 408884 228105 408940 228114
rect 408514 225168 408638 225196
rect 407842 223836 407918 223864
rect 408226 223836 408302 223864
rect 407890 223554 407918 223836
rect 408274 223554 408302 223836
rect 408610 223554 408638 225168
rect 408994 223554 409022 230940
rect 409174 230885 409226 230891
rect 409078 230795 409130 230801
rect 409078 230737 409130 230743
rect 409090 230399 409118 230737
rect 409186 230505 409214 230885
rect 409174 230499 409226 230505
rect 409174 230441 409226 230447
rect 409076 230390 409132 230399
rect 409076 230325 409132 230334
rect 409282 228045 409310 239543
rect 409378 233317 409406 239834
rect 409462 239601 409514 239607
rect 409462 239543 409514 239549
rect 409474 235907 409502 239543
rect 409462 235901 409514 235907
rect 409462 235843 409514 235849
rect 409460 233942 409516 233951
rect 409460 233877 409516 233886
rect 409474 233317 409502 233877
rect 409366 233311 409418 233317
rect 409366 233253 409418 233259
rect 409462 233311 409514 233317
rect 409462 233253 409514 233259
rect 409762 232725 409790 239834
rect 410038 234273 410090 234279
rect 410038 234215 410090 234221
rect 410050 233909 410078 234215
rect 410146 234057 410174 239834
rect 410482 239552 410510 239834
rect 410708 239566 410764 239575
rect 410326 239527 410378 239533
rect 410482 239524 410558 239552
rect 410326 239469 410378 239475
rect 410230 239379 410282 239385
rect 410230 239321 410282 239327
rect 410134 234051 410186 234057
rect 410134 233993 410186 233999
rect 410038 233903 410090 233909
rect 410038 233845 410090 233851
rect 410242 233169 410270 239321
rect 410230 233163 410282 233169
rect 410230 233105 410282 233111
rect 409654 232719 409706 232725
rect 409654 232661 409706 232667
rect 409750 232719 409802 232725
rect 409750 232661 409802 232667
rect 409366 230499 409418 230505
rect 409366 230441 409418 230447
rect 409378 228179 409406 230441
rect 409666 228433 409694 232661
rect 410134 231683 410186 231689
rect 410134 231625 410186 231631
rect 409750 230721 409802 230727
rect 409750 230663 409802 230669
rect 409654 228427 409706 228433
rect 409654 228369 409706 228375
rect 409364 228170 409420 228179
rect 409364 228105 409420 228114
rect 409652 228170 409708 228179
rect 409652 228105 409708 228114
rect 409282 228017 409406 228045
rect 409378 223554 409406 228017
rect 409666 227545 409694 228105
rect 409654 227539 409706 227545
rect 409654 227481 409706 227487
rect 409762 223554 409790 230663
rect 410146 230431 410174 231625
rect 410134 230425 410186 230431
rect 410134 230367 410186 230373
rect 409942 227391 409994 227397
rect 409942 227333 409994 227339
rect 409846 227243 409898 227249
rect 409846 227185 409898 227191
rect 409858 225677 409886 227185
rect 409954 226435 409982 227333
rect 410038 227169 410090 227175
rect 410038 227111 410090 227117
rect 409942 226429 409994 226435
rect 409942 226371 409994 226377
rect 410050 226287 410078 227111
rect 410338 226528 410366 239469
rect 410422 234051 410474 234057
rect 410422 233993 410474 233999
rect 410434 233539 410462 233993
rect 410530 233835 410558 239524
rect 410866 239552 410894 239834
rect 410708 239501 410764 239510
rect 410818 239524 410894 239552
rect 410998 239527 411050 239533
rect 410518 233829 410570 233835
rect 410518 233771 410570 233777
rect 410422 233533 410474 233539
rect 410422 233475 410474 233481
rect 410722 231227 410750 239501
rect 410818 234131 410846 239524
rect 410998 239469 411050 239475
rect 411010 238423 411038 239469
rect 411094 239379 411146 239385
rect 411094 239321 411146 239327
rect 410998 238417 411050 238423
rect 410998 238359 411050 238365
rect 410806 234125 410858 234131
rect 410806 234067 410858 234073
rect 410902 234125 410954 234131
rect 410902 234067 410954 234073
rect 410914 233655 410942 234067
rect 410900 233646 410956 233655
rect 410900 233581 410956 233590
rect 410722 231199 410846 231227
rect 410614 228945 410666 228951
rect 410614 228887 410666 228893
rect 410626 228581 410654 228887
rect 410614 228575 410666 228581
rect 410614 228517 410666 228523
rect 410338 226500 410558 226528
rect 410038 226281 410090 226287
rect 410038 226223 410090 226229
rect 410326 226281 410378 226287
rect 410326 226223 410378 226229
rect 410338 225769 410366 226223
rect 410326 225763 410378 225769
rect 410326 225705 410378 225711
rect 410422 225763 410474 225769
rect 410422 225705 410474 225711
rect 410434 225677 410462 225705
rect 409858 225649 410462 225677
rect 410530 224012 410558 226500
rect 410614 226207 410666 226213
rect 410614 226149 410666 226155
rect 410146 223984 410558 224012
rect 410146 223864 410174 223984
rect 410626 223864 410654 226149
rect 410098 223836 410174 223864
rect 410482 223836 410654 223864
rect 410098 223554 410126 223836
rect 410482 223554 410510 223836
rect 410818 223554 410846 231199
rect 411106 231116 411134 239321
rect 411202 231911 411230 239834
rect 411586 239533 411614 239834
rect 411764 239566 411820 239575
rect 411574 239527 411626 239533
rect 411764 239501 411820 239510
rect 411574 239469 411626 239475
rect 411286 238417 411338 238423
rect 411286 238359 411338 238365
rect 411298 237651 411326 238359
rect 411778 237947 411806 239501
rect 411764 237938 411820 237947
rect 411764 237873 411820 237882
rect 411284 237642 411340 237651
rect 411284 237577 411340 237586
rect 411764 236162 411820 236171
rect 411764 236097 411820 236106
rect 411778 235907 411806 236097
rect 411766 235901 411818 235907
rect 411766 235843 411818 235849
rect 411764 234238 411820 234247
rect 411764 234173 411820 234182
rect 411778 233983 411806 234173
rect 411766 233977 411818 233983
rect 411766 233919 411818 233925
rect 411766 233607 411818 233613
rect 411766 233549 411818 233555
rect 411190 231905 411242 231911
rect 411190 231847 411242 231853
rect 411778 231541 411806 233549
rect 411970 233317 411998 239834
rect 412054 239527 412106 239533
rect 412054 239469 412106 239475
rect 411862 233311 411914 233317
rect 411862 233253 411914 233259
rect 411958 233311 412010 233317
rect 411958 233253 412010 233259
rect 411766 231535 411818 231541
rect 411766 231477 411818 231483
rect 411106 231088 411230 231116
rect 411202 223554 411230 231088
rect 411874 230431 411902 233253
rect 412066 231227 412094 239469
rect 412150 239305 412202 239311
rect 412150 239247 412202 239253
rect 411970 231199 412094 231227
rect 411862 230425 411914 230431
rect 411862 230367 411914 230373
rect 411286 228501 411338 228507
rect 411478 228501 411530 228507
rect 411338 228449 411478 228452
rect 411286 228443 411530 228449
rect 411298 228424 411518 228443
rect 411574 228427 411626 228433
rect 411574 228369 411626 228375
rect 411586 228341 411614 228369
rect 411298 228313 411614 228341
rect 411298 225695 411326 228313
rect 411382 228279 411434 228285
rect 411382 228221 411434 228227
rect 411670 228279 411722 228285
rect 411670 228221 411722 228227
rect 411394 225695 411422 228221
rect 411682 227712 411710 228221
rect 411586 227684 411710 227712
rect 411286 225689 411338 225695
rect 411286 225631 411338 225637
rect 411382 225689 411434 225695
rect 411382 225631 411434 225637
rect 411586 223554 411614 227684
rect 411970 223554 411998 231199
rect 412162 226213 412190 239247
rect 412354 234372 412382 239834
rect 412690 239552 412718 239834
rect 413074 239552 413102 239834
rect 412690 239524 412766 239552
rect 412738 235685 412766 239524
rect 413026 239524 413102 239552
rect 413026 235981 413054 239524
rect 413014 235975 413066 235981
rect 413014 235917 413066 235923
rect 413110 235975 413162 235981
rect 413110 235917 413162 235923
rect 413122 235889 413150 235917
rect 412834 235861 413150 235889
rect 412630 235679 412682 235685
rect 412630 235621 412682 235627
rect 412726 235679 412778 235685
rect 412726 235621 412778 235627
rect 412642 235556 412670 235621
rect 412834 235556 412862 235861
rect 412642 235528 412862 235556
rect 412258 234344 412382 234372
rect 412258 228729 412286 234344
rect 412340 234238 412396 234247
rect 412340 234173 412396 234182
rect 412246 228723 412298 228729
rect 412246 228665 412298 228671
rect 412150 226207 412202 226213
rect 412150 226149 412202 226155
rect 412354 223864 412382 234173
rect 413410 234076 413438 239834
rect 413686 239083 413738 239089
rect 413686 239025 413738 239031
rect 413410 234048 413534 234076
rect 413506 233507 413534 234048
rect 413492 233498 413548 233507
rect 413492 233433 413548 233442
rect 413590 232793 413642 232799
rect 413590 232735 413642 232741
rect 412628 232166 412684 232175
rect 412628 232101 412684 232110
rect 412306 223836 412382 223864
rect 412642 223864 412670 232101
rect 413396 232018 413452 232027
rect 413396 231953 413452 231962
rect 413108 230390 413164 230399
rect 413108 230325 413164 230334
rect 413122 229469 413150 230325
rect 413014 229463 413066 229469
rect 413014 229405 413066 229411
rect 413110 229463 413162 229469
rect 413110 229405 413162 229411
rect 412642 223836 412718 223864
rect 412306 223554 412334 223836
rect 412690 223554 412718 223836
rect 413026 223554 413054 229405
rect 413206 226207 413258 226213
rect 413206 226149 413258 226155
rect 413218 226065 413246 226149
rect 413206 226059 413258 226065
rect 413206 226001 413258 226007
rect 413410 223554 413438 231953
rect 413494 231535 413546 231541
rect 413494 231477 413546 231483
rect 413506 230283 413534 231477
rect 413602 230283 413630 232735
rect 413494 230277 413546 230283
rect 413494 230219 413546 230225
rect 413590 230277 413642 230283
rect 413590 230219 413642 230225
rect 413698 228729 413726 239025
rect 413794 233909 413822 239834
rect 414070 239379 414122 239385
rect 414070 239321 414122 239327
rect 413878 239083 413930 239089
rect 413878 239025 413930 239031
rect 413890 236721 413918 239025
rect 413972 237642 414028 237651
rect 413972 237577 414028 237586
rect 413878 236715 413930 236721
rect 413878 236657 413930 236663
rect 413782 233903 413834 233909
rect 413782 233845 413834 233851
rect 413878 233903 413930 233909
rect 413878 233845 413930 233851
rect 413782 233533 413834 233539
rect 413782 233475 413834 233481
rect 413794 231393 413822 233475
rect 413782 231387 413834 231393
rect 413782 231329 413834 231335
rect 413890 229451 413918 233845
rect 413986 233095 414014 237577
rect 413974 233089 414026 233095
rect 413974 233031 414026 233037
rect 413974 232719 414026 232725
rect 413974 232661 414026 232667
rect 413986 231393 414014 232661
rect 413974 231387 414026 231393
rect 413974 231329 414026 231335
rect 414082 230727 414110 239321
rect 414178 233095 414206 239834
rect 414562 239607 414590 239834
rect 414550 239601 414602 239607
rect 414550 239543 414602 239549
rect 414898 239552 414926 239834
rect 415282 239552 415310 239834
rect 414898 239524 414974 239552
rect 414946 236055 414974 239524
rect 415234 239524 415310 239552
rect 414838 236049 414890 236055
rect 414838 235991 414890 235997
rect 414934 236049 414986 236055
rect 414934 235991 414986 235997
rect 414850 235685 414878 235991
rect 414646 235679 414698 235685
rect 414646 235621 414698 235627
rect 414838 235679 414890 235685
rect 414838 235621 414890 235627
rect 414356 233942 414412 233951
rect 414356 233877 414412 233886
rect 414166 233089 414218 233095
rect 414166 233031 414218 233037
rect 414262 232719 414314 232725
rect 414262 232661 414314 232667
rect 414070 230721 414122 230727
rect 414070 230663 414122 230669
rect 413794 229423 413918 229451
rect 413686 228723 413738 228729
rect 413686 228665 413738 228671
rect 413794 223554 413822 229423
rect 414274 228951 414302 232661
rect 414262 228945 414314 228951
rect 414262 228887 414314 228893
rect 413972 228170 414028 228179
rect 413972 228105 414028 228114
rect 413986 227883 414014 228105
rect 413972 227874 414028 227883
rect 413972 227809 414028 227818
rect 414164 227874 414220 227883
rect 414164 227809 414220 227818
rect 414178 223554 414206 227809
rect 414370 223864 414398 233877
rect 414452 233646 414508 233655
rect 414452 233581 414508 233590
rect 414466 231319 414494 233581
rect 414658 233040 414686 235621
rect 414742 234643 414794 234649
rect 414742 234585 414794 234591
rect 414754 233761 414782 234585
rect 415234 234057 415262 239524
rect 415508 239418 415564 239427
rect 415508 239353 415564 239362
rect 415522 234205 415550 239353
rect 415318 234199 415370 234205
rect 415318 234141 415370 234147
rect 415510 234199 415562 234205
rect 415510 234141 415562 234147
rect 415222 234051 415274 234057
rect 415222 233993 415274 233999
rect 414742 233755 414794 233761
rect 414742 233697 414794 233703
rect 414550 233015 414602 233021
rect 414658 233012 414782 233040
rect 414550 232957 414602 232963
rect 414562 232175 414590 232957
rect 414754 232873 414782 233012
rect 415030 233015 415082 233021
rect 415030 232957 415082 232963
rect 414646 232867 414698 232873
rect 414646 232809 414698 232815
rect 414742 232867 414794 232873
rect 414742 232809 414794 232815
rect 414548 232166 414604 232175
rect 414548 232101 414604 232110
rect 414658 232027 414686 232809
rect 415042 232725 415070 232957
rect 415030 232719 415082 232725
rect 415030 232661 415082 232667
rect 414644 232018 414700 232027
rect 414644 231953 414700 231962
rect 414454 231313 414506 231319
rect 414454 231255 414506 231261
rect 415330 230727 415358 234141
rect 415618 233687 415646 239834
rect 416002 234649 416030 239834
rect 415990 234643 416042 234649
rect 415990 234585 416042 234591
rect 416386 234057 416414 239834
rect 416770 234279 416798 239834
rect 417106 239552 417134 239834
rect 417490 239552 417518 239834
rect 417106 239524 417182 239552
rect 416758 234273 416810 234279
rect 416758 234215 416810 234221
rect 416374 234051 416426 234057
rect 416374 233993 416426 233999
rect 416756 233794 416812 233803
rect 416756 233729 416812 233738
rect 415510 233681 415562 233687
rect 415510 233623 415562 233629
rect 415606 233681 415658 233687
rect 415606 233623 415658 233629
rect 415522 233317 415550 233623
rect 415414 233311 415466 233317
rect 415414 233253 415466 233259
rect 415510 233311 415562 233317
rect 415510 233253 415562 233259
rect 415426 232725 415454 233253
rect 415414 232719 415466 232725
rect 415414 232661 415466 232667
rect 415318 230721 415370 230727
rect 415318 230663 415370 230669
rect 415220 230390 415276 230399
rect 415220 230325 415276 230334
rect 414838 228945 414890 228951
rect 414838 228887 414890 228893
rect 414850 228063 414878 228887
rect 414838 228057 414890 228063
rect 414838 227999 414890 228005
rect 414934 228057 414986 228063
rect 414934 227999 414986 228005
rect 414838 227317 414890 227323
rect 414658 227265 414838 227268
rect 414658 227259 414890 227265
rect 414658 227249 414878 227259
rect 414646 227243 414878 227249
rect 414698 227240 414878 227243
rect 414646 227185 414698 227191
rect 414946 223864 414974 227999
rect 414370 223836 414542 223864
rect 414514 223554 414542 223836
rect 414898 223836 414974 223864
rect 414898 223554 414926 223836
rect 415234 223554 415262 230325
rect 416372 228910 416428 228919
rect 416372 228845 416428 228854
rect 416564 228910 416620 228919
rect 416564 228845 416620 228854
rect 415990 227613 416042 227619
rect 415990 227555 416042 227561
rect 415606 225689 415658 225695
rect 415606 225631 415658 225637
rect 415618 223554 415646 225631
rect 416002 223554 416030 227555
rect 416386 223554 416414 228845
rect 416578 228433 416606 228845
rect 416566 228427 416618 228433
rect 416566 228369 416618 228375
rect 416770 223864 416798 233729
rect 417154 232651 417182 239524
rect 417442 239524 417518 239552
rect 417442 234501 417470 239524
rect 417622 235605 417674 235611
rect 417674 235565 417758 235593
rect 417622 235547 417674 235553
rect 417730 234649 417758 235565
rect 417718 234643 417770 234649
rect 417718 234585 417770 234591
rect 417826 234501 417854 239834
rect 417430 234495 417482 234501
rect 417430 234437 417482 234443
rect 417814 234495 417866 234501
rect 417814 234437 417866 234443
rect 417526 233681 417578 233687
rect 417526 233623 417578 233629
rect 417142 232645 417194 232651
rect 417142 232587 417194 232593
rect 417238 232201 417290 232207
rect 417238 232143 417290 232149
rect 417046 231239 417098 231245
rect 417046 231181 417098 231187
rect 416722 223836 416798 223864
rect 417058 223864 417086 231181
rect 417250 225695 417278 232143
rect 417538 230505 417566 233623
rect 417910 233015 417962 233021
rect 417910 232957 417962 232963
rect 417922 232577 417950 232957
rect 418210 232596 418238 239834
rect 418594 235981 418622 239834
rect 418978 237036 419006 239834
rect 419314 239552 419342 239834
rect 419698 239552 419726 239834
rect 419314 239524 419390 239552
rect 419062 237825 419114 237831
rect 419062 237767 419114 237773
rect 418882 237008 419006 237036
rect 418486 235975 418538 235981
rect 418486 235917 418538 235923
rect 418582 235975 418634 235981
rect 418582 235917 418634 235923
rect 418498 234279 418526 235917
rect 418882 234427 418910 237008
rect 419074 236869 419102 237767
rect 418966 236863 419018 236869
rect 418966 236805 419018 236811
rect 419062 236863 419114 236869
rect 419062 236805 419114 236811
rect 418978 236647 419006 236805
rect 418966 236641 419018 236647
rect 418966 236583 419018 236589
rect 418870 234421 418922 234427
rect 418870 234363 418922 234369
rect 418486 234273 418538 234279
rect 418486 234215 418538 234221
rect 418292 233498 418348 233507
rect 418292 233433 418348 233442
rect 417814 232571 417866 232577
rect 417814 232513 417866 232519
rect 417910 232571 417962 232577
rect 417910 232513 417962 232519
rect 418114 232568 418238 232596
rect 417622 231313 417674 231319
rect 417622 231255 417674 231261
rect 417430 230499 417482 230505
rect 417430 230441 417482 230447
rect 417526 230499 417578 230505
rect 417526 230441 417578 230447
rect 417238 225689 417290 225695
rect 417238 225631 417290 225637
rect 417058 223836 417134 223864
rect 416722 223554 416750 223836
rect 417106 223554 417134 223836
rect 417442 223554 417470 230441
rect 417634 230376 417662 231255
rect 417718 231239 417770 231245
rect 417718 231181 417770 231187
rect 417538 230348 417662 230376
rect 417538 228803 417566 230348
rect 417622 229315 417674 229321
rect 417730 229303 417758 231181
rect 417674 229275 417758 229303
rect 417622 229257 417674 229263
rect 417526 228797 417578 228803
rect 417526 228739 417578 228745
rect 417718 224653 417770 224659
rect 417718 224595 417770 224601
rect 417730 224141 417758 224595
rect 417718 224135 417770 224141
rect 417718 224077 417770 224083
rect 417826 223554 417854 232513
rect 418006 232497 418058 232503
rect 417922 232457 418006 232485
rect 417922 224419 417950 232457
rect 418006 232439 418058 232445
rect 418114 231689 418142 232568
rect 418306 232503 418334 233433
rect 418966 233089 419018 233095
rect 418966 233031 419018 233037
rect 418978 232947 419006 233031
rect 418966 232941 419018 232947
rect 418966 232883 419018 232889
rect 419158 232941 419210 232947
rect 419158 232883 419210 232889
rect 418294 232497 418346 232503
rect 418294 232439 418346 232445
rect 418390 232423 418442 232429
rect 418390 232365 418442 232371
rect 418102 231683 418154 231689
rect 418102 231625 418154 231631
rect 418102 227465 418154 227471
rect 418402 227453 418430 232365
rect 419170 231911 419198 232883
rect 419254 232053 419306 232059
rect 419254 231995 419306 232001
rect 419158 231905 419210 231911
rect 419158 231847 419210 231853
rect 419062 231757 419114 231763
rect 419062 231699 419114 231705
rect 419074 231097 419102 231699
rect 419062 231091 419114 231097
rect 419062 231033 419114 231039
rect 419158 230203 419210 230209
rect 419158 230145 419210 230151
rect 418774 228871 418826 228877
rect 418774 228813 418826 228819
rect 418582 228723 418634 228729
rect 418582 228665 418634 228671
rect 418594 228433 418622 228665
rect 418582 228427 418634 228433
rect 418582 228369 418634 228375
rect 418786 228359 418814 228813
rect 419170 228803 419198 230145
rect 419158 228797 419210 228803
rect 419158 228739 419210 228745
rect 418774 228353 418826 228359
rect 418774 228295 418826 228301
rect 418594 227573 419198 227601
rect 418594 227545 418622 227573
rect 418582 227539 418634 227545
rect 418582 227481 418634 227487
rect 418678 227539 418730 227545
rect 418678 227481 418730 227487
rect 418402 227425 418622 227453
rect 418102 227407 418154 227413
rect 418114 224659 418142 227407
rect 418006 224653 418058 224659
rect 418006 224595 418058 224601
rect 418102 224653 418154 224659
rect 418102 224595 418154 224601
rect 418018 224567 418046 224595
rect 418018 224539 418526 224567
rect 417922 224391 418046 224419
rect 418018 223993 418046 224391
rect 418102 224061 418154 224067
rect 418102 224003 418154 224009
rect 418006 223987 418058 223993
rect 418006 223929 418058 223935
rect 418114 223919 418142 224003
rect 418498 223993 418526 224539
rect 418198 223987 418250 223993
rect 418198 223929 418250 223935
rect 418486 223987 418538 223993
rect 418486 223929 418538 223935
rect 418102 223913 418154 223919
rect 417922 223845 418046 223864
rect 418102 223855 418154 223861
rect 417910 223839 418058 223845
rect 417962 223836 418006 223839
rect 417910 223781 417962 223787
rect 418006 223781 418058 223787
rect 418210 223554 418238 223929
rect 418594 223554 418622 227425
rect 418690 226731 418718 227481
rect 418774 227465 418826 227471
rect 418774 227407 418826 227413
rect 418786 226879 418814 227407
rect 418774 226873 418826 226879
rect 418774 226815 418826 226821
rect 418870 226873 418922 226879
rect 418870 226815 418922 226821
rect 418678 226725 418730 226731
rect 418678 226667 418730 226673
rect 418882 226657 418910 226815
rect 419062 226799 419114 226805
rect 419062 226741 419114 226747
rect 418870 226651 418922 226657
rect 418870 226593 418922 226599
rect 418870 226503 418922 226509
rect 419074 226491 419102 226741
rect 419170 226509 419198 227573
rect 418922 226463 419102 226491
rect 419158 226503 419210 226509
rect 418870 226445 418922 226451
rect 419158 226445 419210 226451
rect 419266 226417 419294 231995
rect 419362 231911 419390 239524
rect 419650 239524 419726 239552
rect 419650 239089 419678 239524
rect 419638 239083 419690 239089
rect 419638 239025 419690 239031
rect 420034 234649 420062 239834
rect 420116 236162 420172 236171
rect 420418 236148 420446 239834
rect 420116 236097 420172 236106
rect 420226 236120 420446 236148
rect 420130 235685 420158 236097
rect 420118 235679 420170 235685
rect 420118 235621 420170 235627
rect 419926 234643 419978 234649
rect 419926 234585 419978 234591
rect 420022 234643 420074 234649
rect 420022 234585 420074 234591
rect 419938 233687 419966 234585
rect 419926 233681 419978 233687
rect 419926 233623 419978 233629
rect 419638 232127 419690 232133
rect 419638 232069 419690 232075
rect 419350 231905 419402 231911
rect 419350 231847 419402 231853
rect 419350 230721 419402 230727
rect 419350 230663 419402 230669
rect 419362 226995 419390 230663
rect 419348 226986 419404 226995
rect 419348 226921 419404 226930
rect 419170 226389 419294 226417
rect 418690 226167 418910 226195
rect 418690 226139 418718 226167
rect 418678 226133 418730 226139
rect 418678 226075 418730 226081
rect 418774 226133 418826 226139
rect 418882 226121 418910 226167
rect 418882 226093 419102 226121
rect 418774 226075 418826 226081
rect 418786 225621 418814 226075
rect 418870 226059 418922 226065
rect 418870 226001 418922 226007
rect 418882 225917 418910 226001
rect 418870 225911 418922 225917
rect 418870 225853 418922 225859
rect 418964 225802 419020 225811
rect 418964 225737 419020 225746
rect 418870 225689 418922 225695
rect 418870 225631 418922 225637
rect 418774 225615 418826 225621
rect 418774 225557 418826 225563
rect 418882 223864 418910 225631
rect 418978 225547 419006 225737
rect 419074 225695 419102 226093
rect 419062 225689 419114 225695
rect 419062 225631 419114 225637
rect 418966 225541 419018 225547
rect 418966 225483 419018 225489
rect 419170 223864 419198 226389
rect 419252 226098 419308 226107
rect 419252 226033 419308 226042
rect 419266 225936 419294 226033
rect 419540 225950 419596 225959
rect 419266 225908 419540 225936
rect 419540 225885 419596 225894
rect 419446 225837 419498 225843
rect 419446 225779 419498 225785
rect 419254 225689 419306 225695
rect 419458 225677 419486 225779
rect 419306 225649 419486 225677
rect 419254 225631 419306 225637
rect 418882 223836 418958 223864
rect 419170 223836 419342 223864
rect 418930 223554 418958 223836
rect 419314 223554 419342 223836
rect 419650 223554 419678 232069
rect 420226 231319 420254 236120
rect 420802 236055 420830 239834
rect 420884 236162 420940 236171
rect 420884 236097 420940 236106
rect 420310 236049 420362 236055
rect 420310 235991 420362 235997
rect 420790 236049 420842 236055
rect 420790 235991 420842 235997
rect 420322 232207 420350 235991
rect 420406 235975 420458 235981
rect 420406 235917 420458 235923
rect 420310 232201 420362 232207
rect 420310 232143 420362 232149
rect 420418 232059 420446 235917
rect 420502 235901 420554 235907
rect 420598 235901 420650 235907
rect 420554 235849 420598 235852
rect 420502 235843 420650 235849
rect 420514 235824 420638 235843
rect 420598 235753 420650 235759
rect 420790 235753 420842 235759
rect 420650 235713 420790 235741
rect 420598 235695 420650 235701
rect 420790 235695 420842 235701
rect 420898 235685 420926 236097
rect 420886 235679 420938 235685
rect 420886 235621 420938 235627
rect 421186 232577 421214 239834
rect 421522 239552 421550 239834
rect 421906 239552 421934 239834
rect 421522 239524 421598 239552
rect 421174 232571 421226 232577
rect 421174 232513 421226 232519
rect 421174 232127 421226 232133
rect 421174 232069 421226 232075
rect 420406 232053 420458 232059
rect 420406 231995 420458 232001
rect 420514 231680 420638 231708
rect 420514 231615 420542 231680
rect 420502 231609 420554 231615
rect 420502 231551 420554 231557
rect 420214 231313 420266 231319
rect 420214 231255 420266 231261
rect 420610 231245 420638 231680
rect 421186 231541 421214 232069
rect 421174 231535 421226 231541
rect 421174 231477 421226 231483
rect 420598 231239 420650 231245
rect 420598 231181 420650 231187
rect 421570 231097 421598 239524
rect 421858 239524 421934 239552
rect 421654 233163 421706 233169
rect 421654 233105 421706 233111
rect 421666 231541 421694 233105
rect 421858 232133 421886 239524
rect 421940 239418 421996 239427
rect 421940 239353 421996 239362
rect 421954 237947 421982 239353
rect 421940 237938 421996 237947
rect 421940 237873 421996 237882
rect 421846 232127 421898 232133
rect 421846 232069 421898 232075
rect 422038 231609 422090 231615
rect 422038 231551 422090 231557
rect 421654 231535 421706 231541
rect 421654 231477 421706 231483
rect 422050 231319 422078 231551
rect 422242 231393 422270 239834
rect 422626 232133 422654 239834
rect 423010 234279 423038 239834
rect 422998 234273 423050 234279
rect 422998 234215 423050 234221
rect 423394 233632 423422 239834
rect 423730 239552 423758 239834
rect 424114 239552 424142 239834
rect 423730 239524 423806 239552
rect 424114 239524 424190 239552
rect 423394 233604 423518 233632
rect 423380 233498 423436 233507
rect 423380 233433 423436 233442
rect 422614 232127 422666 232133
rect 422614 232069 422666 232075
rect 423394 231467 423422 233433
rect 423490 232577 423518 233604
rect 423478 232571 423530 232577
rect 423478 232513 423530 232519
rect 423778 232429 423806 239524
rect 424162 233169 424190 239524
rect 424244 236162 424300 236171
rect 424244 236097 424300 236106
rect 424258 234427 424286 236097
rect 424450 235611 424478 239834
rect 424438 235605 424490 235611
rect 424438 235547 424490 235553
rect 424246 234421 424298 234427
rect 424246 234363 424298 234369
rect 424150 233163 424202 233169
rect 424150 233105 424202 233111
rect 424834 232947 424862 239834
rect 425110 235975 425162 235981
rect 425110 235917 425162 235923
rect 425122 233909 425150 235917
rect 425218 233909 425246 239834
rect 425398 234199 425450 234205
rect 425398 234141 425450 234147
rect 425110 233903 425162 233909
rect 425110 233845 425162 233851
rect 425206 233903 425258 233909
rect 425206 233845 425258 233851
rect 424534 232941 424586 232947
rect 424534 232883 424586 232889
rect 424822 232941 424874 232947
rect 424822 232883 424874 232889
rect 424546 232725 424574 232883
rect 424534 232719 424586 232725
rect 424534 232661 424586 232667
rect 423478 232423 423530 232429
rect 423478 232365 423530 232371
rect 423766 232423 423818 232429
rect 423766 232365 423818 232371
rect 423382 231461 423434 231467
rect 423382 231403 423434 231409
rect 422230 231387 422282 231393
rect 422230 231329 422282 231335
rect 422038 231313 422090 231319
rect 422038 231255 422090 231261
rect 421558 231091 421610 231097
rect 421558 231033 421610 231039
rect 422324 228910 422380 228919
rect 422324 228845 422380 228854
rect 420022 228575 420074 228581
rect 420022 228517 420074 228523
rect 419734 226577 419786 226583
rect 419734 226519 419786 226525
rect 419746 225843 419774 226519
rect 419734 225837 419786 225843
rect 419734 225779 419786 225785
rect 420034 223554 420062 228517
rect 420790 226503 420842 226509
rect 420790 226445 420842 226451
rect 420802 226107 420830 226445
rect 420596 226098 420652 226107
rect 420596 226033 420652 226042
rect 420788 226098 420844 226107
rect 420788 226033 420844 226042
rect 420118 225837 420170 225843
rect 420118 225779 420170 225785
rect 420130 225399 420158 225779
rect 420500 225654 420556 225663
rect 420500 225589 420556 225598
rect 420118 225393 420170 225399
rect 420118 225335 420170 225341
rect 420214 225319 420266 225325
rect 420214 225261 420266 225267
rect 420226 225233 420254 225261
rect 420514 225251 420542 225589
rect 420502 225245 420554 225251
rect 420226 225205 420446 225233
rect 420310 225097 420362 225103
rect 420310 225039 420362 225045
rect 420322 224012 420350 225039
rect 420418 225011 420446 225205
rect 420502 225187 420554 225193
rect 420610 225103 420638 226033
rect 420886 225763 420938 225769
rect 420886 225705 420938 225711
rect 420692 225654 420748 225663
rect 420692 225589 420748 225598
rect 420706 225547 420734 225589
rect 420694 225541 420746 225547
rect 420694 225483 420746 225489
rect 420790 225467 420842 225473
rect 420706 225427 420790 225455
rect 420598 225097 420650 225103
rect 420598 225039 420650 225045
rect 420706 225011 420734 225427
rect 420790 225409 420842 225415
rect 420418 224983 420734 225011
rect 420898 224585 420926 225705
rect 420980 225654 421036 225663
rect 420980 225589 420982 225598
rect 421034 225589 421036 225598
rect 420982 225557 421034 225563
rect 421940 225506 421996 225515
rect 421940 225441 421996 225450
rect 421462 225393 421514 225399
rect 421462 225335 421514 225341
rect 420790 224579 420842 224585
rect 420790 224521 420842 224527
rect 420886 224579 420938 224585
rect 420886 224521 420938 224527
rect 420322 223984 420446 224012
rect 420418 223554 420446 223984
rect 420802 223554 420830 224521
rect 421078 224431 421130 224437
rect 421078 224373 421130 224379
rect 421090 223864 421118 224373
rect 421474 223864 421502 225335
rect 421846 225319 421898 225325
rect 421846 225261 421898 225267
rect 421090 223836 421166 223864
rect 421474 223836 421550 223864
rect 421138 223554 421166 223836
rect 421522 223554 421550 223836
rect 421858 223554 421886 225261
rect 421954 225029 421982 225441
rect 422230 225171 422282 225177
rect 422230 225113 422282 225119
rect 421942 225023 421994 225029
rect 421942 224965 421994 224971
rect 422242 223554 422270 225113
rect 422338 224437 422366 228845
rect 423490 228433 423518 232365
rect 423958 230647 424010 230653
rect 423958 230589 424010 230595
rect 423478 228427 423530 228433
rect 423478 228369 423530 228375
rect 423094 228279 423146 228285
rect 423094 228221 423146 228227
rect 422902 227391 422954 227397
rect 422902 227333 422954 227339
rect 422806 227317 422858 227323
rect 422806 227259 422858 227265
rect 422614 227095 422666 227101
rect 422614 227037 422666 227043
rect 422326 224431 422378 224437
rect 422326 224373 422378 224379
rect 422626 223554 422654 227037
rect 422818 225048 422846 227259
rect 422914 225399 422942 227333
rect 422998 227169 423050 227175
rect 422998 227111 423050 227117
rect 423010 226509 423038 227111
rect 422998 226503 423050 226509
rect 422998 226445 423050 226451
rect 422902 225393 422954 225399
rect 422902 225335 422954 225341
rect 423106 225177 423134 228221
rect 423286 228057 423338 228063
rect 423286 227999 423338 228005
rect 423190 227613 423242 227619
rect 423190 227555 423242 227561
rect 423202 225811 423230 227555
rect 423298 227175 423326 227999
rect 423380 227430 423436 227439
rect 423380 227365 423382 227374
rect 423434 227365 423436 227374
rect 423382 227333 423434 227339
rect 423478 227317 423530 227323
rect 423476 227282 423478 227291
rect 423530 227282 423532 227291
rect 423476 227217 423532 227226
rect 423286 227169 423338 227175
rect 423286 227111 423338 227117
rect 423380 227134 423436 227143
rect 423380 227069 423382 227078
rect 423434 227069 423436 227078
rect 423382 227037 423434 227043
rect 423286 227021 423338 227027
rect 423338 226969 423422 226972
rect 423286 226963 423422 226969
rect 423298 226944 423422 226963
rect 423394 226713 423422 226944
rect 423394 226685 423518 226713
rect 423188 225802 423244 225811
rect 423188 225737 423244 225746
rect 423094 225171 423146 225177
rect 423094 225113 423146 225119
rect 422818 225020 423038 225048
rect 423010 223554 423038 225020
rect 423490 223864 423518 226685
rect 423572 226690 423628 226699
rect 423572 226625 423628 226634
rect 423586 225325 423614 226625
rect 423668 226098 423724 226107
rect 423668 226033 423724 226042
rect 423574 225319 423626 225325
rect 423574 225261 423626 225267
rect 423346 223836 423518 223864
rect 423682 223864 423710 226033
rect 423970 225515 423998 230589
rect 425410 226139 425438 234141
rect 425602 230209 425630 239834
rect 425938 239552 425966 239834
rect 426322 239552 426350 239834
rect 425938 239524 426014 239552
rect 426322 239524 426590 239552
rect 425878 234495 425930 234501
rect 425878 234437 425930 234443
rect 425782 230573 425834 230579
rect 425782 230515 425834 230521
rect 425590 230203 425642 230209
rect 425590 230145 425642 230151
rect 425302 226133 425354 226139
rect 425302 226075 425354 226081
rect 425398 226133 425450 226139
rect 425398 226075 425450 226081
rect 424822 225615 424874 225621
rect 424822 225557 424874 225563
rect 423956 225506 424012 225515
rect 423956 225441 424012 225450
rect 424438 224727 424490 224733
rect 424438 224669 424490 224675
rect 424054 224653 424106 224659
rect 424054 224595 424106 224601
rect 423682 223836 423758 223864
rect 423346 223554 423374 223836
rect 423730 223554 423758 223836
rect 424066 223554 424094 224595
rect 424450 223554 424478 224669
rect 424834 223554 424862 225557
rect 425206 225467 425258 225473
rect 425206 225409 425258 225415
rect 425218 223554 425246 225409
rect 425314 223864 425342 226075
rect 425794 224733 425822 230515
rect 425890 228919 425918 234437
rect 425986 234205 426014 239524
rect 426166 234495 426218 234501
rect 426166 234437 426218 234443
rect 425974 234199 426026 234205
rect 425974 234141 426026 234147
rect 426178 233687 426206 234437
rect 426262 234125 426314 234131
rect 426262 234067 426314 234073
rect 426274 233687 426302 234067
rect 426166 233681 426218 233687
rect 426166 233623 426218 233629
rect 426262 233681 426314 233687
rect 426262 233623 426314 233629
rect 426262 232275 426314 232281
rect 426262 232217 426314 232223
rect 426070 230869 426122 230875
rect 426070 230811 426122 230817
rect 425876 228910 425932 228919
rect 425876 228845 425932 228854
rect 426082 227143 426110 230811
rect 426166 230795 426218 230801
rect 426166 230737 426218 230743
rect 426068 227134 426124 227143
rect 426068 227069 426124 227078
rect 426178 226699 426206 230737
rect 426274 228581 426302 232217
rect 426358 231461 426410 231467
rect 426358 231403 426410 231409
rect 426562 231412 426590 239524
rect 426658 232281 426686 239834
rect 426646 232275 426698 232281
rect 426646 232217 426698 232223
rect 426370 231319 426398 231403
rect 426454 231387 426506 231393
rect 426562 231384 426686 231412
rect 426454 231329 426506 231335
rect 426358 231313 426410 231319
rect 426358 231255 426410 231261
rect 426466 230801 426494 231329
rect 426658 231319 426686 231384
rect 426646 231313 426698 231319
rect 426646 231255 426698 231261
rect 426454 230795 426506 230801
rect 426454 230737 426506 230743
rect 427042 230727 427070 239834
rect 427426 234131 427454 239834
rect 427414 234125 427466 234131
rect 427414 234067 427466 234073
rect 427810 233613 427838 239834
rect 428146 239552 428174 239834
rect 428530 239552 428558 239834
rect 428146 239524 428222 239552
rect 428530 239524 428702 239552
rect 428086 234347 428138 234353
rect 428086 234289 428138 234295
rect 427798 233607 427850 233613
rect 427798 233549 427850 233555
rect 427988 231870 428044 231879
rect 427988 231805 428044 231814
rect 427606 231535 427658 231541
rect 427606 231477 427658 231483
rect 427318 231017 427370 231023
rect 427318 230959 427370 230965
rect 427030 230721 427082 230727
rect 427030 230663 427082 230669
rect 426262 228575 426314 228581
rect 426262 228517 426314 228523
rect 426164 226690 426220 226699
rect 426070 226651 426122 226657
rect 426164 226625 426220 226634
rect 426070 226593 426122 226599
rect 426082 226380 426110 226593
rect 426262 226577 426314 226583
rect 426260 226542 426262 226551
rect 426314 226542 426316 226551
rect 426260 226477 426316 226486
rect 427030 226429 427082 226435
rect 426082 226352 426302 226380
rect 427030 226371 427082 226377
rect 426274 225843 426302 226352
rect 426454 226281 426506 226287
rect 426454 226223 426506 226229
rect 425878 225837 425930 225843
rect 425878 225779 425930 225785
rect 426262 225837 426314 225843
rect 426262 225779 426314 225785
rect 425782 224727 425834 224733
rect 425782 224669 425834 224675
rect 425890 223864 425918 225779
rect 426164 225654 426220 225663
rect 426164 225589 426220 225598
rect 426358 225615 426410 225621
rect 426178 224659 426206 225589
rect 426358 225557 426410 225563
rect 426262 225393 426314 225399
rect 426260 225358 426262 225367
rect 426314 225358 426316 225367
rect 426260 225293 426316 225302
rect 426370 224775 426398 225557
rect 426356 224766 426412 224775
rect 426356 224701 426412 224710
rect 426166 224653 426218 224659
rect 426166 224595 426218 224601
rect 426466 224308 426494 226223
rect 426548 224766 426604 224775
rect 426548 224701 426550 224710
rect 426602 224701 426604 224710
rect 426550 224669 426602 224675
rect 426646 224579 426698 224585
rect 426646 224521 426698 224527
rect 426274 224280 426494 224308
rect 425314 223836 425582 223864
rect 425890 223836 425966 223864
rect 425554 223554 425582 223836
rect 425938 223554 425966 223836
rect 426274 223554 426302 224280
rect 426658 223554 426686 224521
rect 427042 223554 427070 226371
rect 427330 225663 427358 230959
rect 427618 230579 427646 231477
rect 428002 231097 428030 231805
rect 428098 231264 428126 234289
rect 428194 231393 428222 239524
rect 428470 234051 428522 234057
rect 428470 233993 428522 233999
rect 428482 233835 428510 233993
rect 428374 233829 428426 233835
rect 428374 233771 428426 233777
rect 428470 233829 428522 233835
rect 428470 233771 428522 233777
rect 428278 233681 428330 233687
rect 428278 233623 428330 233629
rect 428182 231387 428234 231393
rect 428182 231329 428234 231335
rect 428098 231236 428222 231264
rect 427990 231091 428042 231097
rect 427990 231033 428042 231039
rect 427798 230943 427850 230949
rect 427798 230885 427850 230891
rect 427606 230573 427658 230579
rect 427606 230515 427658 230521
rect 427606 229463 427658 229469
rect 427606 229405 427658 229411
rect 427618 226995 427646 229405
rect 427604 226986 427660 226995
rect 427604 226921 427660 226930
rect 427810 226847 427838 230885
rect 428086 230425 428138 230431
rect 428086 230367 428138 230373
rect 427990 230277 428042 230283
rect 427990 230219 428042 230225
rect 428002 228951 428030 230219
rect 427894 228945 427946 228951
rect 427894 228887 427946 228893
rect 427990 228945 428042 228951
rect 427990 228887 428042 228893
rect 427508 226838 427564 226847
rect 427508 226773 427564 226782
rect 427796 226838 427852 226847
rect 427796 226773 427852 226782
rect 427522 225843 427550 226773
rect 427702 226355 427754 226361
rect 427702 226297 427754 226303
rect 427414 225837 427466 225843
rect 427414 225779 427466 225785
rect 427510 225837 427562 225843
rect 427510 225779 427562 225785
rect 427316 225654 427372 225663
rect 427316 225589 427372 225598
rect 427318 224579 427370 224585
rect 427318 224521 427370 224527
rect 427330 224141 427358 224521
rect 427318 224135 427370 224141
rect 427318 224077 427370 224083
rect 427426 223554 427454 225779
rect 427606 224061 427658 224067
rect 427606 224003 427658 224009
rect 427618 223919 427646 224003
rect 427606 223913 427658 223919
rect 427606 223855 427658 223861
rect 427714 223864 427742 226297
rect 427906 225473 427934 228887
rect 428098 226551 428126 230367
rect 428194 229469 428222 231236
rect 428182 229463 428234 229469
rect 428182 229405 428234 229411
rect 428182 228353 428234 228359
rect 428182 228295 428234 228301
rect 428084 226542 428140 226551
rect 428084 226477 428140 226486
rect 427798 225467 427850 225473
rect 427798 225409 427850 225415
rect 427894 225467 427946 225473
rect 427894 225409 427946 225415
rect 427810 224012 427838 225409
rect 428194 225367 428222 228295
rect 428290 226107 428318 233623
rect 428386 226509 428414 233771
rect 428470 233607 428522 233613
rect 428470 233549 428522 233555
rect 428482 230431 428510 233549
rect 428566 231609 428618 231615
rect 428566 231551 428618 231557
rect 428578 231023 428606 231551
rect 428566 231017 428618 231023
rect 428566 230959 428618 230965
rect 428470 230425 428522 230431
rect 428470 230367 428522 230373
rect 428674 228359 428702 239524
rect 428866 234057 428894 239834
rect 428854 234051 428906 234057
rect 428854 233993 428906 233999
rect 429250 232355 429278 239834
rect 429430 233755 429482 233761
rect 429430 233697 429482 233703
rect 428758 232349 428810 232355
rect 428758 232291 428810 232297
rect 429238 232349 429290 232355
rect 429238 232291 429290 232297
rect 428770 230283 428798 232291
rect 429044 232166 429100 232175
rect 428866 232124 429044 232152
rect 428866 230843 428894 232124
rect 429044 232101 429100 232110
rect 428950 231091 429002 231097
rect 428950 231033 429002 231039
rect 428962 230968 428990 231033
rect 428962 230940 429182 230968
rect 428852 230834 428908 230843
rect 428852 230769 428908 230778
rect 428758 230277 428810 230283
rect 428758 230219 428810 230225
rect 428662 228353 428714 228359
rect 428662 228295 428714 228301
rect 429046 226873 429098 226879
rect 429046 226815 429098 226821
rect 428470 226651 428522 226657
rect 428470 226593 428522 226599
rect 428374 226503 428426 226509
rect 428374 226445 428426 226451
rect 428276 226098 428332 226107
rect 428276 226033 428332 226042
rect 428180 225358 428236 225367
rect 428180 225293 428236 225302
rect 428182 224579 428234 224585
rect 428182 224521 428234 224527
rect 428194 224067 428222 224521
rect 428182 224061 428234 224067
rect 427810 223984 428126 224012
rect 428182 224003 428234 224009
rect 428098 223864 428126 223984
rect 427714 223836 427790 223864
rect 428098 223836 428174 223864
rect 427762 223554 427790 223836
rect 428146 223554 428174 223836
rect 428482 223554 428510 226593
rect 428854 226355 428906 226361
rect 428854 226297 428906 226303
rect 428866 223554 428894 226297
rect 429058 224585 429086 226815
rect 429154 225640 429182 230940
rect 429334 230277 429386 230283
rect 429334 230219 429386 230225
rect 429346 226731 429374 230219
rect 429334 226725 429386 226731
rect 429334 226667 429386 226673
rect 429238 226281 429290 226287
rect 429238 226223 429290 226229
rect 429250 225811 429278 226223
rect 429442 225811 429470 233697
rect 429634 231097 429662 239834
rect 429910 233977 429962 233983
rect 429910 233919 429962 233925
rect 429622 231091 429674 231097
rect 429622 231033 429674 231039
rect 429622 227095 429674 227101
rect 429622 227037 429674 227043
rect 429526 226947 429578 226953
rect 429526 226889 429578 226895
rect 429538 226213 429566 226889
rect 429526 226207 429578 226213
rect 429526 226149 429578 226155
rect 429236 225802 429292 225811
rect 429236 225737 429292 225746
rect 429428 225802 429484 225811
rect 429634 225788 429662 227037
rect 429718 226799 429770 226805
rect 429718 226741 429770 226747
rect 429730 226287 429758 226741
rect 429718 226281 429770 226287
rect 429718 226223 429770 226229
rect 429634 225760 429758 225788
rect 429428 225737 429484 225746
rect 429622 225689 429674 225695
rect 429154 225637 429622 225640
rect 429154 225631 429674 225637
rect 429154 225612 429662 225631
rect 429730 225048 429758 225760
rect 429250 225020 429758 225048
rect 429046 224579 429098 224585
rect 429046 224521 429098 224527
rect 429250 223554 429278 225020
rect 429620 223878 429676 223887
rect 429922 223864 429950 233919
rect 430018 230875 430046 239834
rect 430354 239552 430382 239834
rect 430738 239552 430766 239834
rect 430354 239524 430430 239552
rect 430738 239524 430814 239552
rect 430294 236715 430346 236721
rect 430294 236657 430346 236663
rect 430006 230869 430058 230875
rect 430006 230811 430058 230817
rect 430306 223864 430334 236657
rect 430402 227619 430430 239524
rect 430582 237899 430634 237905
rect 430582 237841 430634 237847
rect 430594 230505 430622 237841
rect 430678 236049 430730 236055
rect 430678 235991 430730 235997
rect 430690 231615 430718 235991
rect 430786 233983 430814 239524
rect 430774 233977 430826 233983
rect 430774 233919 430826 233925
rect 430678 231609 430730 231615
rect 430678 231551 430730 231557
rect 430582 230499 430634 230505
rect 430582 230441 430634 230447
rect 431074 230283 431102 239834
rect 431350 235605 431402 235611
rect 431350 235547 431402 235553
rect 431362 231467 431390 235547
rect 431458 234353 431486 239834
rect 431446 234347 431498 234353
rect 431446 234289 431498 234295
rect 431842 233521 431870 239834
rect 431926 234421 431978 234427
rect 431926 234363 431978 234369
rect 431746 233493 431870 233521
rect 431350 231461 431402 231467
rect 431350 231403 431402 231409
rect 431062 230277 431114 230283
rect 431062 230219 431114 230225
rect 431746 228285 431774 233493
rect 431830 231979 431882 231985
rect 431830 231921 431882 231927
rect 431734 228279 431786 228285
rect 431734 228221 431786 228227
rect 431158 228205 431210 228211
rect 431158 228147 431210 228153
rect 430390 227613 430442 227619
rect 430390 227555 430442 227561
rect 430678 227391 430730 227397
rect 430678 227333 430730 227339
rect 430388 224766 430444 224775
rect 430388 224701 430444 224710
rect 430402 224659 430430 224701
rect 430390 224653 430442 224659
rect 430390 224595 430442 224601
rect 429922 223836 429998 223864
rect 430306 223836 430382 223864
rect 429620 223813 429676 223822
rect 429634 223554 429662 223813
rect 429970 223554 429998 223836
rect 430354 223554 430382 223836
rect 430690 223554 430718 227333
rect 430772 226394 430828 226403
rect 430772 226329 430828 226338
rect 430786 224923 430814 226329
rect 431170 226255 431198 228147
rect 431842 228063 431870 231921
rect 431938 231171 431966 234363
rect 432226 231985 432254 239834
rect 432562 239552 432590 239834
rect 432946 239552 432974 239834
rect 432562 239524 432638 239552
rect 432946 239524 433022 239552
rect 432502 233533 432554 233539
rect 432502 233475 432554 233481
rect 432214 231979 432266 231985
rect 432214 231921 432266 231927
rect 431926 231165 431978 231171
rect 431926 231107 431978 231113
rect 432022 231165 432074 231171
rect 432022 231107 432074 231113
rect 432034 230968 432062 231107
rect 431938 230940 432062 230968
rect 431938 230875 431966 230940
rect 431926 230869 431978 230875
rect 431926 230811 431978 230817
rect 432406 229611 432458 229617
rect 432406 229553 432458 229559
rect 432310 229537 432362 229543
rect 432310 229479 432362 229485
rect 432214 228649 432266 228655
rect 432214 228591 432266 228597
rect 431830 228057 431882 228063
rect 431830 227999 431882 228005
rect 432118 227909 432170 227915
rect 432118 227851 432170 227857
rect 432022 227687 432074 227693
rect 432022 227629 432074 227635
rect 431830 227465 431882 227471
rect 431830 227407 431882 227413
rect 431446 227317 431498 227323
rect 431446 227259 431498 227265
rect 431156 226246 431212 226255
rect 431156 226181 431212 226190
rect 431062 225319 431114 225325
rect 431062 225261 431114 225267
rect 430772 224914 430828 224923
rect 430772 224849 430828 224858
rect 431074 223554 431102 225261
rect 431458 223554 431486 227259
rect 431842 226287 431870 227407
rect 432034 227268 432062 227629
rect 432130 227471 432158 227851
rect 432118 227465 432170 227471
rect 432118 227407 432170 227413
rect 432226 227323 432254 228591
rect 432322 227915 432350 229479
rect 432418 228655 432446 229553
rect 432406 228649 432458 228655
rect 432406 228591 432458 228597
rect 432310 227909 432362 227915
rect 432310 227851 432362 227857
rect 432310 227761 432362 227767
rect 432310 227703 432362 227709
rect 432322 227397 432350 227703
rect 432310 227391 432362 227397
rect 432310 227333 432362 227339
rect 432214 227317 432266 227323
rect 432034 227240 432158 227268
rect 432214 227259 432266 227265
rect 432130 226953 432158 227240
rect 432514 227143 432542 233475
rect 432610 230875 432638 239524
rect 432598 230869 432650 230875
rect 432598 230811 432650 230817
rect 432598 229685 432650 229691
rect 432598 229627 432650 229633
rect 432610 228211 432638 229627
rect 432598 228205 432650 228211
rect 432598 228147 432650 228153
rect 432886 227835 432938 227841
rect 432886 227777 432938 227783
rect 432596 227578 432652 227587
rect 432898 227545 432926 227777
rect 432994 227693 433022 239524
rect 433282 236721 433310 239834
rect 433270 236715 433322 236721
rect 433270 236657 433322 236663
rect 433666 229469 433694 239834
rect 433078 229463 433130 229469
rect 433078 229405 433130 229411
rect 433654 229463 433706 229469
rect 433654 229405 433706 229411
rect 432982 227687 433034 227693
rect 432982 227629 433034 227635
rect 432596 227513 432652 227522
rect 432790 227539 432842 227545
rect 432308 227134 432364 227143
rect 432308 227069 432364 227078
rect 432500 227134 432556 227143
rect 432500 227069 432556 227078
rect 432118 226947 432170 226953
rect 432118 226889 432170 226895
rect 432322 226699 432350 227069
rect 432116 226690 432172 226699
rect 432116 226625 432172 226634
rect 432308 226690 432364 226699
rect 432308 226625 432364 226634
rect 432130 226403 432158 226625
rect 431924 226394 431980 226403
rect 432116 226394 432172 226403
rect 431980 226352 432062 226380
rect 431924 226329 431980 226338
rect 431830 226281 431882 226287
rect 431830 226223 431882 226229
rect 431828 225950 431884 225959
rect 431828 225885 431884 225894
rect 431732 225654 431788 225663
rect 431732 225589 431788 225598
rect 431542 225319 431594 225325
rect 431542 225261 431594 225267
rect 431554 224775 431582 225261
rect 431746 224775 431774 225589
rect 431540 224766 431596 224775
rect 431540 224701 431596 224710
rect 431732 224766 431788 224775
rect 431732 224701 431788 224710
rect 431842 223554 431870 225885
rect 432034 225663 432062 226352
rect 432116 226329 432172 226338
rect 432502 225837 432554 225843
rect 432502 225779 432554 225785
rect 432020 225654 432076 225663
rect 432020 225589 432076 225598
rect 432118 224727 432170 224733
rect 432118 224669 432170 224675
rect 432130 223864 432158 224669
rect 432514 223864 432542 225779
rect 432610 224733 432638 227513
rect 432790 227481 432842 227487
rect 432886 227539 432938 227545
rect 432886 227481 432938 227487
rect 432802 227027 432830 227481
rect 433090 227291 433118 229405
rect 434050 227767 434078 239834
rect 434434 236055 434462 239834
rect 434770 239552 434798 239834
rect 435154 239552 435182 239834
rect 434770 239524 434846 239552
rect 435154 239524 435230 239552
rect 434422 236049 434474 236055
rect 434422 235991 434474 235997
rect 434818 230135 434846 239524
rect 435094 237899 435146 237905
rect 435094 237841 435146 237847
rect 435106 231879 435134 237841
rect 435202 233613 435230 239524
rect 435284 237938 435340 237947
rect 435284 237873 435340 237882
rect 435190 233607 435242 233613
rect 435190 233549 435242 233555
rect 435298 232619 435326 237873
rect 435380 234090 435436 234099
rect 435380 234025 435436 234034
rect 435284 232610 435340 232619
rect 435284 232545 435340 232554
rect 435092 231870 435148 231879
rect 435092 231805 435148 231814
rect 434806 230129 434858 230135
rect 434806 230071 434858 230077
rect 434902 228649 434954 228655
rect 434954 228597 435038 228600
rect 434902 228591 435038 228597
rect 434914 228572 435038 228591
rect 435010 228507 435038 228572
rect 434902 228501 434954 228507
rect 434902 228443 434954 228449
rect 434998 228501 435050 228507
rect 434998 228443 435050 228449
rect 434038 227761 434090 227767
rect 434038 227703 434090 227709
rect 432884 227282 432940 227291
rect 432884 227217 432940 227226
rect 433076 227282 433132 227291
rect 434914 227249 434942 228443
rect 434998 228131 435050 228137
rect 434998 228073 435050 228079
rect 433076 227217 433132 227226
rect 434710 227243 434762 227249
rect 432790 227021 432842 227027
rect 432790 226963 432842 226969
rect 432898 225811 432926 227217
rect 434710 227185 434762 227191
rect 434902 227243 434954 227249
rect 434902 227185 434954 227191
rect 433750 226651 433802 226657
rect 433750 226593 433802 226599
rect 432884 225802 432940 225811
rect 432884 225737 432940 225746
rect 432884 225654 432940 225663
rect 432884 225589 432940 225598
rect 433076 225654 433132 225663
rect 433076 225589 433132 225598
rect 432598 224727 432650 224733
rect 432598 224669 432650 224675
rect 432130 223836 432206 223864
rect 432514 223836 432590 223864
rect 432178 223554 432206 223836
rect 432562 223554 432590 223836
rect 432898 223554 432926 225589
rect 433090 225325 433118 225589
rect 433762 225547 433790 226593
rect 434326 225985 434378 225991
rect 434326 225927 434378 225933
rect 433654 225541 433706 225547
rect 433654 225483 433706 225489
rect 433750 225541 433802 225547
rect 433750 225483 433802 225489
rect 433078 225319 433130 225325
rect 433078 225261 433130 225267
rect 433268 224914 433324 224923
rect 433268 224849 433324 224858
rect 433460 224914 433516 224923
rect 433460 224849 433516 224858
rect 433282 223554 433310 224849
rect 433474 224659 433502 224849
rect 433462 224653 433514 224659
rect 433462 224595 433514 224601
rect 433666 223554 433694 225483
rect 434038 225097 434090 225103
rect 434038 225039 434090 225045
rect 434050 223554 434078 225039
rect 434338 223864 434366 225927
rect 434722 223864 434750 227185
rect 435010 226065 435038 228073
rect 435190 227983 435242 227989
rect 435190 227925 435242 227931
rect 435202 227439 435230 227925
rect 435188 227430 435244 227439
rect 435188 227365 435244 227374
rect 435394 226657 435422 234025
rect 435490 232619 435518 239834
rect 435574 235827 435626 235833
rect 435574 235769 435626 235775
rect 435586 234099 435614 235769
rect 435572 234090 435628 234099
rect 435572 234025 435628 234034
rect 435476 232610 435532 232619
rect 435476 232545 435532 232554
rect 435874 231879 435902 239834
rect 436258 233539 436286 239834
rect 436438 235753 436490 235759
rect 436438 235695 436490 235701
rect 436246 233533 436298 233539
rect 436246 233475 436298 233481
rect 435860 231870 435916 231879
rect 435860 231805 435916 231814
rect 436054 231831 436106 231837
rect 436054 231773 436106 231779
rect 436066 229765 436094 231773
rect 436054 229759 436106 229765
rect 436054 229701 436106 229707
rect 435958 228427 436010 228433
rect 435958 228369 436010 228375
rect 435766 228057 435818 228063
rect 435766 227999 435818 228005
rect 435862 228057 435914 228063
rect 435862 227999 435914 228005
rect 435778 227841 435806 227999
rect 435766 227835 435818 227841
rect 435766 227777 435818 227783
rect 435574 227761 435626 227767
rect 435626 227709 435806 227712
rect 435574 227703 435806 227709
rect 435586 227693 435806 227703
rect 435586 227687 435818 227693
rect 435586 227684 435766 227687
rect 435766 227629 435818 227635
rect 435874 227619 435902 227999
rect 435970 227619 435998 228369
rect 435862 227613 435914 227619
rect 435862 227555 435914 227561
rect 435958 227613 436010 227619
rect 435958 227555 436010 227561
rect 435382 226651 435434 226657
rect 435382 226593 435434 226599
rect 435862 226355 435914 226361
rect 435862 226297 435914 226303
rect 434998 226059 435050 226065
rect 434998 226001 435050 226007
rect 435478 225245 435530 225251
rect 435478 225187 435530 225193
rect 435094 225023 435146 225029
rect 435094 224965 435146 224971
rect 434338 223836 434414 223864
rect 434722 223836 434798 223864
rect 434386 223554 434414 223836
rect 434770 223554 434798 223836
rect 435106 223554 435134 224965
rect 435490 223554 435518 225187
rect 435874 223554 435902 226297
rect 436246 225985 436298 225991
rect 436246 225927 436298 225933
rect 436258 223554 436286 225927
rect 436450 224955 436478 235695
rect 436642 233687 436670 239834
rect 436978 239552 437006 239834
rect 437362 239552 437390 239834
rect 436978 239524 437054 239552
rect 437362 239524 437438 239552
rect 436822 237825 436874 237831
rect 436822 237767 436874 237773
rect 436630 233681 436682 233687
rect 436630 233623 436682 233629
rect 436834 232027 436862 237767
rect 436820 232018 436876 232027
rect 436820 231953 436876 231962
rect 436916 230982 436972 230991
rect 436916 230917 436972 230926
rect 436930 230283 436958 230917
rect 437026 230283 437054 239524
rect 437410 233761 437438 239524
rect 437698 236000 437726 239834
rect 437780 239603 437836 239612
rect 437780 239538 437836 239547
rect 437506 235972 437726 236000
rect 437398 233755 437450 233761
rect 437398 233697 437450 233703
rect 436918 230277 436970 230283
rect 436918 230219 436970 230225
rect 437014 230277 437066 230283
rect 437014 230219 437066 230225
rect 437506 227693 437534 235972
rect 437782 235679 437834 235685
rect 437782 235621 437834 235627
rect 437686 233607 437738 233613
rect 437686 233549 437738 233555
rect 437698 231837 437726 233549
rect 437686 231831 437738 231837
rect 437686 231773 437738 231779
rect 437588 228910 437644 228919
rect 437588 228845 437644 228854
rect 437494 227687 437546 227693
rect 437494 227629 437546 227635
rect 437602 227027 437630 228845
rect 437494 227021 437546 227027
rect 437494 226963 437546 226969
rect 437590 227021 437642 227027
rect 437590 226963 437642 226969
rect 436534 225911 436586 225917
rect 436534 225853 436586 225859
rect 436438 224949 436490 224955
rect 436438 224891 436490 224897
rect 436546 223864 436574 225853
rect 437302 225763 437354 225769
rect 437302 225705 437354 225711
rect 436918 224431 436970 224437
rect 436918 224373 436970 224379
rect 436930 223864 436958 224373
rect 436546 223836 436622 223864
rect 436930 223836 437006 223864
rect 436594 223554 436622 223836
rect 436978 223554 437006 223836
rect 437314 223554 437342 225705
rect 437506 225196 437534 226963
rect 437794 225769 437822 235621
rect 438082 233613 438110 239834
rect 438070 233607 438122 233613
rect 438070 233549 438122 233555
rect 438466 232027 438494 239834
rect 438850 235685 438878 239834
rect 439186 239552 439214 239834
rect 438946 239524 439214 239552
rect 439570 239552 439598 239834
rect 439570 239524 439838 239552
rect 438838 235679 438890 235685
rect 438838 235621 438890 235627
rect 438452 232018 438508 232027
rect 438452 231953 438508 231962
rect 438946 231227 438974 239524
rect 439126 235605 439178 235611
rect 439126 235547 439178 235553
rect 439138 234575 439166 235547
rect 439126 234569 439178 234575
rect 439126 234511 439178 234517
rect 439426 231680 439646 231708
rect 439426 231245 439454 231680
rect 439618 231615 439646 231680
rect 439510 231609 439562 231615
rect 439510 231551 439562 231557
rect 439606 231609 439658 231615
rect 439606 231551 439658 231557
rect 439522 231245 439550 231551
rect 438850 231199 438974 231227
rect 439414 231239 439466 231245
rect 438850 229987 438878 231199
rect 439414 231181 439466 231187
rect 439510 231239 439562 231245
rect 439510 231181 439562 231187
rect 439222 231165 439274 231171
rect 439274 231113 439742 231116
rect 439222 231107 439742 231113
rect 439234 231088 439742 231107
rect 439510 231017 439562 231023
rect 439510 230959 439562 230965
rect 439522 230431 439550 230959
rect 439714 230949 439742 231088
rect 439702 230943 439754 230949
rect 439702 230885 439754 230891
rect 439222 230425 439274 230431
rect 439222 230367 439274 230373
rect 439510 230425 439562 230431
rect 439510 230367 439562 230373
rect 439126 230203 439178 230209
rect 439126 230145 439178 230151
rect 438838 229981 438890 229987
rect 438838 229923 438890 229929
rect 439030 229981 439082 229987
rect 439030 229923 439082 229929
rect 438934 228575 438986 228581
rect 438934 228517 438986 228523
rect 438946 228285 438974 228517
rect 439042 228507 439070 229923
rect 439030 228501 439082 228507
rect 439030 228443 439082 228449
rect 439138 228359 439166 230145
rect 439126 228353 439178 228359
rect 439126 228295 439178 228301
rect 439234 228285 439262 230367
rect 439810 230061 439838 239524
rect 439798 230055 439850 230061
rect 439798 229997 439850 230003
rect 439906 229913 439934 239834
rect 440182 236715 440234 236721
rect 440182 236657 440234 236663
rect 440084 231426 440140 231435
rect 440084 231361 440140 231370
rect 439988 230982 440044 230991
rect 439988 230917 440044 230926
rect 440002 229913 440030 230917
rect 439894 229907 439946 229913
rect 439894 229849 439946 229855
rect 439990 229907 440042 229913
rect 439990 229849 440042 229855
rect 440098 228507 440126 231361
rect 440194 230209 440222 236657
rect 440290 235759 440318 239834
rect 440278 235753 440330 235759
rect 440278 235695 440330 235701
rect 440566 233607 440618 233613
rect 440566 233549 440618 233555
rect 440278 233163 440330 233169
rect 440278 233105 440330 233111
rect 440290 231023 440318 233105
rect 440578 231435 440606 233549
rect 440564 231426 440620 231435
rect 440564 231361 440620 231370
rect 440278 231017 440330 231023
rect 440278 230959 440330 230965
rect 440182 230203 440234 230209
rect 440182 230145 440234 230151
rect 440564 228910 440620 228919
rect 440564 228845 440620 228854
rect 440086 228501 440138 228507
rect 440086 228443 440138 228449
rect 438934 228279 438986 228285
rect 438934 228221 438986 228227
rect 439222 228279 439274 228285
rect 439222 228221 439274 228227
rect 440578 227989 440606 228845
rect 440566 227983 440618 227989
rect 440566 227925 440618 227931
rect 440674 227471 440702 239834
rect 441058 230991 441086 239834
rect 441394 239552 441422 239834
rect 441346 239524 441422 239552
rect 441778 239552 441806 239834
rect 441778 239524 441854 239552
rect 441044 230982 441100 230991
rect 441044 230917 441100 230926
rect 440758 230499 440810 230505
rect 440758 230441 440810 230447
rect 440770 228137 440798 230441
rect 440758 228131 440810 228137
rect 440758 228073 440810 228079
rect 440854 228057 440906 228063
rect 440906 228005 441182 228008
rect 440854 227999 441182 228005
rect 440866 227980 441182 227999
rect 441154 227915 441182 227980
rect 441142 227909 441194 227915
rect 441142 227851 441194 227857
rect 441346 227545 441374 239524
rect 441428 236162 441484 236171
rect 441428 236097 441484 236106
rect 441442 227545 441470 236097
rect 441526 235901 441578 235907
rect 441526 235843 441578 235849
rect 441538 234247 441566 235843
rect 441826 235833 441854 239524
rect 441814 235827 441866 235833
rect 441814 235769 441866 235775
rect 441524 234238 441580 234247
rect 441524 234173 441580 234182
rect 441334 227539 441386 227545
rect 441334 227481 441386 227487
rect 441430 227539 441482 227545
rect 441430 227481 441482 227487
rect 440662 227465 440714 227471
rect 440662 227407 440714 227413
rect 442114 227397 442142 239834
rect 442498 234575 442526 239834
rect 442676 239418 442732 239427
rect 442676 239353 442732 239362
rect 442690 237355 442718 239353
rect 442676 237346 442732 237355
rect 442676 237281 442732 237290
rect 442486 234569 442538 234575
rect 442486 234511 442538 234517
rect 442772 230834 442828 230843
rect 442772 230769 442828 230778
rect 442786 230431 442814 230769
rect 442774 230425 442826 230431
rect 442774 230367 442826 230373
rect 442102 227391 442154 227397
rect 442102 227333 442154 227339
rect 442882 227323 442910 239834
rect 443266 235907 443294 239834
rect 443602 239552 443630 239834
rect 443986 239607 444014 239834
rect 443734 239601 443786 239607
rect 443732 239566 443734 239575
rect 443974 239601 444026 239607
rect 443786 239566 443788 239575
rect 443602 239524 443678 239552
rect 443540 239418 443596 239427
rect 443540 239353 443596 239362
rect 443554 239237 443582 239353
rect 443542 239231 443594 239237
rect 443542 239173 443594 239179
rect 443650 236171 443678 239524
rect 443974 239543 444026 239549
rect 443732 239501 443788 239510
rect 444322 239515 444350 239834
rect 444322 239487 444542 239515
rect 444406 239453 444458 239459
rect 444308 239418 444364 239427
rect 444118 239379 444170 239385
rect 444406 239395 444458 239401
rect 444308 239353 444364 239362
rect 444118 239321 444170 239327
rect 444130 239279 444158 239321
rect 444322 239311 444350 239353
rect 444310 239305 444362 239311
rect 444116 239270 444172 239279
rect 444418 239279 444446 239395
rect 444310 239247 444362 239253
rect 444404 239270 444460 239279
rect 444116 239205 444172 239214
rect 444404 239205 444460 239214
rect 443636 236162 443692 236171
rect 443636 236097 443692 236106
rect 443638 236049 443690 236055
rect 443638 235991 443690 235997
rect 443254 235901 443306 235907
rect 443254 235843 443306 235849
rect 443650 234649 443678 235991
rect 443542 234643 443594 234649
rect 443542 234585 443594 234591
rect 443638 234643 443690 234649
rect 443638 234585 443690 234591
rect 443554 233613 443582 234585
rect 443636 233646 443692 233655
rect 443542 233607 443594 233613
rect 443636 233581 443692 233590
rect 444116 233646 444172 233655
rect 444116 233581 444172 233590
rect 443542 233549 443594 233555
rect 443650 233336 443678 233581
rect 443924 233498 443980 233507
rect 443924 233433 443980 233442
rect 443554 233317 443678 233336
rect 443542 233311 443678 233317
rect 443594 233308 443678 233311
rect 443542 233253 443594 233259
rect 443542 233089 443594 233095
rect 443542 233031 443594 233037
rect 443554 233003 443582 233031
rect 443830 233015 443882 233021
rect 443554 232975 443830 233003
rect 443830 232957 443882 232963
rect 443650 232873 443774 232892
rect 443638 232867 443786 232873
rect 443690 232864 443734 232867
rect 443638 232809 443690 232815
rect 443734 232809 443786 232815
rect 443830 232867 443882 232873
rect 443830 232809 443882 232815
rect 443542 232793 443594 232799
rect 443842 232781 443870 232809
rect 443594 232753 443870 232781
rect 443542 232735 443594 232741
rect 443638 232719 443690 232725
rect 443938 232707 443966 233433
rect 444130 233317 444158 233581
rect 444118 233311 444170 233317
rect 444118 233253 444170 233259
rect 443690 232679 443966 232707
rect 443638 232661 443690 232667
rect 443842 232605 444446 232633
rect 443842 232577 443870 232605
rect 443830 232571 443882 232577
rect 443830 232513 443882 232519
rect 444418 232429 444446 232605
rect 443542 232423 443594 232429
rect 443542 232365 443594 232371
rect 444406 232423 444458 232429
rect 444406 232365 444458 232371
rect 443554 232175 443582 232365
rect 443540 232166 443596 232175
rect 443540 232101 443596 232110
rect 443254 230425 443306 230431
rect 443074 230373 443254 230376
rect 443074 230367 443306 230373
rect 443636 230390 443692 230399
rect 443074 230348 443294 230367
rect 443074 230283 443102 230348
rect 443636 230325 443692 230334
rect 443062 230277 443114 230283
rect 443062 230219 443114 230225
rect 443650 229839 443678 230325
rect 443638 229833 443690 229839
rect 443638 229775 443690 229781
rect 444514 229691 444542 239487
rect 444706 236055 444734 239834
rect 444694 236049 444746 236055
rect 444694 235991 444746 235997
rect 444502 229685 444554 229691
rect 444502 229627 444554 229633
rect 442870 227317 442922 227323
rect 442870 227259 442922 227265
rect 443062 227243 443114 227249
rect 443062 227185 443114 227191
rect 439030 227095 439082 227101
rect 439030 227037 439082 227043
rect 438166 226873 438218 226879
rect 438166 226815 438218 226821
rect 437782 225763 437834 225769
rect 437782 225705 437834 225711
rect 437506 225168 437726 225196
rect 437698 223554 437726 225168
rect 438178 224900 438206 226815
rect 438934 226281 438986 226287
rect 438260 226246 438316 226255
rect 438934 226223 438986 226229
rect 438260 226181 438316 226190
rect 438274 226084 438302 226181
rect 438548 226098 438604 226107
rect 438274 226056 438548 226084
rect 438548 226033 438604 226042
rect 438946 225325 438974 226223
rect 439042 226139 439070 227037
rect 443074 226953 443102 227185
rect 443062 226947 443114 226953
rect 443062 226889 443114 226895
rect 439318 226651 439370 226657
rect 439318 226593 439370 226599
rect 439330 226139 439358 226593
rect 439030 226133 439082 226139
rect 439030 226075 439082 226081
rect 439318 226133 439370 226139
rect 439318 226075 439370 226081
rect 443926 225541 443978 225547
rect 443926 225483 443978 225489
rect 438934 225319 438986 225325
rect 438934 225261 438986 225267
rect 442102 225319 442154 225325
rect 442102 225261 442154 225267
rect 438178 224872 438494 224900
rect 438070 224579 438122 224585
rect 438070 224521 438122 224527
rect 438082 223554 438110 224521
rect 438466 223554 438494 224872
rect 441334 224801 441386 224807
rect 441334 224743 441386 224749
rect 438742 224505 438794 224511
rect 438742 224447 438794 224453
rect 438754 223864 438782 224447
rect 439126 224357 439178 224363
rect 439126 224299 439178 224305
rect 439138 223864 439166 224299
rect 439510 224209 439562 224215
rect 439510 224151 439562 224157
rect 438754 223836 438830 223864
rect 439138 223836 439214 223864
rect 438802 223554 438830 223836
rect 439186 223554 439214 223836
rect 439522 223554 439550 224151
rect 440278 224061 440330 224067
rect 439892 224026 439948 224035
rect 440278 224003 440330 224009
rect 440660 224026 440716 224035
rect 439892 223961 439948 223970
rect 439906 223554 439934 223961
rect 440290 223554 440318 224003
rect 440660 223961 440716 223970
rect 440948 224026 441004 224035
rect 440948 223961 441004 223970
rect 440674 223554 440702 223961
rect 440962 223864 440990 223961
rect 441346 223864 441374 224743
rect 440962 223836 441038 223864
rect 441346 223836 441422 223864
rect 441010 223554 441038 223836
rect 441394 223554 441422 223836
rect 441718 223839 441770 223845
rect 441718 223781 441770 223787
rect 441730 223554 441758 223781
rect 442114 223554 442142 225261
rect 443158 224875 443210 224881
rect 443158 224817 443210 224823
rect 442868 224322 442924 224331
rect 442868 224257 442924 224266
rect 442486 224135 442538 224141
rect 442486 224077 442538 224083
rect 442498 223554 442526 224077
rect 442882 223554 442910 224257
rect 443170 223864 443198 224817
rect 443170 223836 443246 223864
rect 443218 223554 443246 223836
rect 443590 223839 443642 223845
rect 443590 223781 443642 223787
rect 443602 223554 443630 223781
rect 443938 223554 443966 225483
rect 445090 225473 445118 239834
rect 445270 239527 445322 239533
rect 445270 239469 445322 239475
rect 445282 239427 445310 239469
rect 445268 239418 445324 239427
rect 445268 239353 445324 239362
rect 445364 232462 445420 232471
rect 445364 232397 445420 232406
rect 445078 225467 445130 225473
rect 445078 225409 445130 225415
rect 444694 225023 444746 225029
rect 444694 224965 444746 224971
rect 444310 224283 444362 224289
rect 444310 224225 444362 224231
rect 444322 223554 444350 224225
rect 444706 223554 444734 224965
rect 445378 223864 445406 232397
rect 445474 229932 445502 239834
rect 445810 239552 445838 239834
rect 446194 239552 446222 239834
rect 445810 239524 445886 239552
rect 446194 239524 446270 239552
rect 445748 232758 445804 232767
rect 445748 232693 445804 232702
rect 445474 229904 445598 229932
rect 445570 229839 445598 229904
rect 445558 229833 445610 229839
rect 445558 229775 445610 229781
rect 445762 223864 445790 232693
rect 445858 229617 445886 239524
rect 446242 234501 446270 239524
rect 446326 239379 446378 239385
rect 446326 239321 446378 239327
rect 446338 235981 446366 239321
rect 446326 235975 446378 235981
rect 446326 235917 446378 235923
rect 446422 234643 446474 234649
rect 446422 234585 446474 234591
rect 446134 234495 446186 234501
rect 446134 234437 446186 234443
rect 446230 234495 446282 234501
rect 446230 234437 446282 234443
rect 445942 229907 445994 229913
rect 445942 229849 445994 229855
rect 445954 229617 445982 229849
rect 445846 229611 445898 229617
rect 445846 229553 445898 229559
rect 445942 229611 445994 229617
rect 445942 229553 445994 229559
rect 445078 223839 445130 223845
rect 445378 223836 445454 223864
rect 445762 223836 445838 223864
rect 445078 223781 445130 223787
rect 445090 223554 445118 223781
rect 445426 223554 445454 223836
rect 445810 223554 445838 223836
rect 446146 223554 446174 234437
rect 446326 233607 446378 233613
rect 446326 233549 446378 233555
rect 446338 230505 446366 233549
rect 446326 230499 446378 230505
rect 446326 230441 446378 230447
rect 446434 229913 446462 234585
rect 446530 233613 446558 239834
rect 446612 239418 446668 239427
rect 446612 239353 446668 239362
rect 446518 233607 446570 233613
rect 446518 233549 446570 233555
rect 446516 232314 446572 232323
rect 446516 232249 446572 232258
rect 446422 229907 446474 229913
rect 446422 229849 446474 229855
rect 446530 223554 446558 232249
rect 446626 227175 446654 239353
rect 446708 239270 446764 239279
rect 446708 239205 446764 239214
rect 446614 227169 446666 227175
rect 446614 227111 446666 227117
rect 446722 226805 446750 239205
rect 446806 237455 446858 237461
rect 446806 237397 446858 237403
rect 446710 226799 446762 226805
rect 446710 226741 446762 226747
rect 446818 224271 446846 237397
rect 446914 235981 446942 239834
rect 447298 237480 447326 239834
rect 447202 237452 447326 237480
rect 446902 235975 446954 235981
rect 446902 235917 446954 235923
rect 446902 233607 446954 233613
rect 446902 233549 446954 233555
rect 446914 229543 446942 233549
rect 446902 229537 446954 229543
rect 446902 229479 446954 229485
rect 447202 228211 447230 237452
rect 447286 237381 447338 237387
rect 447286 237323 447338 237329
rect 447190 228205 447242 228211
rect 447190 228147 447242 228153
rect 446996 226394 447052 226403
rect 446996 226329 447052 226338
rect 447010 225959 447038 226329
rect 446996 225950 447052 225959
rect 446996 225885 447052 225894
rect 446818 224243 446942 224271
rect 446914 223554 446942 224243
rect 447298 223554 447326 237323
rect 447478 234569 447530 234575
rect 447478 234511 447530 234517
rect 447490 229691 447518 234511
rect 447572 232906 447628 232915
rect 447572 232841 447628 232850
rect 447478 229685 447530 229691
rect 447478 229627 447530 229633
rect 447478 229537 447530 229543
rect 447478 229479 447530 229485
rect 447382 228205 447434 228211
rect 447382 228147 447434 228153
rect 447394 227915 447422 228147
rect 447490 227915 447518 229479
rect 447382 227909 447434 227915
rect 447382 227851 447434 227857
rect 447478 227909 447530 227915
rect 447478 227851 447530 227857
rect 447586 223864 447614 232841
rect 447682 229617 447710 239834
rect 448018 239552 448046 239834
rect 447874 239524 448046 239552
rect 448402 239552 448430 239834
rect 448402 239524 448478 239552
rect 447874 229987 447902 239524
rect 447956 239418 448012 239427
rect 447956 239353 447958 239362
rect 448010 239353 448012 239362
rect 447958 239321 448010 239327
rect 448148 239270 448204 239279
rect 448148 239205 448204 239214
rect 448054 237159 448106 237165
rect 448054 237101 448106 237107
rect 447862 229981 447914 229987
rect 447862 229923 447914 229929
rect 447670 229611 447722 229617
rect 447670 229553 447722 229559
rect 448066 223864 448094 237101
rect 448162 225177 448190 239205
rect 448450 234649 448478 239524
rect 448438 234643 448490 234649
rect 448438 234585 448490 234591
rect 448342 229759 448394 229765
rect 448342 229701 448394 229707
rect 448150 225171 448202 225177
rect 448150 225113 448202 225119
rect 447586 223836 447662 223864
rect 447634 223554 447662 223836
rect 448018 223836 448094 223864
rect 448018 223554 448046 223836
rect 448354 223554 448382 229701
rect 448738 228919 448766 239834
rect 449122 229543 449150 239834
rect 449398 237529 449450 237535
rect 449398 237471 449450 237477
rect 449110 229537 449162 229543
rect 449110 229479 449162 229485
rect 449410 229192 449438 237471
rect 449506 229395 449534 239834
rect 449890 235611 449918 239834
rect 450226 239552 450254 239834
rect 450178 239524 450254 239552
rect 450610 239552 450638 239834
rect 450610 239524 450686 239552
rect 449782 235605 449834 235611
rect 449782 235547 449834 235553
rect 449878 235605 449930 235611
rect 449878 235547 449930 235553
rect 449494 229389 449546 229395
rect 449494 229331 449546 229337
rect 449410 229164 449534 229192
rect 448724 228910 448780 228919
rect 448724 228845 448780 228854
rect 448726 226207 448778 226213
rect 448726 226149 448778 226155
rect 448738 223554 448766 226149
rect 449110 224949 449162 224955
rect 449110 224891 449162 224897
rect 449122 223554 449150 224891
rect 449506 223554 449534 229164
rect 449794 228063 449822 235547
rect 449782 228057 449834 228063
rect 449782 227999 449834 228005
rect 449782 227835 449834 227841
rect 449782 227777 449834 227783
rect 449794 223864 449822 227777
rect 450178 227249 450206 239524
rect 450262 237307 450314 237313
rect 450262 237249 450314 237255
rect 450166 227243 450218 227249
rect 450166 227185 450218 227191
rect 450274 223864 450302 237249
rect 450658 234279 450686 239524
rect 450838 237233 450890 237239
rect 450838 237175 450890 237181
rect 450550 234273 450602 234279
rect 450550 234215 450602 234221
rect 450646 234273 450698 234279
rect 450646 234215 450698 234221
rect 450562 233613 450590 234215
rect 450550 233607 450602 233613
rect 450550 233549 450602 233555
rect 450550 228649 450602 228655
rect 450550 228591 450602 228597
rect 449794 223836 449870 223864
rect 449842 223554 449870 223836
rect 450226 223836 450302 223864
rect 450226 223554 450254 223836
rect 450562 223554 450590 228591
rect 450850 223864 450878 237175
rect 450946 230843 450974 239834
rect 451330 234575 451358 239834
rect 451318 234569 451370 234575
rect 451318 234511 451370 234517
rect 450932 230834 450988 230843
rect 450932 230769 450988 230778
rect 451714 230695 451742 239834
rect 451798 237085 451850 237091
rect 451798 237027 451850 237033
rect 451700 230686 451756 230695
rect 451700 230621 451756 230630
rect 451702 230351 451754 230357
rect 451702 230293 451754 230299
rect 451318 228945 451370 228951
rect 451318 228887 451370 228893
rect 450850 223836 450974 223864
rect 450946 223554 450974 223836
rect 451330 223554 451358 228887
rect 451714 223554 451742 230293
rect 451810 223845 451838 237027
rect 452098 236444 452126 239834
rect 452434 239552 452462 239834
rect 452818 239552 452846 239834
rect 452434 239524 452510 239552
rect 452818 239524 452894 239552
rect 451906 236416 452126 236444
rect 451906 234372 451934 236416
rect 452002 236268 452318 236296
rect 452002 236129 452030 236268
rect 451990 236123 452042 236129
rect 451990 236065 452042 236071
rect 452182 236123 452234 236129
rect 452182 236065 452234 236071
rect 452194 234427 452222 236065
rect 452182 234421 452234 234427
rect 451906 234344 452030 234372
rect 452182 234363 452234 234369
rect 451894 234273 451946 234279
rect 451894 234215 451946 234221
rect 451906 230357 451934 234215
rect 451894 230351 451946 230357
rect 451894 230293 451946 230299
rect 452002 229395 452030 234344
rect 452084 231130 452140 231139
rect 452084 231065 452140 231074
rect 452098 229987 452126 231065
rect 452086 229981 452138 229987
rect 452086 229923 452138 229929
rect 451990 229389 452042 229395
rect 451990 229331 452042 229337
rect 452290 228951 452318 236268
rect 452278 228945 452330 228951
rect 452278 228887 452330 228893
rect 452374 226725 452426 226731
rect 452374 226667 452426 226673
rect 452386 223864 452414 226667
rect 452482 224733 452510 239524
rect 452866 234427 452894 239524
rect 452854 234421 452906 234427
rect 452854 234363 452906 234369
rect 453154 228896 453182 239834
rect 453430 236641 453482 236647
rect 453430 236583 453482 236589
rect 453442 236000 453470 236583
rect 453538 236129 453566 239834
rect 453814 236937 453866 236943
rect 453814 236879 453866 236885
rect 453526 236123 453578 236129
rect 453526 236065 453578 236071
rect 453826 236000 453854 236879
rect 453922 236129 453950 239834
rect 454006 239601 454058 239607
rect 454006 239543 454058 239549
rect 453910 236123 453962 236129
rect 453910 236065 453962 236071
rect 453442 235972 453566 236000
rect 453826 235972 453950 236000
rect 453332 232462 453388 232471
rect 453332 232397 453334 232406
rect 453386 232397 453388 232406
rect 453430 232423 453482 232429
rect 453334 232365 453386 232371
rect 453430 232365 453482 232371
rect 453442 232175 453470 232365
rect 453428 232166 453484 232175
rect 453428 232101 453484 232110
rect 453058 228868 453182 228896
rect 452758 228501 452810 228507
rect 452758 228443 452810 228449
rect 452470 224727 452522 224733
rect 452470 224669 452522 224675
rect 451798 223839 451850 223845
rect 451798 223781 451850 223787
rect 452038 223839 452090 223845
rect 452386 223836 452462 223864
rect 452038 223781 452090 223787
rect 452050 223554 452078 223781
rect 452434 223554 452462 223836
rect 452770 223554 452798 228443
rect 453058 228327 453086 228868
rect 453142 228723 453194 228729
rect 453142 228665 453194 228671
rect 453044 228318 453100 228327
rect 453044 228253 453100 228262
rect 453154 223554 453182 228665
rect 453538 223554 453566 235972
rect 453622 233533 453674 233539
rect 453622 233475 453674 233481
rect 453634 229765 453662 233475
rect 453718 232571 453770 232577
rect 453718 232513 453770 232519
rect 453730 232471 453758 232513
rect 453716 232462 453772 232471
rect 453716 232397 453772 232406
rect 453622 229759 453674 229765
rect 453622 229701 453674 229707
rect 453922 223554 453950 235972
rect 454018 232175 454046 239543
rect 454004 232166 454060 232175
rect 454004 232101 454060 232110
rect 454198 231757 454250 231763
rect 454198 231699 454250 231705
rect 454210 223864 454238 231699
rect 454306 226065 454334 239834
rect 454642 239552 454670 239834
rect 454642 239524 454718 239552
rect 454582 233015 454634 233021
rect 454582 232957 454634 232963
rect 454294 226059 454346 226065
rect 454294 226001 454346 226007
rect 454210 223836 454286 223864
rect 454258 223554 454286 223836
rect 454594 223827 454622 232957
rect 454690 230135 454718 239524
rect 454966 236863 455018 236869
rect 454966 236805 455018 236811
rect 454678 230129 454730 230135
rect 454678 230071 454730 230077
rect 454594 223799 454670 223827
rect 454642 223554 454670 223799
rect 454978 223554 455006 236805
rect 455458 236795 455486 257747
rect 457954 239163 457982 275488
rect 459094 269497 459146 269503
rect 459094 269439 459146 269445
rect 459106 267547 459134 269439
rect 459286 268905 459338 268911
rect 459286 268847 459338 268853
rect 459298 268689 459326 268847
rect 459286 268683 459338 268689
rect 459286 268625 459338 268631
rect 459092 267538 459148 267547
rect 459092 267473 459148 267482
rect 459490 260549 459518 275502
rect 460628 273754 460684 273763
rect 460628 273689 460684 273698
rect 460642 273467 460670 273689
rect 460628 273458 460684 273467
rect 460628 273393 460684 273402
rect 460738 263139 460766 275502
rect 460822 268979 460874 268985
rect 460822 268921 460874 268927
rect 460834 268837 460862 268921
rect 460822 268831 460874 268837
rect 460822 268773 460874 268779
rect 461890 267579 461918 275502
rect 462850 275488 463152 275516
rect 463714 275488 464304 275516
rect 461878 267573 461930 267579
rect 461878 267515 461930 267521
rect 460822 266907 460874 266913
rect 460822 266849 460874 266855
rect 460834 266691 460862 266849
rect 460822 266685 460874 266691
rect 460822 266627 460874 266633
rect 460726 263133 460778 263139
rect 460726 263075 460778 263081
rect 459478 260543 459530 260549
rect 459478 260485 459530 260491
rect 462850 257811 462878 275488
rect 460822 257805 460874 257811
rect 460822 257747 460874 257753
rect 462838 257805 462890 257811
rect 462838 257747 462890 257753
rect 457942 239157 457994 239163
rect 457942 239099 457994 239105
rect 460834 237017 460862 257747
rect 463714 238127 463742 275488
rect 465538 269471 465566 275502
rect 465524 269462 465580 269471
rect 465524 269397 465580 269406
rect 466594 262103 466622 275502
rect 467842 263213 467870 275502
rect 468994 267505 469022 275502
rect 469364 269166 469420 269175
rect 469364 269101 469366 269110
rect 469418 269101 469420 269110
rect 469366 269069 469418 269075
rect 468982 267499 469034 267505
rect 468982 267441 469034 267447
rect 470146 267399 470174 275502
rect 471106 275488 471408 275516
rect 470806 269053 470858 269059
rect 470806 268995 470858 269001
rect 470818 268911 470846 268995
rect 470806 268905 470858 268911
rect 470806 268847 470858 268853
rect 470132 267390 470188 267399
rect 470132 267325 470188 267334
rect 467830 263207 467882 263213
rect 467830 263149 467882 263155
rect 466582 262097 466634 262103
rect 466582 262039 466634 262045
rect 471106 257811 471134 275488
rect 472546 270211 472574 275502
rect 472532 270202 472588 270211
rect 472532 270137 472588 270146
rect 473794 261955 473822 275502
rect 474946 263287 474974 275502
rect 476194 268245 476222 275502
rect 476182 268239 476234 268245
rect 476182 268181 476234 268187
rect 474934 263281 474986 263287
rect 474934 263223 474986 263229
rect 477346 262029 477374 275502
rect 478594 263361 478622 275502
rect 479746 268319 479774 275502
rect 480884 269166 480940 269175
rect 480884 269101 480886 269110
rect 480938 269101 480940 269110
rect 480886 269069 480938 269075
rect 479734 268313 479786 268319
rect 479734 268255 479786 268261
rect 480694 267351 480746 267357
rect 480694 267293 480746 267299
rect 480706 266839 480734 267293
rect 480994 267251 481022 275502
rect 481186 275488 482160 275516
rect 483010 275488 483312 275516
rect 480980 267242 481036 267251
rect 480980 267177 481036 267186
rect 480694 266833 480746 266839
rect 480694 266775 480746 266781
rect 480790 266759 480842 266765
rect 480790 266701 480842 266707
rect 480802 266321 480830 266701
rect 480790 266315 480842 266321
rect 480790 266257 480842 266263
rect 478582 263355 478634 263361
rect 478582 263297 478634 263303
rect 477334 262023 477386 262029
rect 477334 261965 477386 261971
rect 473782 261949 473834 261955
rect 473782 261891 473834 261897
rect 469462 257805 469514 257811
rect 469462 257747 469514 257753
rect 471094 257805 471146 257811
rect 471094 257747 471146 257753
rect 480982 257805 481034 257811
rect 480982 257747 481034 257753
rect 469366 255659 469418 255665
rect 469366 255601 469418 255607
rect 469378 255517 469406 255601
rect 469366 255511 469418 255517
rect 469366 255453 469418 255459
rect 469474 238275 469502 257747
rect 469462 238269 469514 238275
rect 469462 238211 469514 238217
rect 463702 238121 463754 238127
rect 463702 238063 463754 238069
rect 477814 237751 477866 237757
rect 477814 237693 477866 237699
rect 477430 237677 477482 237683
rect 477430 237619 477482 237625
rect 460822 237011 460874 237017
rect 460822 236953 460874 236959
rect 455446 236789 455498 236795
rect 455446 236731 455498 236737
rect 475606 234347 475658 234353
rect 475606 234289 475658 234295
rect 470038 234199 470090 234205
rect 470038 234141 470090 234147
rect 469366 233903 469418 233909
rect 469366 233845 469418 233851
rect 456118 233829 456170 233835
rect 456118 233771 456170 233777
rect 456130 233169 456158 233771
rect 466582 233681 466634 233687
rect 466582 233623 466634 233629
rect 460820 233498 460876 233507
rect 460820 233433 460876 233442
rect 456406 233237 456458 233243
rect 456406 233179 456458 233185
rect 456118 233163 456170 233169
rect 456118 233105 456170 233111
rect 455350 232867 455402 232873
rect 455350 232809 455402 232815
rect 455362 223554 455390 232809
rect 456118 230647 456170 230653
rect 456118 230589 456170 230595
rect 456130 229321 456158 230589
rect 456118 229315 456170 229321
rect 456118 229257 456170 229263
rect 456118 228797 456170 228803
rect 456118 228739 456170 228745
rect 455734 227539 455786 227545
rect 455734 227481 455786 227487
rect 455746 223554 455774 227481
rect 456130 223554 456158 228739
rect 456418 223864 456446 233179
rect 458326 231683 458378 231689
rect 458326 231625 458378 231631
rect 457942 230573 457994 230579
rect 457942 230515 457994 230521
rect 457558 228945 457610 228951
rect 457558 228887 457610 228893
rect 456790 228871 456842 228877
rect 456790 228813 456842 228819
rect 456802 223864 456830 228813
rect 457174 225763 457226 225769
rect 457174 225705 457226 225711
rect 456418 223836 456494 223864
rect 456802 223836 456878 223864
rect 456466 223554 456494 223836
rect 456850 223554 456878 223836
rect 457186 223554 457214 225705
rect 457570 223554 457598 228887
rect 457954 223554 457982 230515
rect 458338 223554 458366 231625
rect 458614 231609 458666 231615
rect 458614 231551 458666 231557
rect 458626 223864 458654 231551
rect 460150 231535 460202 231541
rect 460150 231477 460202 231483
rect 459286 229685 459338 229691
rect 459286 229627 459338 229633
rect 459298 228507 459326 229627
rect 459286 228501 459338 228507
rect 459286 228443 459338 228449
rect 459766 228131 459818 228137
rect 459766 228073 459818 228079
rect 459382 228057 459434 228063
rect 459382 227999 459434 228005
rect 458998 227095 459050 227101
rect 458998 227037 459050 227043
rect 459010 223864 459038 227037
rect 458626 223836 458702 223864
rect 459010 223836 459086 223864
rect 458674 223554 458702 223836
rect 459058 223554 459086 223836
rect 459394 223554 459422 227999
rect 459778 223554 459806 228073
rect 460162 223554 460190 231477
rect 460534 226281 460586 226287
rect 460534 226223 460586 226229
rect 460546 223554 460574 226223
rect 460834 223864 460862 233433
rect 463414 233163 463466 233169
rect 463414 233105 463466 233111
rect 462358 233089 462410 233095
rect 462358 233031 462410 233037
rect 461590 232793 461642 232799
rect 461590 232735 461642 232741
rect 461206 232719 461258 232725
rect 461206 232661 461258 232667
rect 461218 223864 461246 232661
rect 460834 223836 460910 223864
rect 461218 223836 461294 223864
rect 460882 223554 460910 223836
rect 461266 223554 461294 223836
rect 461602 223554 461630 232735
rect 461974 227613 462026 227619
rect 461974 227555 462026 227561
rect 461986 223554 462014 227555
rect 462370 223554 462398 233031
rect 462742 232201 462794 232207
rect 462742 232143 462794 232149
rect 462754 223554 462782 232143
rect 463126 230351 463178 230357
rect 463126 230293 463178 230299
rect 463138 229321 463166 230293
rect 463030 229315 463082 229321
rect 463030 229257 463082 229263
rect 463126 229315 463178 229321
rect 463126 229257 463178 229263
rect 463042 223864 463070 229257
rect 463426 223864 463454 233105
rect 463798 232497 463850 232503
rect 463798 232439 463850 232445
rect 463042 223836 463118 223864
rect 463426 223836 463502 223864
rect 463090 223554 463118 223836
rect 463474 223554 463502 223836
rect 463810 223554 463838 232439
rect 464566 232053 464618 232059
rect 464566 231995 464618 232001
rect 464182 227021 464234 227027
rect 464182 226963 464234 226969
rect 464194 223554 464222 226963
rect 464578 223554 464606 231995
rect 466594 231911 466622 233623
rect 467158 233607 467210 233613
rect 467158 233549 467210 233555
rect 466774 232127 466826 232133
rect 466774 232069 466826 232075
rect 464950 231905 465002 231911
rect 464950 231847 465002 231853
rect 466582 231905 466634 231911
rect 466582 231847 466634 231853
rect 464962 223554 464990 231847
rect 465622 231239 465674 231245
rect 465622 231181 465674 231187
rect 465238 230499 465290 230505
rect 465238 230441 465290 230447
rect 465250 223864 465278 230441
rect 465634 223864 465662 231181
rect 466006 231091 466058 231097
rect 466006 231033 466058 231039
rect 465250 223836 465326 223864
rect 465634 223836 465710 223864
rect 465298 223554 465326 223836
rect 465682 223554 465710 223836
rect 466018 223554 466046 231033
rect 466390 230795 466442 230801
rect 466390 230737 466442 230743
rect 466402 223554 466430 230737
rect 466786 223554 466814 232069
rect 467170 223554 467198 233549
rect 468982 232941 469034 232947
rect 468982 232883 469034 232889
rect 467350 232571 467402 232577
rect 467350 232513 467402 232519
rect 467362 224012 467390 232513
rect 467830 232423 467882 232429
rect 467830 232365 467882 232371
rect 467362 223984 467582 224012
rect 467554 223716 467582 223984
rect 467842 223864 467870 232365
rect 468598 231461 468650 231467
rect 468598 231403 468650 231409
rect 468214 231017 468266 231023
rect 468214 230959 468266 230965
rect 467842 223836 467918 223864
rect 467506 223688 467582 223716
rect 467506 223554 467534 223688
rect 467890 223554 467918 223836
rect 468226 223554 468254 230959
rect 468610 223554 468638 231403
rect 468994 223554 469022 232883
rect 469378 223554 469406 233845
rect 469654 228353 469706 228359
rect 469654 228295 469706 228301
rect 469666 223864 469694 228295
rect 470050 223864 470078 234141
rect 471574 234125 471626 234131
rect 471574 234067 471626 234073
rect 470614 234051 470666 234057
rect 470614 233993 470666 233999
rect 470626 233095 470654 233993
rect 470614 233089 470666 233095
rect 470614 233031 470666 233037
rect 470806 232275 470858 232281
rect 470806 232217 470858 232223
rect 470422 231313 470474 231319
rect 470422 231255 470474 231261
rect 469666 223836 469742 223864
rect 470050 223836 470126 223864
rect 469714 223554 469742 223836
rect 470098 223554 470126 223836
rect 470434 223554 470462 231255
rect 470818 223554 470846 232217
rect 471190 230721 471242 230727
rect 471190 230663 471242 230669
rect 471202 223554 471230 230663
rect 471586 223554 471614 234067
rect 474838 233977 474890 233983
rect 474838 233919 474890 233925
rect 473014 233089 473066 233095
rect 473014 233031 473066 233037
rect 472246 231387 472298 231393
rect 472246 231329 472298 231335
rect 471862 228279 471914 228285
rect 471862 228221 471914 228227
rect 471874 223864 471902 228221
rect 472258 223864 472286 231329
rect 472630 228427 472682 228433
rect 472630 228369 472682 228375
rect 471874 223836 471950 223864
rect 472258 223836 472334 223864
rect 471922 223554 471950 223836
rect 472306 223554 472334 223836
rect 472642 223554 472670 228369
rect 473026 223554 473054 233031
rect 473398 232349 473450 232355
rect 473398 232291 473450 232297
rect 473410 223554 473438 232291
rect 473782 231165 473834 231171
rect 473782 231107 473834 231113
rect 473794 223554 473822 231107
rect 474070 230943 474122 230949
rect 474070 230885 474122 230891
rect 474082 223864 474110 230885
rect 474454 228205 474506 228211
rect 474454 228147 474506 228153
rect 474466 223864 474494 228147
rect 474082 223836 474158 223864
rect 474466 223836 474542 223864
rect 474130 223554 474158 223836
rect 474514 223554 474542 223836
rect 474850 223554 474878 233919
rect 475126 233755 475178 233761
rect 475126 233697 475178 233703
rect 475138 232059 475166 233697
rect 475126 232053 475178 232059
rect 475126 231995 475178 232001
rect 475222 227909 475274 227915
rect 475222 227851 475274 227857
rect 475234 223554 475262 227851
rect 475618 223554 475646 234289
rect 476278 231979 476330 231985
rect 476278 231921 476330 231927
rect 475990 228575 476042 228581
rect 475990 228517 476042 228523
rect 476002 223554 476030 228517
rect 476290 223864 476318 231921
rect 476662 230869 476714 230875
rect 476662 230811 476714 230817
rect 476674 223864 476702 230811
rect 477046 227983 477098 227989
rect 477046 227925 477098 227931
rect 476290 223836 476366 223864
rect 476674 223836 476750 223864
rect 476338 223554 476366 223836
rect 476722 223554 476750 223836
rect 477058 223554 477086 227925
rect 477442 223554 477470 237619
rect 477526 229167 477578 229173
rect 477526 229109 477578 229115
rect 477538 229025 477566 229109
rect 477526 229019 477578 229025
rect 477526 228961 477578 228967
rect 477826 223554 477854 237693
rect 478198 237603 478250 237609
rect 478198 237545 478250 237551
rect 478210 223554 478238 237545
rect 479638 236567 479690 236573
rect 479638 236509 479690 236515
rect 479254 236493 479306 236499
rect 479254 236435 479306 236441
rect 478870 236419 478922 236425
rect 478870 236361 478922 236367
rect 478486 236345 478538 236351
rect 478486 236287 478538 236293
rect 478498 223864 478526 236287
rect 478882 223864 478910 236361
rect 478498 223836 478574 223864
rect 478882 223836 478958 223864
rect 478546 223554 478574 223836
rect 478930 223554 478958 223836
rect 479266 223554 479294 236435
rect 479446 229463 479498 229469
rect 479446 229405 479498 229411
rect 479458 229247 479486 229405
rect 479446 229241 479498 229247
rect 479446 229183 479498 229189
rect 479650 223554 479678 236509
rect 480692 234978 480748 234987
rect 480692 234913 480748 234922
rect 480020 234830 480076 234839
rect 480020 234765 480076 234774
rect 480034 223554 480062 234765
rect 480406 229981 480458 229987
rect 480406 229923 480458 229929
rect 480418 223554 480446 229923
rect 480706 223864 480734 234913
rect 480994 224183 481022 257747
rect 481186 238497 481214 275488
rect 483010 257811 483038 275488
rect 484450 261881 484478 275502
rect 485206 266907 485258 266913
rect 485206 266849 485258 266855
rect 485218 266247 485246 266849
rect 485206 266241 485258 266247
rect 485206 266183 485258 266189
rect 485602 263435 485630 275502
rect 486850 268393 486878 275502
rect 487042 275488 488016 275516
rect 488962 275488 489264 275516
rect 489634 275488 490416 275516
rect 486838 268387 486890 268393
rect 486838 268329 486890 268335
rect 485590 263429 485642 263435
rect 485590 263371 485642 263377
rect 484438 261875 484490 261881
rect 484438 261817 484490 261823
rect 482998 257805 483050 257811
rect 482998 257747 483050 257753
rect 486838 257805 486890 257811
rect 486838 257747 486890 257753
rect 486850 238571 486878 257747
rect 486838 238565 486890 238571
rect 486838 238507 486890 238513
rect 481174 238491 481226 238497
rect 481174 238433 481226 238439
rect 485494 237973 485546 237979
rect 485494 237915 485546 237921
rect 482614 236271 482666 236277
rect 482614 236213 482666 236219
rect 481076 234682 481132 234691
rect 481076 234617 481132 234626
rect 480980 224174 481036 224183
rect 480980 224109 481036 224118
rect 481090 223864 481118 234617
rect 481846 233459 481898 233465
rect 481846 233401 481898 233407
rect 481462 233311 481514 233317
rect 481462 233253 481514 233259
rect 480706 223836 480782 223864
rect 481090 223836 481166 223864
rect 480754 223554 480782 223836
rect 481138 223554 481166 223836
rect 481474 223554 481502 233253
rect 481858 223554 481886 233401
rect 482230 233385 482282 233391
rect 482230 233327 482282 233333
rect 482242 223554 482270 233327
rect 482626 223554 482654 236213
rect 482902 236197 482954 236203
rect 482902 236139 482954 236145
rect 482914 223864 482942 236139
rect 485108 235422 485164 235431
rect 485108 235357 485164 235366
rect 483668 235274 483724 235283
rect 483668 235209 483724 235218
rect 483284 228170 483340 228179
rect 483284 228105 483340 228114
rect 483298 223864 483326 228105
rect 482914 223836 482990 223864
rect 483298 223836 483374 223864
rect 482962 223554 482990 223836
rect 483346 223554 483374 223836
rect 483682 223554 483710 235209
rect 484436 235126 484492 235135
rect 484436 235061 484492 235070
rect 483862 230203 483914 230209
rect 483862 230145 483914 230151
rect 483874 223845 483902 230145
rect 484054 226133 484106 226139
rect 484054 226075 484106 226081
rect 483862 223839 483914 223845
rect 483862 223781 483914 223787
rect 484066 223554 484094 226075
rect 484450 223554 484478 235061
rect 484820 228466 484876 228475
rect 484820 228401 484876 228410
rect 484834 223554 484862 228401
rect 485122 223864 485150 235357
rect 485506 223864 485534 237915
rect 487042 236467 487070 275488
rect 488962 257811 488990 275488
rect 488950 257805 489002 257811
rect 488950 257747 489002 257753
rect 489634 237628 489662 275488
rect 489718 269127 489770 269133
rect 489718 269069 489770 269075
rect 489730 268911 489758 269069
rect 489718 268905 489770 268911
rect 489718 268847 489770 268853
rect 489814 267351 489866 267357
rect 489814 267293 489866 267299
rect 489826 266839 489854 267293
rect 489814 266833 489866 266839
rect 489814 266775 489866 266781
rect 489718 266759 489770 266765
rect 489718 266701 489770 266707
rect 489730 266321 489758 266701
rect 489718 266315 489770 266321
rect 489718 266257 489770 266263
rect 491650 261807 491678 275502
rect 492802 263509 492830 275502
rect 494050 268467 494078 275502
rect 494818 275488 495216 275516
rect 495490 275488 496464 275516
rect 497314 275488 497616 275516
rect 494038 268461 494090 268467
rect 494038 268403 494090 268409
rect 492790 263503 492842 263509
rect 492790 263445 492842 263451
rect 491638 261801 491690 261807
rect 491638 261743 491690 261749
rect 494818 257811 494846 275488
rect 495286 266907 495338 266913
rect 495286 266849 495338 266855
rect 495298 266247 495326 266849
rect 495286 266241 495338 266247
rect 495286 266183 495338 266189
rect 492694 257805 492746 257811
rect 492694 257747 492746 257753
rect 494806 257805 494858 257811
rect 494806 257747 494858 257753
rect 495382 257805 495434 257811
rect 495382 257747 495434 257753
rect 490966 255733 491018 255739
rect 490966 255675 491018 255681
rect 490978 255591 491006 255675
rect 490966 255585 491018 255591
rect 490966 255527 491018 255533
rect 489634 237600 489758 237628
rect 487028 236458 487084 236467
rect 487028 236393 487084 236402
rect 486644 236014 486700 236023
rect 486644 235949 486700 235958
rect 485876 235570 485932 235579
rect 485876 235505 485932 235514
rect 485122 223836 485198 223864
rect 485506 223836 485582 223864
rect 485170 223554 485198 223836
rect 485554 223554 485582 223836
rect 485890 223554 485918 235505
rect 486260 229206 486316 229215
rect 486260 229141 486316 229150
rect 486274 223554 486302 229141
rect 486658 223554 486686 235949
rect 488084 235866 488140 235875
rect 488084 235801 488140 235810
rect 487316 235718 487372 235727
rect 487316 235653 487372 235662
rect 487028 229354 487084 229363
rect 487028 229289 487084 229298
rect 487042 223554 487070 229289
rect 487330 223864 487358 235653
rect 487700 229058 487756 229067
rect 487700 228993 487756 229002
rect 487714 223864 487742 228993
rect 487330 223836 487406 223864
rect 487714 223836 487790 223864
rect 487378 223554 487406 223836
rect 487762 223554 487790 223836
rect 488098 223554 488126 235801
rect 488854 235087 488906 235093
rect 488854 235029 488906 235035
rect 488468 230538 488524 230547
rect 488468 230473 488524 230482
rect 488482 223554 488510 230473
rect 488866 223554 488894 235029
rect 489620 231278 489676 231287
rect 489620 231213 489676 231222
rect 489238 229019 489290 229025
rect 489238 228961 489290 228967
rect 489250 223554 489278 228961
rect 489634 223864 489662 231213
rect 489730 225399 489758 237600
rect 492706 236319 492734 257747
rect 495286 256177 495338 256183
rect 495286 256119 495338 256125
rect 495298 253593 495326 256119
rect 495286 253587 495338 253593
rect 495286 253529 495338 253535
rect 492692 236310 492748 236319
rect 492692 236245 492748 236254
rect 494998 236049 495050 236055
rect 494998 235991 495050 235997
rect 493750 235901 493802 235907
rect 493750 235843 493802 235849
rect 493558 235827 493610 235833
rect 493558 235769 493610 235775
rect 491734 235531 491786 235537
rect 491734 235473 491786 235479
rect 491062 235161 491114 235167
rect 491062 235103 491114 235109
rect 490294 234865 490346 234871
rect 490294 234807 490346 234813
rect 489910 229167 489962 229173
rect 489910 229109 489962 229115
rect 489718 225393 489770 225399
rect 489718 225335 489770 225341
rect 489586 223836 489662 223864
rect 489922 223864 489950 229109
rect 489922 223836 489998 223864
rect 489586 223554 489614 223836
rect 489970 223554 489998 223836
rect 490306 223554 490334 234807
rect 490678 228945 490730 228951
rect 490678 228887 490730 228893
rect 490690 223554 490718 228887
rect 491074 223554 491102 235103
rect 491446 229093 491498 229099
rect 491446 229035 491498 229041
rect 491458 223554 491486 229035
rect 491746 223864 491774 235473
rect 493270 235013 493322 235019
rect 493270 234955 493322 234961
rect 492502 234717 492554 234723
rect 492502 234659 492554 234665
rect 492116 231574 492172 231583
rect 492116 231509 492172 231518
rect 492130 223864 492158 231509
rect 491746 223836 491822 223864
rect 492130 223836 492206 223864
rect 491794 223554 491822 223836
rect 492178 223554 492206 223836
rect 492514 223554 492542 234659
rect 492884 229946 492940 229955
rect 492884 229881 492940 229890
rect 492898 223554 492926 229881
rect 493282 223554 493310 234955
rect 493570 229173 493598 235769
rect 493558 229167 493610 229173
rect 493558 229109 493610 229115
rect 493762 228803 493790 235843
rect 494806 235753 494858 235759
rect 494806 235695 494858 235701
rect 494422 235679 494474 235685
rect 494422 235621 494474 235627
rect 494038 235235 494090 235241
rect 494038 235177 494090 235183
rect 493942 234495 493994 234501
rect 493942 234437 493994 234443
rect 493954 229099 493982 234437
rect 493942 229093 493994 229099
rect 493942 229035 493994 229041
rect 493750 228797 493802 228803
rect 493652 228762 493708 228771
rect 493750 228739 493802 228745
rect 493652 228697 493708 228706
rect 493666 223554 493694 228697
rect 494050 223864 494078 235177
rect 494324 230094 494380 230103
rect 494324 230029 494380 230038
rect 494002 223836 494078 223864
rect 494338 223864 494366 230029
rect 494434 229987 494462 235621
rect 494710 235383 494762 235389
rect 494710 235325 494762 235331
rect 494422 229981 494474 229987
rect 494422 229923 494474 229929
rect 494338 223836 494414 223864
rect 494002 223554 494030 223836
rect 494386 223554 494414 223836
rect 494722 223554 494750 235325
rect 494818 229469 494846 235695
rect 494806 229463 494858 229469
rect 494806 229405 494858 229411
rect 495010 228951 495038 235991
rect 495092 233202 495148 233211
rect 495092 233137 495148 233146
rect 494998 228945 495050 228951
rect 494998 228887 495050 228893
rect 495106 223554 495134 233137
rect 495298 230431 495326 253529
rect 495394 234099 495422 257747
rect 495490 238719 495518 275488
rect 497314 257811 497342 275488
rect 498274 267052 498590 267080
rect 498274 266987 498302 267052
rect 498562 266987 498590 267052
rect 498262 266981 498314 266987
rect 498262 266923 498314 266929
rect 498358 266981 498410 266987
rect 498550 266981 498602 266987
rect 498410 266929 498494 266932
rect 498358 266923 498494 266929
rect 498550 266923 498602 266929
rect 498370 266904 498494 266923
rect 498466 266321 498494 266904
rect 498454 266315 498506 266321
rect 498454 266257 498506 266263
rect 498850 261585 498878 275502
rect 499702 269053 499754 269059
rect 499702 268995 499754 269001
rect 499714 268467 499742 268995
rect 499702 268461 499754 268467
rect 499702 268403 499754 268409
rect 499906 264915 499934 275502
rect 501154 268541 501182 275502
rect 501346 275488 502320 275516
rect 503170 275488 503472 275516
rect 504034 275488 504720 275516
rect 501142 268535 501194 268541
rect 501142 268477 501194 268483
rect 499894 264909 499946 264915
rect 499894 264851 499946 264857
rect 498838 261579 498890 261585
rect 498838 261521 498890 261527
rect 497302 257805 497354 257811
rect 497302 257747 497354 257753
rect 501238 257805 501290 257811
rect 501238 257747 501290 257753
rect 501142 255733 501194 255739
rect 501140 255698 501142 255707
rect 501194 255698 501196 255707
rect 501140 255633 501196 255642
rect 501250 238867 501278 257747
rect 501238 238861 501290 238867
rect 501238 238803 501290 238809
rect 495478 238713 495530 238719
rect 495478 238655 495530 238661
rect 501346 238645 501374 275488
rect 503170 257811 503198 275488
rect 503158 257805 503210 257811
rect 503158 257747 503210 257753
rect 501334 238639 501386 238645
rect 501334 238581 501386 238587
rect 504034 238053 504062 275488
rect 505858 261511 505886 275502
rect 506914 275488 507120 275516
rect 506914 264841 506942 275488
rect 508258 268615 508286 275502
rect 509218 275488 509520 275516
rect 509890 275488 510672 275516
rect 511618 275488 511920 275516
rect 512962 275488 513072 275516
rect 514018 275488 514320 275516
rect 515170 275488 515472 275516
rect 508342 270533 508394 270539
rect 508342 270475 508394 270481
rect 508246 268609 508298 268615
rect 508246 268551 508298 268557
rect 506902 264835 506954 264841
rect 506902 264777 506954 264783
rect 505846 261505 505898 261511
rect 505846 261447 505898 261453
rect 507094 257805 507146 257811
rect 507094 257747 507146 257753
rect 507106 238793 507134 257747
rect 508354 253445 508382 270475
rect 508438 267869 508490 267875
rect 508438 267811 508490 267817
rect 508450 256183 508478 267811
rect 509218 257811 509246 275488
rect 509782 269053 509834 269059
rect 509698 269013 509782 269041
rect 509698 268985 509726 269013
rect 509782 268995 509834 269001
rect 509686 268979 509738 268985
rect 509686 268921 509738 268927
rect 509206 257805 509258 257811
rect 509206 257747 509258 257753
rect 509782 257805 509834 257811
rect 509782 257747 509834 257753
rect 508438 256177 508490 256183
rect 508438 256119 508490 256125
rect 508342 253439 508394 253445
rect 508342 253381 508394 253387
rect 507094 238787 507146 238793
rect 507094 238729 507146 238735
rect 504022 238047 504074 238053
rect 504022 237989 504074 237995
rect 501142 236123 501194 236129
rect 501142 236065 501194 236071
rect 497878 235975 497930 235981
rect 497878 235917 497930 235923
rect 497686 235457 497738 235463
rect 497686 235399 497738 235405
rect 496918 235309 496970 235315
rect 496918 235251 496970 235257
rect 496150 234939 496202 234945
rect 496150 234881 496202 234887
rect 495478 234791 495530 234797
rect 495478 234733 495530 234739
rect 495380 234090 495436 234099
rect 495380 234025 495436 234034
rect 495190 230425 495242 230431
rect 495190 230367 495242 230373
rect 495286 230425 495338 230431
rect 495286 230367 495338 230373
rect 495202 230209 495230 230367
rect 495190 230203 495242 230209
rect 495190 230145 495242 230151
rect 495490 223554 495518 234733
rect 495860 227726 495916 227735
rect 495860 227661 495916 227670
rect 495874 223554 495902 227661
rect 496162 223864 496190 234881
rect 496532 229798 496588 229807
rect 496532 229733 496588 229742
rect 496546 223864 496574 229733
rect 496162 223836 496238 223864
rect 496546 223836 496622 223864
rect 496210 223554 496238 223836
rect 496594 223554 496622 223836
rect 496930 223554 496958 235251
rect 497300 228614 497356 228623
rect 497300 228549 497356 228558
rect 497314 223554 497342 228549
rect 497698 223554 497726 235399
rect 497890 229025 497918 235917
rect 498070 234643 498122 234649
rect 498070 234585 498122 234591
rect 497878 229019 497930 229025
rect 497878 228961 497930 228967
rect 498082 228877 498110 234585
rect 499702 234569 499754 234575
rect 499702 234511 499754 234517
rect 499892 234534 499948 234543
rect 499606 234421 499658 234427
rect 499606 234363 499658 234369
rect 499124 233350 499180 233359
rect 499124 233285 499180 233294
rect 498356 233054 498412 233063
rect 498356 232989 498412 232998
rect 498164 231722 498220 231731
rect 498164 231657 498220 231666
rect 498070 228871 498122 228877
rect 498070 228813 498122 228819
rect 498178 223864 498206 231657
rect 498082 223836 498206 223864
rect 498370 223864 498398 232989
rect 498740 230242 498796 230251
rect 498740 230177 498796 230186
rect 498754 223864 498782 230177
rect 498370 223836 498446 223864
rect 498754 223836 498830 223864
rect 498082 223554 498110 223836
rect 498418 223554 498446 223836
rect 498802 223554 498830 223836
rect 499138 223554 499166 233285
rect 499508 229502 499564 229511
rect 499508 229437 499564 229446
rect 499522 223554 499550 229437
rect 499618 228655 499646 234363
rect 499606 228649 499658 228655
rect 499606 228591 499658 228597
rect 499714 228285 499742 234511
rect 499892 234469 499948 234478
rect 499702 228279 499754 228285
rect 499702 228221 499754 228227
rect 499906 223554 499934 234469
rect 500660 234386 500716 234395
rect 500660 234321 500716 234330
rect 500276 229650 500332 229659
rect 500276 229585 500332 229594
rect 500290 223554 500318 229585
rect 500674 223864 500702 234321
rect 500950 230425 501002 230431
rect 500950 230367 501002 230373
rect 500626 223836 500702 223864
rect 500962 223864 500990 230367
rect 501154 229691 501182 236065
rect 506902 235605 506954 235611
rect 506902 235547 506954 235553
rect 503924 232610 503980 232619
rect 503924 232545 503980 232554
rect 503542 231831 503594 231837
rect 503542 231773 503594 231779
rect 501718 230277 501770 230283
rect 501718 230219 501770 230225
rect 501334 230129 501386 230135
rect 501334 230071 501386 230077
rect 501142 229685 501194 229691
rect 501142 229627 501194 229633
rect 501046 227613 501098 227619
rect 501046 227555 501098 227561
rect 501058 224183 501086 227555
rect 501044 224174 501100 224183
rect 501044 224109 501100 224118
rect 500962 223836 501038 223864
rect 500626 223554 500654 223836
rect 501010 223554 501038 223836
rect 501346 223554 501374 230071
rect 501730 223554 501758 230219
rect 502774 229907 502826 229913
rect 502774 229849 502826 229855
rect 502102 229241 502154 229247
rect 502102 229183 502154 229189
rect 502114 223554 502142 229183
rect 502486 227761 502538 227767
rect 502486 227703 502538 227709
rect 502498 223554 502526 227703
rect 502786 223864 502814 229849
rect 502786 223836 502862 223864
rect 502834 223554 502862 223836
rect 503206 223839 503258 223845
rect 503206 223781 503258 223787
rect 503218 223554 503246 223781
rect 503554 223554 503582 231773
rect 503938 223554 503966 232545
rect 505750 232053 505802 232059
rect 505750 231995 505802 232001
rect 504982 231905 505034 231911
rect 504308 231870 504364 231879
rect 504982 231847 505034 231853
rect 504308 231805 504364 231814
rect 504322 223554 504350 231805
rect 504694 229759 504746 229765
rect 504694 229701 504746 229707
rect 504706 223554 504734 229701
rect 504994 223864 505022 231847
rect 505366 230203 505418 230209
rect 505366 230145 505418 230151
rect 505378 223864 505406 230145
rect 504994 223836 505070 223864
rect 505378 223836 505454 223864
rect 505042 223554 505070 223836
rect 505426 223554 505454 223836
rect 505762 223554 505790 231995
rect 506516 231426 506572 231435
rect 506516 231361 506572 231370
rect 506134 227687 506186 227693
rect 506134 227629 506186 227635
rect 506146 223554 506174 227629
rect 506530 223554 506558 231361
rect 506914 227693 506942 235547
rect 506996 232018 507052 232027
rect 506996 231953 507052 231962
rect 506902 227687 506954 227693
rect 506902 227629 506954 227635
rect 507010 227564 507038 231953
rect 508340 230982 508396 230991
rect 508340 230917 508396 230926
rect 507574 230055 507626 230061
rect 507574 229997 507626 230003
rect 507190 229981 507242 229987
rect 507190 229923 507242 229929
rect 506914 227536 507038 227564
rect 506914 223554 506942 227536
rect 507202 223864 507230 229923
rect 507586 223864 507614 229997
rect 507958 229463 508010 229469
rect 507958 229405 508010 229411
rect 507202 223836 507278 223864
rect 507586 223836 507662 223864
rect 507250 223554 507278 223836
rect 507634 223554 507662 223836
rect 507970 223554 507998 229405
rect 508354 223554 508382 230917
rect 508726 229167 508778 229173
rect 508726 229109 508778 229115
rect 508738 223554 508766 229109
rect 509398 228797 509450 228803
rect 509398 228739 509450 228745
rect 509110 228501 509162 228507
rect 509110 228443 509162 228449
rect 509122 223554 509150 228443
rect 509410 223864 509438 228739
rect 509794 224479 509822 257747
rect 509890 238095 509918 275488
rect 511618 257811 511646 275488
rect 512758 275047 512810 275053
rect 512758 274989 512810 274995
rect 512770 267875 512798 274989
rect 512758 267869 512810 267875
rect 512758 267811 512810 267817
rect 511606 257805 511658 257811
rect 511606 257747 511658 257753
rect 512854 257805 512906 257811
rect 512854 257747 512906 257753
rect 512662 257731 512714 257737
rect 512662 257673 512714 257679
rect 509876 238086 509932 238095
rect 509876 238021 509932 238030
rect 509876 232166 509932 232175
rect 509876 232101 509932 232110
rect 509780 224470 509836 224479
rect 509780 224405 509836 224414
rect 509890 223864 509918 232101
rect 510550 229833 510602 229839
rect 510550 229775 510602 229781
rect 510166 228945 510218 228951
rect 510166 228887 510218 228893
rect 509410 223836 509486 223864
rect 509458 223554 509486 223836
rect 509842 223836 509918 223864
rect 509842 223554 509870 223836
rect 510178 223554 510206 228887
rect 510562 223554 510590 229775
rect 511606 229611 511658 229617
rect 511606 229553 511658 229559
rect 510934 229093 510986 229099
rect 510934 229035 510986 229041
rect 510946 223554 510974 229035
rect 511318 229019 511370 229025
rect 511318 228961 511370 228967
rect 511330 223554 511358 228961
rect 511618 223864 511646 229553
rect 512374 229537 512426 229543
rect 512374 229479 512426 229485
rect 511990 228871 512042 228877
rect 511990 228813 512042 228819
rect 512002 223864 512030 228813
rect 511618 223836 511694 223864
rect 512002 223836 512078 223864
rect 511666 223554 511694 223836
rect 512050 223554 512078 223836
rect 512386 223554 512414 229479
rect 512674 225769 512702 257673
rect 512866 238243 512894 257747
rect 512962 238941 512990 275488
rect 514018 257811 514046 275488
rect 514964 262210 515020 262219
rect 514964 262145 515020 262154
rect 514006 257805 514058 257811
rect 514006 257747 514058 257753
rect 512950 238935 513002 238941
rect 512950 238877 513002 238883
rect 512852 238234 512908 238243
rect 512852 238169 512908 238178
rect 514582 229685 514634 229691
rect 514582 229627 514634 229633
rect 513814 229389 513866 229395
rect 513814 229331 513866 229337
rect 513142 229315 513194 229321
rect 513142 229257 513194 229263
rect 512758 227687 512810 227693
rect 512758 227629 512810 227635
rect 512662 225763 512714 225769
rect 512662 225705 512714 225711
rect 512770 223554 512798 227629
rect 513154 223554 513182 229257
rect 513526 228279 513578 228285
rect 513526 228221 513578 228227
rect 513538 223554 513566 228221
rect 513826 223864 513854 229331
rect 514198 228649 514250 228655
rect 514198 228591 514250 228597
rect 514210 223864 514238 228591
rect 513826 223836 513902 223864
rect 514210 223836 514286 223864
rect 513874 223554 513902 223836
rect 514258 223554 514286 223836
rect 514594 223554 514622 229627
rect 514978 223554 515006 262145
rect 515170 257737 515198 275488
rect 516514 261437 516542 275502
rect 517762 264693 517790 275502
rect 518914 268467 518942 275502
rect 519874 275488 520176 275516
rect 518902 268461 518954 268467
rect 518902 268403 518954 268409
rect 517750 264687 517802 264693
rect 517750 264629 517802 264635
rect 516502 261431 516554 261437
rect 516502 261373 516554 261379
rect 515158 257731 515210 257737
rect 515158 257673 515210 257679
rect 519874 255295 519902 275488
rect 518422 255289 518474 255295
rect 518422 255231 518474 255237
rect 519862 255289 519914 255295
rect 519862 255231 519914 255237
rect 518434 239015 518462 255231
rect 518422 239009 518474 239015
rect 518422 238951 518474 238957
rect 521314 224627 521342 275502
rect 522562 274609 522590 275502
rect 522262 274603 522314 274609
rect 522262 274545 522314 274551
rect 522550 274603 522602 274609
rect 522550 274545 522602 274551
rect 521974 270607 522026 270613
rect 521974 270549 522026 270555
rect 521398 267943 521450 267949
rect 521398 267885 521450 267891
rect 521410 225621 521438 267885
rect 521986 260623 522014 270549
rect 522274 267949 522302 274545
rect 522262 267943 522314 267949
rect 522262 267885 522314 267891
rect 523714 261289 523742 275502
rect 524962 264767 524990 275502
rect 526114 269207 526142 275502
rect 527266 275488 527376 275516
rect 528226 275488 528528 275516
rect 529474 275488 529776 275516
rect 526102 269201 526154 269207
rect 526102 269143 526154 269149
rect 524950 264761 525002 264767
rect 524950 264703 525002 264709
rect 523702 261283 523754 261289
rect 523702 261225 523754 261231
rect 521974 260617 522026 260623
rect 521974 260559 522026 260565
rect 527062 257805 527114 257811
rect 527062 257747 527114 257753
rect 527074 226583 527102 257747
rect 527158 257731 527210 257737
rect 527158 257673 527210 257679
rect 527170 227397 527198 257673
rect 527266 238201 527294 275488
rect 528226 257811 528254 275488
rect 528214 257805 528266 257811
rect 528214 257747 528266 257753
rect 529474 257737 529502 275488
rect 529844 273458 529900 273467
rect 529900 273416 530078 273444
rect 529844 273393 529900 273402
rect 530050 273319 530078 273416
rect 530036 273310 530092 273319
rect 530036 273245 530092 273254
rect 530914 261215 530942 275502
rect 532066 264619 532094 275502
rect 533218 268911 533246 275502
rect 533410 275488 534384 275516
rect 535330 275488 535632 275516
rect 535714 275488 536784 275516
rect 533206 268905 533258 268911
rect 533206 268847 533258 268853
rect 532054 264613 532106 264619
rect 532054 264555 532106 264561
rect 530902 261209 530954 261215
rect 530902 261151 530954 261157
rect 533014 257805 533066 257811
rect 533014 257747 533066 257753
rect 529462 257731 529514 257737
rect 529462 257673 529514 257679
rect 532918 247741 532970 247747
rect 532918 247683 532970 247689
rect 532930 238349 532958 247683
rect 532918 238343 532970 238349
rect 532918 238285 532970 238291
rect 527254 238195 527306 238201
rect 527254 238137 527306 238143
rect 533026 237905 533054 257747
rect 533410 247747 533438 275488
rect 535330 257811 535358 275488
rect 535714 267283 535742 275488
rect 535702 267277 535754 267283
rect 535702 267219 535754 267225
rect 536182 267277 536234 267283
rect 536182 267219 536234 267225
rect 535510 266833 535562 266839
rect 535606 266833 535658 266839
rect 535562 266781 535606 266784
rect 535510 266775 535658 266781
rect 535522 266756 535646 266775
rect 535510 266685 535562 266691
rect 535426 266645 535510 266673
rect 535426 266321 535454 266645
rect 535510 266627 535562 266633
rect 535798 266611 535850 266617
rect 535990 266611 536042 266617
rect 535850 266571 535990 266599
rect 535798 266553 535850 266559
rect 535990 266553 536042 266559
rect 535702 266537 535754 266543
rect 535702 266479 535754 266485
rect 535414 266315 535466 266321
rect 535414 266257 535466 266263
rect 535714 266247 535742 266479
rect 535702 266241 535754 266247
rect 535702 266183 535754 266189
rect 536194 263583 536222 267219
rect 535702 263577 535754 263583
rect 535702 263519 535754 263525
rect 536182 263577 536234 263583
rect 536182 263519 536234 263525
rect 535318 257805 535370 257811
rect 535318 257747 535370 257753
rect 533398 247741 533450 247747
rect 533398 247683 533450 247689
rect 533014 237899 533066 237905
rect 533014 237841 533066 237847
rect 535714 234247 535742 263519
rect 538018 261141 538046 275502
rect 538484 267242 538540 267251
rect 538484 267177 538540 267186
rect 538498 266691 538526 267177
rect 538486 266685 538538 266691
rect 538486 266627 538538 266633
rect 539170 264545 539198 275502
rect 540418 270687 540446 275502
rect 541584 275488 542078 275516
rect 540406 270681 540458 270687
rect 540406 270623 540458 270629
rect 541750 266315 541802 266321
rect 541750 266257 541802 266263
rect 541462 266167 541514 266173
rect 541462 266109 541514 266115
rect 539158 264539 539210 264545
rect 539158 264481 539210 264487
rect 538006 261135 538058 261141
rect 538006 261077 538058 261083
rect 541474 255813 541502 266109
rect 541654 257805 541706 257811
rect 541654 257747 541706 257753
rect 541462 255807 541514 255813
rect 541462 255749 541514 255755
rect 538484 255661 538540 255670
rect 538484 255596 538540 255605
rect 541462 249147 541514 249153
rect 541462 249089 541514 249095
rect 541474 238423 541502 249089
rect 541558 247741 541610 247747
rect 541558 247683 541610 247689
rect 541462 238417 541514 238423
rect 541462 238359 541514 238365
rect 541570 237831 541598 247683
rect 541666 239681 541694 257747
rect 541762 247747 541790 266257
rect 542050 266173 542078 275488
rect 542818 266321 542846 275502
rect 543682 275488 543984 275516
rect 542806 266315 542858 266321
rect 542806 266257 542858 266263
rect 542038 266167 542090 266173
rect 542038 266109 542090 266115
rect 543682 257811 543710 275488
rect 545218 260147 545246 275502
rect 545686 266537 545738 266543
rect 545686 266479 545738 266485
rect 545698 266247 545726 266479
rect 545686 266241 545738 266247
rect 545686 266183 545738 266189
rect 546370 264397 546398 275502
rect 547522 267431 547550 275502
rect 548770 268763 548798 275502
rect 548758 268757 548810 268763
rect 548758 268699 548810 268705
rect 547510 267425 547562 267431
rect 547510 267367 547562 267373
rect 546358 264391 546410 264397
rect 546358 264333 546410 264339
rect 549826 261067 549854 275502
rect 551074 270613 551102 275502
rect 551062 270607 551114 270613
rect 551062 270549 551114 270555
rect 552226 269133 552254 275502
rect 552214 269127 552266 269133
rect 552214 269069 552266 269075
rect 549814 261061 549866 261067
rect 549814 261003 549866 261009
rect 553474 260993 553502 275502
rect 554626 261733 554654 275502
rect 555874 266807 555902 275502
rect 555860 266798 555916 266807
rect 555860 266733 555916 266742
rect 554614 261727 554666 261733
rect 554614 261669 554666 261675
rect 553462 260987 553514 260993
rect 553462 260929 553514 260935
rect 557026 260295 557054 275502
rect 558274 264471 558302 275502
rect 559426 267103 559454 275502
rect 559412 267094 559468 267103
rect 559412 267029 559468 267038
rect 558262 264465 558314 264471
rect 558262 264407 558314 264413
rect 560674 260443 560702 275502
rect 561524 267242 561580 267251
rect 561524 267177 561580 267186
rect 561538 266691 561566 267177
rect 561526 266685 561578 266691
rect 561526 266627 561578 266633
rect 561826 261659 561854 275502
rect 562978 266955 563006 275502
rect 564226 270465 564254 275502
rect 564214 270459 564266 270465
rect 564214 270401 564266 270407
rect 562964 266946 563020 266955
rect 562964 266881 563020 266890
rect 565378 264249 565406 275502
rect 566530 270539 566558 275502
rect 566518 270533 566570 270539
rect 566518 270475 566570 270481
rect 567682 270391 567710 275502
rect 567670 270385 567722 270391
rect 567670 270327 567722 270333
rect 568930 264323 568958 275502
rect 570082 266659 570110 275502
rect 570262 266907 570314 266913
rect 570262 266849 570314 266855
rect 570274 266691 570302 266849
rect 570262 266685 570314 266691
rect 570068 266650 570124 266659
rect 570262 266627 570314 266633
rect 570068 266585 570124 266594
rect 568918 264317 568970 264323
rect 568918 264259 568970 264265
rect 565366 264243 565418 264249
rect 565366 264185 565418 264191
rect 561814 261653 561866 261659
rect 561814 261595 561866 261601
rect 571330 260697 571358 275502
rect 572482 264175 572510 275502
rect 573730 266511 573758 275502
rect 573716 266502 573772 266511
rect 573716 266437 573772 266446
rect 572470 264169 572522 264175
rect 572470 264111 572522 264117
rect 574882 260845 574910 275502
rect 576130 264101 576158 275502
rect 577282 270317 577310 275502
rect 577270 270311 577322 270317
rect 577270 270253 577322 270259
rect 578434 270169 578462 275502
rect 578422 270163 578474 270169
rect 578422 270105 578474 270111
rect 576118 264095 576170 264101
rect 576118 264037 576170 264043
rect 579682 264027 579710 275502
rect 580834 270243 580862 275502
rect 580822 270237 580874 270243
rect 580822 270179 580874 270185
rect 582082 270095 582110 275502
rect 582070 270089 582122 270095
rect 582070 270031 582122 270037
rect 579670 264021 579722 264027
rect 579670 263963 579722 263969
rect 583138 263879 583166 275502
rect 583126 263873 583178 263879
rect 583126 263815 583178 263821
rect 584386 262071 584414 275502
rect 585538 270021 585566 275502
rect 585526 270015 585578 270021
rect 585526 269957 585578 269963
rect 586786 263953 586814 275502
rect 587938 266363 587966 275502
rect 589186 269947 589214 275502
rect 589174 269941 589226 269947
rect 589174 269883 589226 269889
rect 590230 266833 590282 266839
rect 590228 266798 590230 266807
rect 590282 266798 590284 266807
rect 590134 266759 590186 266765
rect 590228 266733 590284 266742
rect 590134 266701 590186 266707
rect 590146 266659 590174 266701
rect 590132 266650 590188 266659
rect 590132 266585 590188 266594
rect 587924 266354 587980 266363
rect 587924 266289 587980 266298
rect 586774 263947 586826 263953
rect 586774 263889 586826 263895
rect 584372 262062 584428 262071
rect 584372 261997 584428 262006
rect 574870 260839 574922 260845
rect 574870 260781 574922 260787
rect 571318 260691 571370 260697
rect 571318 260633 571370 260639
rect 560660 260434 560716 260443
rect 560660 260369 560716 260378
rect 557012 260286 557068 260295
rect 557012 260221 557068 260230
rect 545204 260138 545260 260147
rect 545204 260073 545260 260082
rect 590338 259513 590366 275502
rect 590518 266833 590570 266839
rect 590516 266798 590518 266807
rect 590570 266798 590572 266807
rect 590516 266733 590572 266742
rect 590614 266759 590666 266765
rect 590614 266701 590666 266707
rect 590626 266659 590654 266701
rect 590612 266650 590668 266659
rect 590612 266585 590668 266594
rect 591586 261923 591614 275502
rect 592738 263805 592766 275502
rect 593890 265433 593918 275502
rect 593878 265427 593930 265433
rect 593878 265369 593930 265375
rect 592726 263799 592778 263805
rect 592726 263741 592778 263747
rect 591572 261914 591628 261923
rect 591572 261849 591628 261858
rect 595138 261775 595166 275502
rect 596290 269799 596318 275502
rect 596278 269793 596330 269799
rect 596278 269735 596330 269741
rect 597538 266025 597566 275502
rect 598690 269873 598718 275502
rect 598678 269867 598730 269873
rect 598678 269809 598730 269815
rect 599842 269725 599870 275502
rect 599830 269719 599882 269725
rect 599830 269661 599882 269667
rect 600994 267209 601022 275502
rect 600982 267203 601034 267209
rect 600982 267145 601034 267151
rect 597526 266019 597578 266025
rect 597526 265961 597578 265967
rect 595124 261766 595180 261775
rect 595124 261701 595180 261710
rect 602242 261627 602270 275502
rect 603394 269651 603422 275502
rect 603382 269645 603434 269651
rect 603382 269587 603434 269593
rect 604642 267135 604670 275502
rect 605794 269429 605822 275502
rect 605782 269423 605834 269429
rect 605782 269365 605834 269371
rect 604630 267129 604682 267135
rect 604630 267071 604682 267077
rect 607042 264587 607070 275502
rect 608194 267061 608222 275502
rect 608182 267055 608234 267061
rect 608182 266997 608234 267003
rect 607028 264578 607084 264587
rect 607028 264513 607084 264522
rect 602228 261618 602284 261627
rect 602228 261553 602284 261562
rect 609346 261479 609374 275502
rect 610486 267129 610538 267135
rect 610486 267071 610538 267077
rect 610294 267055 610346 267061
rect 610294 266997 610346 267003
rect 610306 266765 610334 266997
rect 610498 266913 610526 267071
rect 610486 266907 610538 266913
rect 610486 266849 610538 266855
rect 610390 266833 610442 266839
rect 610388 266798 610390 266807
rect 610442 266798 610444 266807
rect 610294 266759 610346 266765
rect 610388 266733 610444 266742
rect 610294 266701 610346 266707
rect 610594 264439 610622 275502
rect 611746 266987 611774 275502
rect 612022 267055 612074 267061
rect 612022 266997 612074 267003
rect 611734 266981 611786 266987
rect 611734 266923 611786 266929
rect 610678 266833 610730 266839
rect 610676 266798 610678 266807
rect 610730 266798 610732 266807
rect 612034 266765 612062 266997
rect 610676 266733 610732 266742
rect 612022 266759 612074 266765
rect 612022 266701 612074 266707
rect 610580 264430 610636 264439
rect 610580 264365 610636 264374
rect 609332 261470 609388 261479
rect 609332 261405 609388 261414
rect 612994 261331 613022 275502
rect 614146 264291 614174 275502
rect 614132 264282 614188 264291
rect 614132 264217 614188 264226
rect 612980 261322 613036 261331
rect 612980 261257 613036 261266
rect 615394 260919 615422 275502
rect 616450 269355 616478 275502
rect 616438 269349 616490 269355
rect 616438 269291 616490 269297
rect 617698 264143 617726 275502
rect 617684 264134 617740 264143
rect 617684 264069 617740 264078
rect 615382 260913 615434 260919
rect 615382 260855 615434 260861
rect 618850 260771 618878 275502
rect 620098 269503 620126 275502
rect 621250 269577 621278 275502
rect 621238 269571 621290 269577
rect 621238 269513 621290 269519
rect 620086 269497 620138 269503
rect 620086 269439 620138 269445
rect 622102 267795 622154 267801
rect 622102 267737 622154 267743
rect 621910 267129 621962 267135
rect 621910 267071 621962 267077
rect 621922 266895 621950 267071
rect 622114 266895 622142 267737
rect 621922 266867 622142 266895
rect 622498 266099 622526 275502
rect 622486 266093 622538 266099
rect 622486 266035 622538 266041
rect 623650 261183 623678 275502
rect 624802 263731 624830 275502
rect 626050 266839 626078 275502
rect 626038 266833 626090 266839
rect 626038 266775 626090 266781
rect 624790 263725 624842 263731
rect 624790 263667 624842 263673
rect 623636 261174 623692 261183
rect 623636 261109 623692 261118
rect 627202 261035 627230 275502
rect 628450 263657 628478 275502
rect 629602 266765 629630 275502
rect 629590 266759 629642 266765
rect 629590 266701 629642 266707
rect 628438 263651 628490 263657
rect 628438 263593 628490 263599
rect 627188 261026 627244 261035
rect 627188 260961 627244 260970
rect 618838 260765 618890 260771
rect 618838 260707 618890 260713
rect 590326 259507 590378 259513
rect 590326 259449 590378 259455
rect 630658 259236 630686 275636
rect 632002 263995 632030 275502
rect 633154 267801 633182 275502
rect 633142 267795 633194 267801
rect 633142 267737 633194 267743
rect 631988 263986 632044 263995
rect 631988 263921 632044 263930
rect 634306 260887 634334 275502
rect 635554 263847 635582 275502
rect 636706 266617 636734 275502
rect 637666 275488 637968 275516
rect 636694 266611 636746 266617
rect 636694 266553 636746 266559
rect 635540 263838 635596 263847
rect 635540 263773 635596 263782
rect 634292 260878 634348 260887
rect 634292 260813 634348 260822
rect 630658 259208 630782 259236
rect 543670 257805 543722 257811
rect 543670 257747 543722 257753
rect 630754 256257 630782 259208
rect 637666 256331 637694 275488
rect 639106 263699 639134 275502
rect 640258 266543 640286 275502
rect 640246 266537 640298 266543
rect 640246 266479 640298 266485
rect 639092 263690 639148 263699
rect 639092 263625 639148 263634
rect 641506 260739 641534 275502
rect 642658 263551 642686 275502
rect 643906 266469 643934 275502
rect 643894 266463 643946 266469
rect 643894 266405 643946 266411
rect 642644 263542 642700 263551
rect 642644 263477 642700 263486
rect 641492 260730 641548 260739
rect 641492 260665 641548 260674
rect 645058 260591 645086 275502
rect 645142 273419 645194 273425
rect 645142 273361 645194 273367
rect 645154 273171 645182 273361
rect 645140 273162 645196 273171
rect 645140 273097 645196 273106
rect 646306 262177 646334 275502
rect 647458 266395 647486 275502
rect 648706 269281 648734 275502
rect 649378 275053 649406 980505
rect 649474 953337 649502 980727
rect 649462 953331 649514 953337
rect 649462 953273 649514 953279
rect 649462 927431 649514 927437
rect 649462 927373 649514 927379
rect 649366 275047 649418 275053
rect 649366 274989 649418 274995
rect 648694 269275 648746 269281
rect 648694 269217 648746 269223
rect 647446 266389 647498 266395
rect 647446 266331 647498 266337
rect 646294 262171 646346 262177
rect 646294 262113 646346 262119
rect 645044 260582 645100 260591
rect 645044 260517 645100 260526
rect 640726 256399 640778 256405
rect 640726 256341 640778 256347
rect 637654 256325 637706 256331
rect 637654 256267 637706 256273
rect 630742 256251 630794 256257
rect 630742 256193 630794 256199
rect 622004 255846 622060 255855
rect 541846 255807 541898 255813
rect 622004 255781 622060 255790
rect 541846 255749 541898 255755
rect 541858 249153 541886 255749
rect 622018 255739 622046 255781
rect 570166 255733 570218 255739
rect 590518 255733 590570 255739
rect 570218 255681 570398 255684
rect 570166 255675 570398 255681
rect 570178 255665 570398 255675
rect 590338 255681 590518 255684
rect 601942 255733 601994 255739
rect 590338 255675 590570 255681
rect 601940 255698 601942 255707
rect 622006 255733 622058 255739
rect 601994 255698 601996 255707
rect 590338 255665 590558 255675
rect 570178 255659 570410 255665
rect 570178 255656 570358 255659
rect 570358 255601 570410 255607
rect 590326 255659 590558 255665
rect 590378 255656 590558 255659
rect 622006 255675 622058 255681
rect 630646 255733 630698 255739
rect 630698 255681 630878 255684
rect 630646 255675 630878 255681
rect 630658 255665 630878 255675
rect 630658 255659 630890 255665
rect 630658 255656 630838 255659
rect 601940 255633 601996 255642
rect 590326 255601 590378 255607
rect 630838 255601 630890 255607
rect 541846 249147 541898 249153
rect 541846 249089 541898 249095
rect 541750 247741 541802 247747
rect 541750 247683 541802 247689
rect 541654 239675 541706 239681
rect 541654 239617 541706 239623
rect 541558 237825 541610 237831
rect 541558 237767 541610 237773
rect 535700 234238 535756 234247
rect 535700 234173 535756 234182
rect 633814 229611 633866 229617
rect 633814 229553 633866 229559
rect 633142 229537 633194 229543
rect 633142 229479 633194 229485
rect 632758 229463 632810 229469
rect 632758 229405 632810 229411
rect 632374 229389 632426 229395
rect 632374 229331 632426 229337
rect 631990 229315 632042 229321
rect 631990 229257 632042 229263
rect 631606 229241 631658 229247
rect 631606 229183 631658 229189
rect 631318 229167 631370 229173
rect 631318 229109 631370 229115
rect 541366 229019 541418 229025
rect 541366 228961 541418 228967
rect 541378 227619 541406 228961
rect 539638 227613 539690 227619
rect 539638 227555 539690 227561
rect 541366 227613 541418 227619
rect 541366 227555 541418 227561
rect 527158 227391 527210 227397
rect 527158 227333 527210 227339
rect 527062 226577 527114 226583
rect 527062 226519 527114 226525
rect 521398 225615 521450 225621
rect 521398 225557 521450 225563
rect 521300 224618 521356 224627
rect 521300 224553 521356 224562
rect 539650 223554 539678 227555
rect 631330 224035 631358 229109
rect 631316 224026 631372 224035
rect 631316 223961 631372 223970
rect 631330 223864 631358 223961
rect 631618 223887 631646 229183
rect 632002 224183 632030 229257
rect 631988 224174 632044 224183
rect 631988 224109 632044 224118
rect 631282 223836 631358 223864
rect 631604 223878 631660 223887
rect 631282 223554 631310 223836
rect 631604 223813 631660 223822
rect 631618 223554 631646 223813
rect 632002 223554 632030 224109
rect 632386 223887 632414 229331
rect 632770 223887 632798 229405
rect 633154 223887 633182 229479
rect 633526 229093 633578 229099
rect 633526 229035 633578 229041
rect 633538 224035 633566 229035
rect 633524 224026 633580 224035
rect 633524 223961 633580 223970
rect 632372 223878 632428 223887
rect 632372 223813 632428 223822
rect 632756 223878 632812 223887
rect 632756 223813 632812 223822
rect 633140 223878 633196 223887
rect 633538 223864 633566 223961
rect 633140 223813 633196 223822
rect 633490 223836 633566 223864
rect 632386 223554 632414 223813
rect 632770 223554 632798 223813
rect 633154 223716 633182 223813
rect 633106 223688 633182 223716
rect 633106 223554 633134 223688
rect 633490 223554 633518 223836
rect 204982 223099 205034 223105
rect 204982 223041 205034 223047
rect 633826 222976 633854 229553
rect 204898 222948 205152 222976
rect 633826 222962 634142 222976
rect 633840 222948 634142 222962
rect 204886 222877 204938 222883
rect 204886 222819 204938 222825
rect 204898 207417 204926 222819
rect 204994 222703 205022 222948
rect 204980 222694 205036 222703
rect 204980 222629 205036 222638
rect 204886 207411 204938 207417
rect 204886 207353 204938 207359
rect 204982 132523 205034 132529
rect 204982 132465 205034 132471
rect 204886 112395 204938 112401
rect 204886 112337 204938 112343
rect 204898 96436 204926 112337
rect 204994 96565 205022 132465
rect 204982 96559 205034 96565
rect 204982 96501 205034 96507
rect 204898 96408 205022 96436
rect 204886 96337 204938 96343
rect 204886 96279 204938 96285
rect 204898 86691 204926 96279
rect 204884 86682 204940 86691
rect 204884 86617 204940 86626
rect 204886 86569 204938 86575
rect 204886 86511 204938 86517
rect 204790 58967 204842 58973
rect 204790 58909 204842 58915
rect 204692 58858 204748 58867
rect 204692 58793 204748 58802
rect 204610 58668 204734 58696
rect 204596 58414 204652 58423
rect 204596 58349 204652 58358
rect 204502 57339 204554 57345
rect 204502 57281 204554 57287
rect 204500 57230 204556 57239
rect 204500 57165 204556 57174
rect 204514 53423 204542 57165
rect 204502 53417 204554 53423
rect 204502 53359 204554 53365
rect 204610 53275 204638 58349
rect 204706 56309 204734 58668
rect 204694 56303 204746 56309
rect 204694 56245 204746 56251
rect 204692 56194 204748 56203
rect 204692 56129 204748 56138
rect 204502 53269 204554 53275
rect 204502 53211 204554 53217
rect 204598 53269 204650 53275
rect 204598 53211 204650 53217
rect 204406 53121 204458 53127
rect 204308 53086 204364 53095
rect 204406 53063 204458 53069
rect 204514 53072 204542 53211
rect 204514 53044 204638 53072
rect 204308 53021 204364 53030
rect 204226 52896 204542 52924
rect 204514 51721 204542 52896
rect 204502 51715 204554 51721
rect 204502 51657 204554 51663
rect 204610 51647 204638 53044
rect 204706 52091 204734 56129
rect 204788 55158 204844 55167
rect 204788 55093 204844 55102
rect 204694 52085 204746 52091
rect 204694 52027 204746 52033
rect 204802 51943 204830 55093
rect 204898 54575 204926 86511
rect 204994 59121 205022 96408
rect 634006 92341 634058 92347
rect 634006 92283 634058 92289
rect 204982 59115 205034 59121
rect 204982 59057 205034 59063
rect 204982 58967 205034 58973
rect 204982 58909 205034 58915
rect 204994 54829 205022 58909
rect 204982 54823 205034 54829
rect 204982 54765 205034 54771
rect 204980 54714 205036 54723
rect 204980 54649 205036 54658
rect 204884 54566 204940 54575
rect 204884 54501 204940 54510
rect 204994 53941 205022 54649
rect 634018 54404 634046 92283
rect 633840 54376 634046 54404
rect 210356 54270 210412 54279
rect 205942 54231 205994 54237
rect 214772 54270 214828 54279
rect 210412 54228 210480 54256
rect 214704 54228 214772 54256
rect 210356 54205 210412 54214
rect 214964 54270 215020 54279
rect 214896 54228 214964 54256
rect 214772 54205 214828 54214
rect 627092 54270 627148 54279
rect 215170 54237 215280 54256
rect 214964 54205 215020 54214
rect 215158 54231 215280 54237
rect 205942 54173 205994 54179
rect 215210 54228 215280 54231
rect 626880 54228 627092 54256
rect 629588 54270 629644 54279
rect 629424 54228 629588 54256
rect 627092 54205 627148 54214
rect 632016 54237 632318 54256
rect 632016 54231 632330 54237
rect 632016 54228 632278 54231
rect 629588 54205 629644 54214
rect 215158 54173 215210 54179
rect 632278 54173 632330 54179
rect 204982 53935 205034 53941
rect 204982 53877 205034 53883
rect 204898 53784 205152 53812
rect 204790 51937 204842 51943
rect 204692 51902 204748 51911
rect 204790 51879 204842 51885
rect 204692 51837 204748 51846
rect 204598 51641 204650 51647
rect 204034 51564 204542 51592
rect 204598 51583 204650 51589
rect 204514 48613 204542 51564
rect 204706 48687 204734 51837
rect 204694 48681 204746 48687
rect 204694 48623 204746 48629
rect 204502 48607 204554 48613
rect 204502 48549 204554 48555
rect 203830 48533 203882 48539
rect 203830 48475 203882 48481
rect 203734 48459 203786 48465
rect 203734 48401 203786 48407
rect 203446 48237 203498 48243
rect 203446 48179 203498 48185
rect 203350 47941 203402 47947
rect 203350 47883 203402 47889
rect 203254 47867 203306 47873
rect 203254 47809 203306 47815
rect 202486 46609 202538 46615
rect 202486 46551 202538 46557
rect 202294 46461 202346 46467
rect 202294 46403 202346 46409
rect 202198 46165 202250 46171
rect 202198 46107 202250 46113
rect 201334 42169 201386 42175
rect 201334 42111 201386 42117
rect 187604 41838 187660 41847
rect 187344 41796 187604 41824
rect 194324 41838 194380 41847
rect 194064 41796 194324 41824
rect 187604 41773 187660 41782
rect 194324 41773 194380 41782
rect 204898 40811 204926 53784
rect 205330 53516 205358 53798
rect 205330 53488 205406 53516
rect 205270 53121 205322 53127
rect 205270 53063 205322 53069
rect 205174 52085 205226 52091
rect 205174 52027 205226 52033
rect 205078 51937 205130 51943
rect 205078 51879 205130 51885
rect 205090 45399 205118 51879
rect 205076 45390 205132 45399
rect 205076 45325 205132 45334
rect 205186 45209 205214 52027
rect 205174 45203 205226 45209
rect 205174 45145 205226 45151
rect 205282 44839 205310 53063
rect 205378 52091 205406 53488
rect 205366 52085 205418 52091
rect 205366 52027 205418 52033
rect 205474 45103 205502 53798
rect 205558 53269 205610 53275
rect 205558 53211 205610 53217
rect 205460 45094 205516 45103
rect 205460 45029 205516 45038
rect 205270 44833 205322 44839
rect 205270 44775 205322 44781
rect 205570 44691 205598 53211
rect 205666 52207 205694 53798
rect 205762 53784 205872 53812
rect 205652 52198 205708 52207
rect 205652 52133 205708 52142
rect 205762 44955 205790 53784
rect 205846 53121 205898 53127
rect 205844 53086 205846 53095
rect 205898 53086 205900 53095
rect 205844 53021 205900 53030
rect 205954 51869 205982 54173
rect 206326 54157 206378 54163
rect 214966 54157 215018 54163
rect 208532 54122 208588 54131
rect 206378 54105 206448 54108
rect 206326 54099 206448 54105
rect 206338 54080 206448 54099
rect 212564 54122 212620 54131
rect 208588 54080 208656 54108
rect 208532 54057 208588 54066
rect 633718 54157 633770 54163
rect 632948 54122 633004 54131
rect 214966 54099 215018 54105
rect 212564 54057 212620 54066
rect 214774 54083 214826 54089
rect 208148 53974 208204 53983
rect 206134 53935 206186 53941
rect 208204 53932 208272 53960
rect 208148 53909 208204 53918
rect 206134 53877 206186 53883
rect 206050 51943 206078 53798
rect 206038 51937 206090 51943
rect 206038 51879 206090 51885
rect 205942 51863 205994 51869
rect 205942 51805 205994 51811
rect 206146 45251 206174 53877
rect 206326 53861 206378 53867
rect 210740 53826 210796 53835
rect 206326 53803 206378 53809
rect 206242 45547 206270 53798
rect 206338 53664 206366 53803
rect 206338 53636 206558 53664
rect 206530 53423 206558 53636
rect 206326 53417 206378 53423
rect 206326 53359 206378 53365
rect 206518 53417 206570 53423
rect 206518 53359 206570 53365
rect 206228 45538 206284 45547
rect 206228 45473 206284 45482
rect 206132 45242 206188 45251
rect 206132 45177 206188 45186
rect 205748 44946 205804 44955
rect 205748 44881 205804 44890
rect 206338 44807 206366 53359
rect 206324 44798 206380 44807
rect 206324 44733 206380 44742
rect 205558 44685 205610 44691
rect 205558 44627 205610 44633
rect 206626 42397 206654 53798
rect 206708 53530 206764 53539
rect 206708 53465 206764 53474
rect 206722 53095 206750 53465
rect 206708 53086 206764 53095
rect 206708 53021 206764 53030
rect 206818 52059 206846 53798
rect 206976 53784 207038 53812
rect 206900 53382 206956 53391
rect 206900 53317 206956 53326
rect 206914 53275 206942 53317
rect 206902 53269 206954 53275
rect 206902 53211 206954 53217
rect 206804 52050 206860 52059
rect 206804 51985 206860 51994
rect 207010 45135 207038 53784
rect 207154 53664 207182 53798
rect 207106 53650 207182 53664
rect 207092 53641 207182 53650
rect 207148 53636 207182 53641
rect 207092 53576 207148 53585
rect 207346 53516 207374 53798
rect 207490 53784 207552 53812
rect 207490 53645 207518 53784
rect 207478 53639 207530 53645
rect 207478 53581 207530 53587
rect 207574 53639 207626 53645
rect 207574 53581 207626 53587
rect 207586 53539 207614 53581
rect 207572 53530 207628 53539
rect 207346 53488 207422 53516
rect 206998 45129 207050 45135
rect 206998 45071 207050 45077
rect 207394 45061 207422 53488
rect 207572 53465 207628 53474
rect 207382 45055 207434 45061
rect 207382 44997 207434 45003
rect 206614 42391 206666 42397
rect 206614 42333 206666 42339
rect 207682 42101 207710 53798
rect 207874 52355 207902 53798
rect 207860 52346 207916 52355
rect 207860 52281 207916 52290
rect 207956 46574 208012 46583
rect 207956 46509 208012 46518
rect 207860 46426 207916 46435
rect 207860 46361 207862 46370
rect 207914 46361 207916 46370
rect 207862 46329 207914 46335
rect 207970 46319 207998 46509
rect 207958 46313 208010 46319
rect 207958 46255 208010 46261
rect 208066 44987 208094 53798
rect 208342 47497 208394 47503
rect 208342 47439 208394 47445
rect 208354 46541 208382 47439
rect 208342 46535 208394 46541
rect 208342 46477 208394 46483
rect 208054 44981 208106 44987
rect 208054 44923 208106 44929
rect 207670 42095 207722 42101
rect 207670 42037 207722 42043
rect 208450 41731 208478 53798
rect 208726 47867 208778 47873
rect 208726 47809 208778 47815
rect 208738 47577 208766 47809
rect 208726 47571 208778 47577
rect 208726 47513 208778 47519
rect 208534 46609 208586 46615
rect 208532 46574 208534 46583
rect 208586 46574 208588 46583
rect 208532 46509 208588 46518
rect 208834 44659 208862 53798
rect 209026 53539 209054 53798
rect 209184 53784 209246 53812
rect 209012 53530 209068 53539
rect 209012 53465 209068 53474
rect 208918 48681 208970 48687
rect 208918 48623 208970 48629
rect 208930 47947 208958 48623
rect 208918 47941 208970 47947
rect 208918 47883 208970 47889
rect 209218 44913 209246 53784
rect 209362 53664 209390 53798
rect 209314 53636 209390 53664
rect 209314 53391 209342 53636
rect 209554 53516 209582 53798
rect 209746 53645 209774 53798
rect 209734 53639 209786 53645
rect 209734 53581 209786 53587
rect 209554 53488 209630 53516
rect 209300 53382 209356 53391
rect 209300 53317 209356 53326
rect 209302 48459 209354 48465
rect 209302 48401 209354 48407
rect 209314 47429 209342 48401
rect 209302 47423 209354 47429
rect 209302 47365 209354 47371
rect 209398 47423 209450 47429
rect 209398 47365 209450 47371
rect 209410 46837 209438 47365
rect 209398 46831 209450 46837
rect 209398 46773 209450 46779
rect 209206 44907 209258 44913
rect 209206 44849 209258 44855
rect 209602 44765 209630 53488
rect 209890 52683 209918 53798
rect 210082 53571 210110 53798
rect 210070 53565 210122 53571
rect 210070 53507 210122 53513
rect 210274 53349 210302 53798
rect 210262 53343 210314 53349
rect 210262 53285 210314 53291
rect 210658 53201 210686 53798
rect 210740 53761 210796 53770
rect 210754 53645 210782 53761
rect 210742 53639 210794 53645
rect 210742 53581 210794 53587
rect 210646 53195 210698 53201
rect 210646 53137 210698 53143
rect 209878 52677 209930 52683
rect 209878 52619 209930 52625
rect 210850 51869 210878 53798
rect 211042 53053 211070 53798
rect 211234 53423 211262 53798
rect 211392 53784 211454 53812
rect 211222 53417 211274 53423
rect 211222 53359 211274 53365
rect 211030 53047 211082 53053
rect 211030 52989 211082 52995
rect 211426 52609 211454 53784
rect 211570 53645 211598 53798
rect 211558 53639 211610 53645
rect 211558 53581 211610 53587
rect 211762 53516 211790 53798
rect 211954 53645 211982 53798
rect 211942 53639 211994 53645
rect 211942 53581 211994 53587
rect 211714 53488 211790 53516
rect 211714 52905 211742 53488
rect 211702 52899 211754 52905
rect 211702 52841 211754 52847
rect 212098 52757 212126 53798
rect 212086 52751 212138 52757
rect 212086 52693 212138 52699
rect 211414 52603 211466 52609
rect 211414 52545 211466 52551
rect 210838 51863 210890 51869
rect 210838 51805 210890 51811
rect 212290 51721 212318 53798
rect 212482 52017 212510 53798
rect 212578 53539 212606 54057
rect 214774 54025 214826 54031
rect 212564 53530 212620 53539
rect 212564 53465 212620 53474
rect 212674 52017 212702 53798
rect 212866 53497 212894 53798
rect 212854 53491 212906 53497
rect 212854 53433 212906 53439
rect 212470 52011 212522 52017
rect 212470 51953 212522 51959
rect 212662 52011 212714 52017
rect 212662 51953 212714 51959
rect 212278 51715 212330 51721
rect 212278 51657 212330 51663
rect 213058 51647 213086 53798
rect 213250 52979 213278 53798
rect 213442 53645 213470 53798
rect 213600 53784 213662 53812
rect 213430 53639 213482 53645
rect 213430 53581 213482 53587
rect 213238 52973 213290 52979
rect 213238 52915 213290 52921
rect 213634 52535 213662 53784
rect 213778 53516 213806 53798
rect 213970 53516 213998 53798
rect 214162 53645 214190 53798
rect 214150 53639 214202 53645
rect 214150 53581 214202 53587
rect 213730 53488 213806 53516
rect 213922 53488 213998 53516
rect 213730 52947 213758 53488
rect 213716 52938 213772 52947
rect 213716 52873 213772 52882
rect 213922 52831 213950 53488
rect 213910 52825 213962 52831
rect 213910 52767 213962 52773
rect 213622 52529 213674 52535
rect 213622 52471 213674 52477
rect 213046 51641 213098 51647
rect 213046 51583 213098 51589
rect 214306 48983 214334 53798
rect 214498 53539 214526 53798
rect 214786 53645 214814 54025
rect 214774 53639 214826 53645
rect 214774 53581 214826 53587
rect 214484 53530 214540 53539
rect 214484 53465 214540 53474
rect 214978 51911 215006 54099
rect 632784 54080 632948 54108
rect 633120 54089 633374 54108
rect 633504 54105 633718 54108
rect 633504 54099 633770 54105
rect 633120 54083 633386 54089
rect 633120 54080 633334 54083
rect 632948 54057 633004 54066
rect 633504 54080 633758 54099
rect 633334 54025 633386 54031
rect 632566 54009 632618 54015
rect 628532 53974 628588 53983
rect 215808 53932 215870 53960
rect 628368 53932 628532 53960
rect 214964 51902 215020 51911
rect 214964 51837 215020 51846
rect 214294 48977 214346 48983
rect 214294 48919 214346 48925
rect 215074 48909 215102 53798
rect 215254 51567 215306 51573
rect 215254 51509 215306 51515
rect 215062 48903 215114 48909
rect 215062 48845 215114 48851
rect 215158 48903 215210 48909
rect 215158 48845 215210 48851
rect 211606 48237 211658 48243
rect 211606 48179 211658 48185
rect 211618 47873 211646 48179
rect 211606 47867 211658 47873
rect 211606 47809 211658 47815
rect 215170 46763 215198 48845
rect 215266 46763 215294 51509
rect 215458 48835 215486 53798
rect 215650 53645 215678 53798
rect 215638 53639 215690 53645
rect 215638 53581 215690 53587
rect 215842 53275 215870 53932
rect 631632 53941 631934 53960
rect 632400 53957 632566 53960
rect 632400 53951 632618 53957
rect 631632 53935 631946 53941
rect 631632 53932 631894 53935
rect 628532 53909 628588 53918
rect 632400 53932 632606 53951
rect 631894 53877 631946 53883
rect 629302 53861 629354 53867
rect 215986 53516 216014 53798
rect 216178 53516 216206 53798
rect 215986 53488 216062 53516
rect 215830 53269 215882 53275
rect 215830 53211 215882 53217
rect 215446 48829 215498 48835
rect 215446 48771 215498 48777
rect 216034 48169 216062 53488
rect 216130 53488 216206 53516
rect 216322 53784 216384 53812
rect 216130 48243 216158 53488
rect 216322 48983 216350 53784
rect 216310 48977 216362 48983
rect 216310 48919 216362 48925
rect 216118 48237 216170 48243
rect 216118 48179 216170 48185
rect 216022 48163 216074 48169
rect 216022 48105 216074 48111
rect 216514 48095 216542 53798
rect 216502 48089 216554 48095
rect 216502 48031 216554 48037
rect 216598 48089 216650 48095
rect 216598 48031 216650 48037
rect 209686 46757 209738 46763
rect 209686 46699 209738 46705
rect 215158 46757 215210 46763
rect 215158 46699 215210 46705
rect 215254 46757 215306 46763
rect 215254 46699 215306 46705
rect 209698 46435 209726 46699
rect 216610 46615 216638 48031
rect 216706 46615 216734 53798
rect 216898 48539 216926 53798
rect 217090 48803 217118 53798
rect 217076 48794 217132 48803
rect 217076 48729 217132 48738
rect 216886 48533 216938 48539
rect 216886 48475 216938 48481
rect 217282 48391 217310 53798
rect 217474 48951 217502 53798
rect 217460 48942 217516 48951
rect 217460 48877 217516 48886
rect 217666 48613 217694 53798
rect 217654 48607 217706 48613
rect 217654 48549 217706 48555
rect 217270 48385 217322 48391
rect 217270 48327 217322 48333
rect 217858 46911 217886 53798
rect 218016 53784 218078 53812
rect 218050 52503 218078 53784
rect 218194 53516 218222 53798
rect 218386 53516 218414 53798
rect 218194 53488 218270 53516
rect 218036 52494 218092 52503
rect 218036 52429 218092 52438
rect 218242 51763 218270 53488
rect 218338 53488 218414 53516
rect 218338 53095 218366 53488
rect 218324 53086 218380 53095
rect 218324 53021 218380 53030
rect 218722 52387 218750 53798
rect 218710 52381 218762 52387
rect 218710 52323 218762 52329
rect 218228 51754 218284 51763
rect 218228 51689 218284 51698
rect 219106 47873 219134 53798
rect 219094 47867 219146 47873
rect 219094 47809 219146 47815
rect 219490 47799 219518 53798
rect 219478 47793 219530 47799
rect 219478 47735 219530 47741
rect 219874 47577 219902 53798
rect 220224 53784 220286 53812
rect 220258 52651 220286 53784
rect 220594 53516 220622 53798
rect 220546 53488 220622 53516
rect 220546 52799 220574 53488
rect 220532 52790 220588 52799
rect 220532 52725 220588 52734
rect 220244 52642 220300 52651
rect 220244 52577 220300 52586
rect 219862 47571 219914 47577
rect 219862 47513 219914 47519
rect 217846 46905 217898 46911
rect 217846 46847 217898 46853
rect 216598 46609 216650 46615
rect 216598 46551 216650 46557
rect 216694 46609 216746 46615
rect 216694 46551 216746 46557
rect 220930 46541 220958 53798
rect 221314 52239 221342 53798
rect 221302 52233 221354 52239
rect 221302 52175 221354 52181
rect 221698 47947 221726 53798
rect 221686 47941 221738 47947
rect 221686 47883 221738 47889
rect 221782 46683 221834 46689
rect 221782 46625 221834 46631
rect 221794 46541 221822 46625
rect 220918 46535 220970 46541
rect 220918 46477 220970 46483
rect 221782 46535 221834 46541
rect 221782 46477 221834 46483
rect 209684 46426 209740 46435
rect 209684 46361 209740 46370
rect 222082 46171 222110 53798
rect 222178 53784 222432 53812
rect 222562 53784 222816 53812
rect 222178 46467 222206 53784
rect 222562 52461 222590 53784
rect 222550 52455 222602 52461
rect 222550 52397 222602 52403
rect 223138 46763 223166 53798
rect 223522 52313 223550 53798
rect 223510 52307 223562 52313
rect 223510 52249 223562 52255
rect 223126 46757 223178 46763
rect 223126 46699 223178 46705
rect 222166 46461 222218 46467
rect 222166 46403 222218 46409
rect 223906 46245 223934 53798
rect 224290 52165 224318 53798
rect 224640 53784 224702 53812
rect 224278 52159 224330 52165
rect 224278 52101 224330 52107
rect 224674 46393 224702 53784
rect 224770 53784 225024 53812
rect 224770 48095 224798 53784
rect 224758 48089 224810 48095
rect 224758 48031 224810 48037
rect 224662 46387 224714 46393
rect 224662 46329 224714 46335
rect 225346 46319 225374 53798
rect 225730 49797 225758 53798
rect 226114 49871 226142 53798
rect 226102 49865 226154 49871
rect 226102 49807 226154 49813
rect 225718 49791 225770 49797
rect 225718 49733 225770 49739
rect 226498 49575 226526 53798
rect 226594 53784 226848 53812
rect 226978 53784 227232 53812
rect 226486 49569 226538 49575
rect 226486 49511 226538 49517
rect 226594 48909 226622 53784
rect 226978 49945 227006 53784
rect 227554 50315 227582 53798
rect 227938 53127 227966 53798
rect 227926 53121 227978 53127
rect 227926 53063 227978 53069
rect 227542 50309 227594 50315
rect 227542 50251 227594 50257
rect 226966 49939 227018 49945
rect 226966 49881 227018 49887
rect 226582 48903 226634 48909
rect 226582 48845 226634 48851
rect 228322 46541 228350 53798
rect 228706 50167 228734 53798
rect 228802 53784 229056 53812
rect 229186 53784 229440 53812
rect 228802 50241 228830 53784
rect 228790 50235 228842 50241
rect 228790 50177 228842 50183
rect 228694 50161 228746 50167
rect 228694 50103 228746 50109
rect 229186 50093 229214 53784
rect 229174 50087 229226 50093
rect 229174 50029 229226 50035
rect 229762 47651 229790 53798
rect 230146 50019 230174 53798
rect 230134 50013 230186 50019
rect 230134 49955 230186 49961
rect 230530 48021 230558 53798
rect 230914 50759 230942 53798
rect 231010 53784 231264 53812
rect 231394 53784 231648 53812
rect 230902 50753 230954 50759
rect 230902 50695 230954 50701
rect 231010 50537 231038 53784
rect 230998 50531 231050 50537
rect 230998 50473 231050 50479
rect 231394 50389 231422 53784
rect 231382 50383 231434 50389
rect 231382 50325 231434 50331
rect 230518 48015 230570 48021
rect 230518 47957 230570 47963
rect 231970 47725 231998 53798
rect 232354 50611 232382 53798
rect 232738 50685 232766 53798
rect 232726 50679 232778 50685
rect 232726 50621 232778 50627
rect 232342 50605 232394 50611
rect 232342 50547 232394 50553
rect 233122 50463 233150 53798
rect 233314 53784 233472 53812
rect 233602 53784 233856 53812
rect 233110 50457 233162 50463
rect 233110 50399 233162 50405
rect 231958 47719 232010 47725
rect 231958 47661 232010 47667
rect 229750 47645 229802 47651
rect 229750 47587 229802 47593
rect 233314 46837 233342 53784
rect 233602 47429 233630 53784
rect 234178 51055 234206 53798
rect 234562 51129 234590 53798
rect 234550 51123 234602 51129
rect 234550 51065 234602 51071
rect 234166 51049 234218 51055
rect 234166 50991 234218 50997
rect 234946 50981 234974 53798
rect 234934 50975 234986 50981
rect 234934 50917 234986 50923
rect 235330 50833 235358 53798
rect 235426 53784 235680 53812
rect 235810 53784 236064 53812
rect 235318 50827 235370 50833
rect 235318 50769 235370 50775
rect 235426 48465 235454 53784
rect 235810 50907 235838 53784
rect 236386 51277 236414 53798
rect 236374 51271 236426 51277
rect 236374 51213 236426 51219
rect 235798 50901 235850 50907
rect 235798 50843 235850 50849
rect 235414 48459 235466 48465
rect 235414 48401 235466 48407
rect 236770 47915 236798 53798
rect 237154 51351 237182 53798
rect 237142 51345 237194 51351
rect 237142 51287 237194 51293
rect 237538 51203 237566 53798
rect 237634 53784 237888 53812
rect 238018 53784 238272 53812
rect 237526 51197 237578 51203
rect 237526 51139 237578 51145
rect 237634 49205 237662 53784
rect 238018 51425 238046 53784
rect 238006 51419 238058 51425
rect 238006 51361 238058 51367
rect 237622 49199 237674 49205
rect 237622 49141 237674 49147
rect 238594 48063 238622 53798
rect 238978 49353 239006 53798
rect 238966 49347 239018 49353
rect 238966 49289 239018 49295
rect 239362 48211 239390 53798
rect 239746 49649 239774 53798
rect 239842 53784 240096 53812
rect 240226 53784 240480 53812
rect 239842 51171 239870 53784
rect 239828 51162 239884 51171
rect 239828 51097 239884 51106
rect 239734 49643 239786 49649
rect 239734 49585 239786 49591
rect 239348 48202 239404 48211
rect 239348 48137 239404 48146
rect 238580 48054 238636 48063
rect 238580 47989 238636 47998
rect 236756 47906 236812 47915
rect 236756 47841 236812 47850
rect 240226 47619 240254 53784
rect 240802 49279 240830 53798
rect 241186 49501 241214 53798
rect 241174 49495 241226 49501
rect 241174 49437 241226 49443
rect 240790 49273 240842 49279
rect 240790 49215 240842 49221
rect 241570 47767 241598 53798
rect 241954 49723 241982 53798
rect 242050 53784 242304 53812
rect 242434 53784 242688 53812
rect 242050 51023 242078 53784
rect 242036 51014 242092 51023
rect 242036 50949 242092 50958
rect 241942 49717 241994 49723
rect 241942 49659 241994 49665
rect 242434 48359 242462 53784
rect 243010 51319 243038 53798
rect 242996 51310 243052 51319
rect 242996 51245 243052 51254
rect 243394 48507 243422 53798
rect 243778 48655 243806 53798
rect 244162 50875 244190 53798
rect 244148 50866 244204 50875
rect 244148 50801 244204 50810
rect 264884 50422 264940 50431
rect 264884 50357 264940 50366
rect 264898 48983 264926 50357
rect 627202 48983 627230 53798
rect 627600 53784 627806 53812
rect 627778 53497 627806 53784
rect 627766 53491 627818 53497
rect 627766 53433 627818 53439
rect 264886 48977 264938 48983
rect 264886 48919 264938 48925
rect 627190 48977 627242 48983
rect 627190 48919 627242 48925
rect 243764 48646 243820 48655
rect 243764 48581 243820 48590
rect 243380 48498 243436 48507
rect 243380 48433 243436 48442
rect 242420 48350 242476 48359
rect 242420 48285 242476 48294
rect 241556 47758 241612 47767
rect 627970 47725 627998 53798
rect 628704 53784 628958 53812
rect 629088 53809 629302 53812
rect 630644 53826 630700 53835
rect 629088 53803 629354 53809
rect 629088 53784 629342 53803
rect 629808 53784 630110 53812
rect 630192 53793 630398 53812
rect 630192 53787 630410 53793
rect 630192 53784 630358 53787
rect 628930 48317 628958 53784
rect 630082 53719 630110 53784
rect 630576 53784 630644 53812
rect 630912 53784 631166 53812
rect 631296 53784 631550 53812
rect 630644 53761 630700 53770
rect 630358 53729 630410 53735
rect 630070 53713 630122 53719
rect 630070 53655 630122 53661
rect 631138 53571 631166 53784
rect 631522 53645 631550 53784
rect 631510 53639 631562 53645
rect 631510 53581 631562 53587
rect 631126 53565 631178 53571
rect 631126 53507 631178 53513
rect 634114 52091 634142 222948
rect 639668 222398 639724 222407
rect 639668 222333 639724 222342
rect 639380 221806 639436 221815
rect 639380 221741 639436 221750
rect 635254 92859 635306 92865
rect 635254 92801 635306 92807
rect 635062 92785 635114 92791
rect 635062 92727 635114 92733
rect 634966 92563 635018 92569
rect 634966 92505 635018 92511
rect 634774 76505 634826 76511
rect 634774 76447 634826 76453
rect 634786 53867 634814 76447
rect 634870 76431 634922 76437
rect 634870 76373 634922 76379
rect 634882 53983 634910 76373
rect 634978 54237 635006 92505
rect 635074 54279 635102 92727
rect 635158 92415 635210 92421
rect 635158 92357 635210 92363
rect 635060 54270 635116 54279
rect 634966 54231 635018 54237
rect 635060 54205 635116 54214
rect 634966 54173 635018 54179
rect 634868 53974 634924 53983
rect 634868 53909 634924 53918
rect 634774 53861 634826 53867
rect 634774 53803 634826 53809
rect 635170 53719 635198 92357
rect 635266 53793 635294 92801
rect 635350 92637 635402 92643
rect 635350 92579 635402 92585
rect 635362 54427 635390 92579
rect 635446 92489 635498 92495
rect 635446 92431 635498 92437
rect 635348 54418 635404 54427
rect 635348 54353 635404 54362
rect 635458 53941 635486 92431
rect 635542 87827 635594 87833
rect 635542 87769 635594 87775
rect 635446 53935 635498 53941
rect 635446 53877 635498 53883
rect 635254 53787 635306 53793
rect 635254 53729 635306 53735
rect 635158 53713 635210 53719
rect 635158 53655 635210 53661
rect 634102 52085 634154 52091
rect 634102 52027 634154 52033
rect 628918 48311 628970 48317
rect 628918 48253 628970 48259
rect 241556 47693 241612 47702
rect 627958 47719 628010 47725
rect 627958 47661 628010 47667
rect 240212 47610 240268 47619
rect 240212 47545 240268 47554
rect 233590 47423 233642 47429
rect 233590 47365 233642 47371
rect 233302 46831 233354 46837
rect 233302 46773 233354 46779
rect 228310 46535 228362 46541
rect 228310 46477 228362 46483
rect 225334 46313 225386 46319
rect 225334 46255 225386 46261
rect 223894 46239 223946 46245
rect 223894 46181 223946 46187
rect 222070 46165 222122 46171
rect 222070 46107 222122 46113
rect 403126 45203 403178 45209
rect 403126 45145 403178 45151
rect 209590 44759 209642 44765
rect 209590 44701 209642 44707
rect 208820 44650 208876 44659
rect 208820 44585 208876 44594
rect 302516 43318 302572 43327
rect 302516 43253 302572 43262
rect 306740 43318 306796 43327
rect 306740 43253 306796 43262
rect 361748 43318 361804 43327
rect 361748 43253 361804 43262
rect 364916 43318 364972 43327
rect 364916 43253 364972 43262
rect 302530 42120 302558 43253
rect 306754 42120 306782 43253
rect 357140 43170 357196 43179
rect 357140 43105 357196 43114
rect 310102 42391 310154 42397
rect 310102 42333 310154 42339
rect 302530 42092 302688 42120
rect 306754 42092 307008 42120
rect 310114 42106 310142 42333
rect 357154 42120 357182 43105
rect 357154 42092 357456 42120
rect 361762 42106 361790 43253
rect 364930 42106 364958 43253
rect 403138 41953 403166 45145
rect 408886 45129 408938 45135
rect 408886 45071 408938 45077
rect 406294 45055 406346 45061
rect 406294 44997 406346 45003
rect 405238 42169 405290 42175
rect 405290 42117 405552 42120
rect 405238 42111 405552 42117
rect 405250 42092 405552 42111
rect 403126 41947 403178 41953
rect 403126 41889 403178 41895
rect 406306 41847 406334 44997
rect 408898 42143 408926 45071
rect 446518 44981 446570 44987
rect 446518 44923 446570 44929
rect 408884 42134 408940 42143
rect 408884 42069 408940 42078
rect 416276 42134 416332 42143
rect 416332 42092 416592 42120
rect 416276 42069 416332 42078
rect 406292 41838 406348 41847
rect 406292 41773 406348 41782
rect 410804 41838 410860 41847
rect 410860 41796 411120 41824
rect 410804 41773 410860 41782
rect 208438 41725 208490 41731
rect 208438 41667 208490 41673
rect 204884 40802 204940 40811
rect 204884 40737 204940 40746
rect 138164 40210 138220 40219
rect 138164 40145 138220 40154
rect 446530 37439 446558 44923
rect 499990 44907 500042 44913
rect 499990 44849 500042 44855
rect 465620 44798 465676 44807
rect 465620 44733 465676 44742
rect 460066 42101 460368 42120
rect 460054 42095 460368 42101
rect 460106 42092 460368 42095
rect 460054 42037 460106 42043
rect 459190 42021 459242 42027
rect 459190 41963 459242 41969
rect 463702 42021 463754 42027
rect 463754 41969 464016 41972
rect 463702 41963 464016 41969
rect 459202 37439 459230 41963
rect 463714 41944 464016 41963
rect 465634 41824 465662 44733
rect 471092 42134 471148 42143
rect 471148 42092 471408 42120
rect 471092 42069 471148 42078
rect 465634 41796 465936 41824
rect 500002 40399 500030 44849
rect 508246 44833 508298 44839
rect 508246 44775 508298 44781
rect 508258 43285 508286 44775
rect 523894 44759 523946 44765
rect 523894 44701 523946 44707
rect 521206 44685 521258 44691
rect 521206 44627 521258 44633
rect 521588 44650 521644 44659
rect 508246 43279 508298 43285
rect 508246 43221 508298 43227
rect 520342 43205 520394 43211
rect 520342 43147 520394 43153
rect 520354 42120 520382 43147
rect 521218 42143 521246 44627
rect 521588 44585 521644 44594
rect 521204 42134 521260 42143
rect 520354 42092 520656 42120
rect 521602 42120 521630 44585
rect 523906 43179 523934 44701
rect 635554 44691 635582 87769
rect 635638 83683 635690 83689
rect 635638 83625 635690 83631
rect 635650 53645 635678 83625
rect 635734 83609 635786 83615
rect 635734 83551 635786 83557
rect 635638 53639 635690 53645
rect 635638 53581 635690 53587
rect 635746 53497 635774 83551
rect 635926 80797 635978 80803
rect 635926 80739 635978 80745
rect 635830 80723 635882 80729
rect 635830 80665 635882 80671
rect 635842 54015 635870 80665
rect 635830 54009 635882 54015
rect 635830 53951 635882 53957
rect 635938 53571 635966 80739
rect 636310 76801 636362 76807
rect 636310 76743 636362 76749
rect 636022 76727 636074 76733
rect 636022 76669 636074 76675
rect 636034 54089 636062 76669
rect 636214 76653 636266 76659
rect 636214 76595 636266 76601
rect 636118 76579 636170 76585
rect 636118 76521 636170 76527
rect 636022 54083 636074 54089
rect 636022 54025 636074 54031
rect 635926 53565 635978 53571
rect 635926 53507 635978 53513
rect 635734 53491 635786 53497
rect 635734 53433 635786 53439
rect 636130 48983 636158 76521
rect 636226 54163 636254 76595
rect 636214 54157 636266 54163
rect 636214 54099 636266 54105
rect 636322 53835 636350 76743
rect 636406 76357 636458 76363
rect 636406 76299 636458 76305
rect 636418 54131 636446 76299
rect 636404 54122 636460 54131
rect 636404 54057 636460 54066
rect 636308 53826 636364 53835
rect 636308 53761 636364 53770
rect 636118 48977 636170 48983
rect 636118 48919 636170 48925
rect 639394 48169 639422 221741
rect 639574 195867 639626 195873
rect 639574 195809 639626 195815
rect 639586 54681 639614 195809
rect 639574 54675 639626 54681
rect 639574 54617 639626 54623
rect 639682 51943 639710 222333
rect 640738 221815 640766 256341
rect 642260 255698 642316 255707
rect 642260 255633 642262 255642
rect 642314 255633 642316 255642
rect 642262 255601 642314 255607
rect 649474 229469 649502 927373
rect 649570 846079 649598 989755
rect 649750 980859 649802 980865
rect 649750 980801 649802 980807
rect 649556 846070 649612 846079
rect 649556 846005 649612 846014
rect 649558 748869 649610 748875
rect 649558 748811 649610 748817
rect 649570 229543 649598 748811
rect 649654 702767 649706 702773
rect 649654 702709 649706 702715
rect 649558 229537 649610 229543
rect 649558 229479 649610 229485
rect 649462 229463 649514 229469
rect 649462 229405 649514 229411
rect 649666 222439 649694 702709
rect 649762 676873 649790 980801
rect 649858 752099 649886 990643
rect 649942 989369 649994 989375
rect 649942 989311 649994 989317
rect 649954 799163 649982 989311
rect 650050 892847 650078 994005
rect 650902 992181 650954 992187
rect 650902 992123 650954 992129
rect 650134 984929 650186 984935
rect 650134 984871 650186 984877
rect 650036 892838 650092 892847
rect 650036 892773 650092 892782
rect 649940 799154 649996 799163
rect 649940 799089 649996 799098
rect 649844 752090 649900 752099
rect 649844 752025 649900 752034
rect 650146 705331 650174 984871
rect 650132 705322 650188 705331
rect 650132 705257 650188 705266
rect 649750 676867 649802 676873
rect 649750 676809 649802 676815
rect 649750 656739 649802 656745
rect 649750 656681 649802 656687
rect 649762 229099 649790 656681
rect 649846 613523 649898 613529
rect 649846 613465 649898 613471
rect 649858 229617 649886 613465
rect 649942 567421 649994 567427
rect 649942 567363 649994 567369
rect 649846 229611 649898 229617
rect 649846 229553 649898 229559
rect 649954 229173 649982 567363
rect 650038 521319 650090 521325
rect 650038 521261 650090 521267
rect 649942 229167 649994 229173
rect 649942 229109 649994 229115
rect 649750 229093 649802 229099
rect 649750 229035 649802 229041
rect 641014 222433 641066 222439
rect 641012 222398 641014 222407
rect 649654 222433 649706 222439
rect 641066 222398 641068 222407
rect 649654 222375 649706 222381
rect 641012 222333 641068 222342
rect 640724 221806 640780 221815
rect 640724 221741 640780 221750
rect 641302 221397 641354 221403
rect 639860 221362 639916 221371
rect 639860 221297 639916 221306
rect 641300 221362 641302 221371
rect 641354 221362 641356 221371
rect 641300 221297 641356 221306
rect 639764 211002 639820 211011
rect 639764 210937 639820 210946
rect 639778 210303 639806 210937
rect 639766 210297 639818 210303
rect 639766 210239 639818 210245
rect 639778 52017 639806 210239
rect 639766 52011 639818 52017
rect 639766 51953 639818 51959
rect 639670 51937 639722 51943
rect 639670 51879 639722 51885
rect 639382 48163 639434 48169
rect 639382 48105 639434 48111
rect 639874 46615 639902 221297
rect 650050 220811 650078 521261
rect 650134 478177 650186 478183
rect 650134 478119 650186 478125
rect 650146 229247 650174 478119
rect 650230 391745 650282 391751
rect 650230 391687 650282 391693
rect 650242 229321 650270 391687
rect 650326 345643 650378 345649
rect 650326 345585 650378 345591
rect 650230 229315 650282 229321
rect 650230 229257 650282 229263
rect 650134 229241 650186 229247
rect 650134 229183 650186 229189
rect 650338 221403 650366 345585
rect 650422 299615 650474 299621
rect 650422 299557 650474 299563
rect 650434 229395 650462 299557
rect 650422 229389 650474 229395
rect 650422 229331 650474 229337
rect 650914 229025 650942 992123
rect 652246 983671 652298 983677
rect 652246 983613 652298 983619
rect 652258 939129 652286 983613
rect 652342 983597 652394 983603
rect 652342 983539 652394 983545
rect 652354 943199 652382 983539
rect 652438 983523 652490 983529
rect 652438 983465 652490 983471
rect 652342 943193 652394 943199
rect 652342 943135 652394 943141
rect 652450 941941 652478 983465
rect 673942 980711 673994 980717
rect 673942 980653 673994 980659
rect 655124 974386 655180 974395
rect 655124 974321 655180 974330
rect 653686 953331 653738 953337
rect 653686 953273 653738 953279
rect 653698 947436 653726 953273
rect 654356 951002 654412 951011
rect 654356 950937 654412 950946
rect 653698 947408 653822 947436
rect 652438 941935 652490 941941
rect 652438 941877 652490 941883
rect 653794 939319 653822 947408
rect 654370 942089 654398 950937
rect 655138 944679 655166 974321
rect 673954 967587 673982 980653
rect 674518 980637 674570 980643
rect 674518 980579 674570 980585
rect 673940 967578 673996 967587
rect 673940 967513 673996 967522
rect 655220 962694 655276 962703
rect 655220 962629 655276 962638
rect 655234 944901 655262 962629
rect 674530 960573 674558 980579
rect 675106 966722 675408 966750
rect 675106 965663 675134 966722
rect 675778 965663 675806 966070
rect 675092 965654 675148 965663
rect 675092 965589 675148 965598
rect 675764 965654 675820 965663
rect 675764 965589 675820 965598
rect 675106 965421 675408 965449
rect 675106 964923 675134 965421
rect 675092 964914 675148 964923
rect 675092 964849 675148 964858
rect 675106 963581 675408 963609
rect 675106 962851 675134 963581
rect 675202 963022 675408 963050
rect 675092 962842 675148 962851
rect 675092 962777 675148 962786
rect 675202 962555 675230 963022
rect 675188 962546 675244 962555
rect 675188 962481 675244 962490
rect 675394 962259 675422 962399
rect 675380 962250 675436 962259
rect 675380 962185 675436 962194
rect 675778 961519 675806 961778
rect 675764 961510 675820 961519
rect 675764 961445 675820 961454
rect 675490 961075 675518 961186
rect 675476 961066 675532 961075
rect 675476 961001 675532 961010
rect 674530 960559 675696 960573
rect 674530 960545 675710 960559
rect 675682 960187 675710 960545
rect 675668 960178 675724 960187
rect 675668 960113 675724 960122
rect 675490 959035 675518 959262
rect 673942 959029 673994 959035
rect 673942 958971 673994 958977
rect 675478 959029 675530 959035
rect 675478 958971 675530 958977
rect 669526 954737 669578 954743
rect 669526 954679 669578 954685
rect 655222 944895 655274 944901
rect 655222 944837 655274 944843
rect 655126 944673 655178 944679
rect 655126 944615 655178 944621
rect 654358 942083 654410 942089
rect 654358 942025 654410 942031
rect 653780 939310 653836 939319
rect 653780 939245 653836 939254
rect 652246 939123 652298 939129
rect 652246 939065 652298 939071
rect 654454 927505 654506 927511
rect 654452 927470 654454 927479
rect 666742 927505 666794 927511
rect 654506 927470 654508 927479
rect 666742 927447 666794 927453
rect 654452 927405 654508 927414
rect 654452 915778 654508 915787
rect 654452 915713 654508 915722
rect 654466 913007 654494 915713
rect 654454 913001 654506 913007
rect 654454 912943 654506 912949
rect 660982 913001 661034 913007
rect 660982 912943 661034 912949
rect 654452 904086 654508 904095
rect 654452 904021 654508 904030
rect 654466 901537 654494 904021
rect 654454 901531 654506 901537
rect 654454 901473 654506 901479
rect 654452 880554 654508 880563
rect 654452 880489 654508 880498
rect 654466 878449 654494 880489
rect 654454 878443 654506 878449
rect 654454 878385 654506 878391
rect 660886 878443 660938 878449
rect 660886 878385 660938 878391
rect 654452 868862 654508 868871
rect 654452 868797 654508 868806
rect 654466 867349 654494 868797
rect 654454 867343 654506 867349
rect 654454 867285 654506 867291
rect 654452 857170 654508 857179
rect 654452 857105 654508 857114
rect 654466 855435 654494 857105
rect 654454 855429 654506 855435
rect 654454 855371 654506 855377
rect 654452 833638 654508 833647
rect 654452 833573 654508 833582
rect 654466 832421 654494 833573
rect 654454 832415 654506 832421
rect 654454 832357 654506 832363
rect 654452 821946 654508 821955
rect 654452 821881 654508 821890
rect 654466 820877 654494 821881
rect 654454 820871 654506 820877
rect 654454 820813 654506 820819
rect 654452 810254 654508 810263
rect 654452 810189 654508 810198
rect 654466 809333 654494 810189
rect 654454 809327 654506 809333
rect 654454 809269 654506 809275
rect 654452 786722 654508 786731
rect 654452 786657 654508 786666
rect 654466 786319 654494 786657
rect 654454 786313 654506 786319
rect 654454 786255 654506 786261
rect 654452 775030 654508 775039
rect 654452 774965 654508 774974
rect 654466 774775 654494 774965
rect 654454 774769 654506 774775
rect 654454 774711 654506 774717
rect 654452 763338 654508 763347
rect 654452 763273 654454 763282
rect 654506 763273 654508 763282
rect 654454 763241 654506 763247
rect 654452 739806 654508 739815
rect 654452 739741 654508 739750
rect 654466 737331 654494 739741
rect 654454 737325 654506 737331
rect 654454 737267 654506 737273
rect 655124 728114 655180 728123
rect 655124 728049 655180 728058
rect 654452 716274 654508 716283
rect 654452 716209 654508 716218
rect 654466 714317 654494 716209
rect 654454 714311 654506 714317
rect 654454 714253 654506 714259
rect 654836 692890 654892 692899
rect 654836 692825 654892 692834
rect 654850 691303 654878 692825
rect 654838 691297 654890 691303
rect 654838 691239 654890 691245
rect 653686 676867 653738 676873
rect 653686 676809 653738 676815
rect 653698 673932 653726 676809
rect 653698 673904 653822 673932
rect 653794 658415 653822 673904
rect 654452 669358 654508 669367
rect 654452 669293 654508 669302
rect 654466 668215 654494 669293
rect 654454 668209 654506 668215
rect 654454 668151 654506 668157
rect 653780 658406 653836 658415
rect 653780 658341 653836 658350
rect 654452 645974 654508 645983
rect 654452 645909 654508 645918
rect 654466 645201 654494 645909
rect 654454 645195 654506 645201
rect 654454 645137 654506 645143
rect 654452 622442 654508 622451
rect 654452 622377 654508 622386
rect 654466 622113 654494 622377
rect 654454 622107 654506 622113
rect 654454 622049 654506 622055
rect 654454 613449 654506 613455
rect 654454 613391 654506 613397
rect 654466 610759 654494 613391
rect 654452 610750 654508 610759
rect 654452 610685 654508 610694
rect 654452 599354 654508 599363
rect 654452 599289 654508 599298
rect 654466 599099 654494 599289
rect 654454 599093 654506 599099
rect 654454 599035 654506 599041
rect 654452 587218 654508 587227
rect 654452 587153 654508 587162
rect 654466 585113 654494 587153
rect 654454 585107 654506 585113
rect 654454 585049 654506 585055
rect 655138 584817 655166 728049
rect 660898 721939 660926 878385
rect 660994 767819 661022 912943
rect 663958 901531 664010 901537
rect 663958 901473 664010 901479
rect 663766 867343 663818 867349
rect 663766 867285 663818 867291
rect 661174 855429 661226 855435
rect 661174 855371 661226 855377
rect 660982 767813 661034 767819
rect 660982 767755 661034 767761
rect 661078 763299 661130 763305
rect 661078 763241 661130 763247
rect 660982 737399 661034 737405
rect 660982 737341 661034 737347
rect 660886 721933 660938 721939
rect 660886 721875 660938 721881
rect 655316 681198 655372 681207
rect 655316 681133 655372 681142
rect 655220 634282 655276 634291
rect 655220 634217 655276 634226
rect 655126 584811 655178 584817
rect 655126 584753 655178 584759
rect 654452 575526 654508 575535
rect 654452 575461 654508 575470
rect 654466 573199 654494 575461
rect 654454 573193 654506 573199
rect 654454 573135 654506 573141
rect 654454 564461 654506 564467
rect 654454 564403 654506 564409
rect 654466 563843 654494 564403
rect 654452 563834 654508 563843
rect 654452 563769 654508 563778
rect 654452 552142 654508 552151
rect 654452 552077 654508 552086
rect 654466 550185 654494 552077
rect 654454 550179 654506 550185
rect 654454 550121 654506 550127
rect 655124 540302 655180 540311
rect 655124 540237 655180 540246
rect 654452 528610 654508 528619
rect 654452 528545 654508 528554
rect 654466 527097 654494 528545
rect 654454 527091 654506 527097
rect 654454 527033 654506 527039
rect 654454 517989 654506 517995
rect 654454 517931 654506 517937
rect 654466 516927 654494 517931
rect 654452 516918 654508 516927
rect 654452 516853 654508 516862
rect 654452 505226 654508 505235
rect 654452 505161 654508 505170
rect 654466 504083 654494 505161
rect 654454 504077 654506 504083
rect 654454 504019 654506 504025
rect 654452 493386 654508 493395
rect 654452 493321 654508 493330
rect 654466 492539 654494 493321
rect 654454 492533 654506 492539
rect 654454 492475 654506 492481
rect 654452 481694 654508 481703
rect 654452 481629 654508 481638
rect 654466 480995 654494 481629
rect 654454 480989 654506 480995
rect 654454 480931 654506 480937
rect 654454 470037 654506 470043
rect 654452 470002 654454 470011
rect 654506 470002 654508 470011
rect 654452 469937 654508 469946
rect 654356 458310 654412 458319
rect 654356 458245 654412 458254
rect 654370 457981 654398 458245
rect 654358 457975 654410 457981
rect 654358 457917 654410 457923
rect 654452 446470 654508 446479
rect 654452 446405 654454 446414
rect 654506 446405 654508 446414
rect 654454 446373 654506 446379
rect 654356 434778 654412 434787
rect 654356 434713 654412 434722
rect 654370 432081 654398 434713
rect 654358 432075 654410 432081
rect 654358 432017 654410 432023
rect 654454 423343 654506 423349
rect 654454 423285 654506 423291
rect 654466 423095 654494 423285
rect 654452 423086 654508 423095
rect 654452 423021 654508 423030
rect 655028 411246 655084 411255
rect 655028 411181 655084 411190
rect 655042 408993 655070 411181
rect 655030 408987 655082 408993
rect 655030 408929 655082 408935
rect 654452 399554 654508 399563
rect 654452 399489 654508 399498
rect 654466 397523 654494 399489
rect 654454 397517 654506 397523
rect 654454 397459 654506 397465
rect 653876 387862 653932 387871
rect 653876 387797 653932 387806
rect 653890 385979 653918 387797
rect 653878 385973 653930 385979
rect 653878 385915 653930 385921
rect 654166 377241 654218 377247
rect 654166 377183 654218 377189
rect 654178 376179 654206 377183
rect 654164 376170 654220 376179
rect 654164 376105 654220 376114
rect 654452 364330 654508 364339
rect 654452 364265 654508 364274
rect 654466 363409 654494 364265
rect 654454 363403 654506 363409
rect 654454 363345 654506 363351
rect 655138 363113 655166 540237
rect 655234 495573 655262 634217
rect 655330 541527 655358 681133
rect 660886 555877 660938 555883
rect 660886 555819 660938 555825
rect 655318 541521 655370 541527
rect 655318 541463 655370 541469
rect 655222 495567 655274 495573
rect 655222 495509 655274 495515
rect 655126 363107 655178 363113
rect 655126 363049 655178 363055
rect 655316 352638 655372 352647
rect 655316 352573 655372 352582
rect 654164 340946 654220 340955
rect 654164 340881 654220 340890
rect 654178 339877 654206 340881
rect 654166 339871 654218 339877
rect 654166 339813 654218 339819
rect 653974 329807 654026 329813
rect 653974 329749 654026 329755
rect 653986 329263 654014 329749
rect 653972 329254 654028 329263
rect 653972 329189 654028 329198
rect 655124 317414 655180 317423
rect 655124 317349 655180 317358
rect 653782 282447 653834 282453
rect 653782 282389 653834 282395
rect 653794 282347 653822 282389
rect 653780 282338 653836 282347
rect 653780 282273 653836 282282
rect 650902 229019 650954 229025
rect 650902 228961 650954 228967
rect 650326 221397 650378 221403
rect 650326 221339 650378 221345
rect 641302 220805 641354 220811
rect 639956 220770 640012 220779
rect 639956 220705 640012 220714
rect 641300 220770 641302 220779
rect 650038 220805 650090 220811
rect 641354 220770 641356 220779
rect 650038 220747 650090 220753
rect 641300 220705 641356 220714
rect 639970 195873 639998 220705
rect 639958 195867 640010 195873
rect 639958 195809 640010 195815
rect 641494 167229 641546 167235
rect 641494 167171 641546 167177
rect 641506 165871 641534 167171
rect 642068 166898 642124 166907
rect 642068 166833 642124 166842
rect 641492 165862 641548 165871
rect 641492 165797 641548 165806
rect 642082 164201 642110 166833
rect 642164 166454 642220 166463
rect 642164 166389 642220 166398
rect 642178 164275 642206 166389
rect 642166 164269 642218 164275
rect 642166 164211 642218 164217
rect 642070 164195 642122 164201
rect 642070 164137 642122 164143
rect 640148 150026 640204 150035
rect 640148 149961 640204 149970
rect 640162 149845 640190 149961
rect 640150 149839 640202 149845
rect 640150 149781 640202 149787
rect 643606 149839 643658 149845
rect 643606 149781 643658 149787
rect 642164 143514 642220 143523
rect 642164 143449 642220 143458
rect 642178 142593 642206 143449
rect 642166 142587 642218 142593
rect 642166 142529 642218 142535
rect 640726 135409 640778 135415
rect 640726 135351 640778 135357
rect 640738 120139 640766 135351
rect 643618 132529 643646 149781
rect 655138 138449 655166 317349
rect 655220 305722 655276 305731
rect 655220 305657 655276 305666
rect 655234 138597 655262 305657
rect 655330 184403 655358 352573
rect 655412 294030 655468 294039
rect 655412 293965 655468 293974
rect 655318 184397 655370 184403
rect 655318 184339 655370 184345
rect 655222 138591 655274 138597
rect 655222 138533 655274 138539
rect 655126 138443 655178 138449
rect 655126 138385 655178 138391
rect 655426 135637 655454 293965
rect 660898 282453 660926 555819
rect 660994 470043 661022 737341
rect 661090 630623 661118 763241
rect 661186 720903 661214 855371
rect 663778 722531 663806 867285
rect 663862 780541 663914 780547
rect 663862 780483 663914 780489
rect 663766 722525 663818 722531
rect 663766 722467 663818 722473
rect 661174 720897 661226 720903
rect 661174 720839 661226 720845
rect 661270 668209 661322 668215
rect 661270 668151 661322 668157
rect 661078 630617 661130 630623
rect 661078 630559 661130 630565
rect 661174 585107 661226 585113
rect 661174 585049 661226 585055
rect 661078 550179 661130 550185
rect 661078 550121 661130 550127
rect 660982 470037 661034 470043
rect 660982 469979 661034 469985
rect 660982 457975 661034 457981
rect 660982 457917 661034 457923
rect 660886 282447 660938 282453
rect 660886 282389 660938 282395
rect 660994 274091 661022 457917
rect 661090 363927 661118 550121
rect 661186 409955 661214 585049
rect 661282 540787 661310 668151
rect 663766 602127 663818 602133
rect 663766 602069 663818 602075
rect 661270 540781 661322 540787
rect 661270 540723 661322 540729
rect 661174 409949 661226 409955
rect 661174 409891 661226 409897
rect 661078 363921 661130 363927
rect 661078 363863 661130 363869
rect 661174 363403 661226 363409
rect 661174 363345 661226 363351
rect 660982 274085 661034 274091
rect 660982 274027 661034 274033
rect 661186 183959 661214 363345
rect 663778 329813 663806 602069
rect 663874 517995 663902 780483
rect 663970 765895 663998 901473
rect 666646 865345 666698 865351
rect 666646 865287 666698 865293
rect 664054 809327 664106 809333
rect 664054 809269 664106 809275
rect 663958 765889 664010 765895
rect 663958 765831 664010 765837
rect 663958 737325 664010 737331
rect 663958 737267 664010 737273
rect 663970 586371 663998 737267
rect 664066 675911 664094 809269
rect 664150 714311 664202 714317
rect 664150 714253 664202 714259
rect 664054 675905 664106 675911
rect 664054 675847 664106 675853
rect 663958 586365 664010 586371
rect 663958 586307 664010 586313
rect 664162 585483 664190 714253
rect 664150 585477 664202 585483
rect 664150 585419 664202 585425
rect 663958 573193 664010 573199
rect 663958 573135 664010 573141
rect 663862 517989 663914 517995
rect 663862 517931 663914 517937
rect 663862 492533 663914 492539
rect 663862 492475 663914 492481
rect 663766 329807 663818 329813
rect 663766 329749 663818 329755
rect 663874 319971 663902 492475
rect 663970 408475 663998 573135
rect 666658 564467 666686 865287
rect 666754 766931 666782 927447
rect 667030 820871 667082 820877
rect 667030 820813 667082 820819
rect 666838 786313 666890 786319
rect 666838 786255 666890 786261
rect 666742 766925 666794 766931
rect 666742 766867 666794 766873
rect 666742 645269 666794 645275
rect 666742 645211 666794 645217
rect 666646 564461 666698 564467
rect 666646 564403 666698 564409
rect 666646 504077 666698 504083
rect 666646 504019 666698 504025
rect 664054 432075 664106 432081
rect 664054 432017 664106 432023
rect 663958 408469 664010 408475
rect 663958 408411 664010 408417
rect 663958 397517 664010 397523
rect 663958 397459 664010 397465
rect 663862 319965 663914 319971
rect 663862 319907 663914 319913
rect 662326 255659 662378 255665
rect 662326 255601 662378 255607
rect 662338 255559 662366 255601
rect 662324 255550 662380 255559
rect 662324 255485 662380 255494
rect 663970 229543 663998 397459
rect 664066 273351 664094 432017
rect 666658 318935 666686 504019
rect 666754 377247 666782 645211
rect 666850 631807 666878 786255
rect 666934 691297 666986 691303
rect 666934 691239 666986 691245
rect 666838 631801 666890 631807
rect 666838 631743 666890 631749
rect 666838 599093 666890 599099
rect 666838 599035 666890 599041
rect 666850 409363 666878 599035
rect 666946 541379 666974 691239
rect 667042 677539 667070 820813
rect 667030 677533 667082 677539
rect 667030 677475 667082 677481
rect 669538 613455 669566 954679
rect 672886 943193 672938 943199
rect 672886 943135 672938 943141
rect 672310 942601 672362 942607
rect 672310 942543 672362 942549
rect 669718 832415 669770 832421
rect 669718 832357 669770 832363
rect 669622 686265 669674 686271
rect 669622 686207 669674 686213
rect 669526 613449 669578 613455
rect 669526 613391 669578 613397
rect 666934 541373 666986 541379
rect 666934 541315 666986 541321
rect 666934 480989 666986 480995
rect 666934 480931 666986 480937
rect 666838 409357 666890 409363
rect 666838 409299 666890 409305
rect 666742 377241 666794 377247
rect 666742 377183 666794 377189
rect 666742 339871 666794 339877
rect 666742 339813 666794 339819
rect 666646 318929 666698 318935
rect 666646 318871 666698 318877
rect 665204 273606 665260 273615
rect 665204 273541 665260 273550
rect 665218 273425 665246 273541
rect 665206 273419 665258 273425
rect 665206 273361 665258 273367
rect 664054 273345 664106 273351
rect 664054 273287 664106 273293
rect 663958 229537 664010 229543
rect 663958 229479 664010 229485
rect 661174 183953 661226 183959
rect 661174 183895 661226 183901
rect 666754 182923 666782 339813
rect 666946 318343 666974 480931
rect 669634 423349 669662 686207
rect 669730 676503 669758 832357
rect 672214 783501 672266 783507
rect 672214 783443 672266 783449
rect 672022 779357 672074 779363
rect 672022 779299 672074 779305
rect 669814 774769 669866 774775
rect 669814 774711 669866 774717
rect 669718 676497 669770 676503
rect 669718 676439 669770 676445
rect 669718 645195 669770 645201
rect 669718 645137 669770 645143
rect 669730 497349 669758 645137
rect 669826 632547 669854 774711
rect 670966 763225 671018 763231
rect 670966 763167 671018 763173
rect 670978 717129 671006 763167
rect 671926 719047 671978 719053
rect 671926 718989 671978 718995
rect 670966 717123 671018 717129
rect 670966 717065 671018 717071
rect 670966 699955 671018 699961
rect 670966 699897 671018 699903
rect 670978 673173 671006 699897
rect 671938 674875 671966 718989
rect 672034 709063 672062 779299
rect 672118 778617 672170 778623
rect 672118 778559 672170 778565
rect 672022 709057 672074 709063
rect 672022 708999 672074 709005
rect 672130 706843 672158 778559
rect 672226 710543 672254 783443
rect 672322 765303 672350 942543
rect 672898 941867 672926 943135
rect 673844 941974 673900 941983
rect 673844 941909 673900 941918
rect 673858 941867 673886 941909
rect 672886 941861 672938 941867
rect 672886 941803 672938 941809
rect 673846 941861 673898 941867
rect 673846 941803 673898 941809
rect 672502 782317 672554 782323
rect 672502 782259 672554 782265
rect 672406 777655 672458 777661
rect 672406 777597 672458 777603
rect 672310 765297 672362 765303
rect 672310 765239 672362 765245
rect 672310 733625 672362 733631
rect 672310 733567 672362 733573
rect 672214 710537 672266 710543
rect 672214 710479 672266 710485
rect 672118 706837 672170 706843
rect 672118 706779 672170 706785
rect 672214 692925 672266 692931
rect 672214 692867 672266 692873
rect 672118 688633 672170 688639
rect 672118 688575 672170 688581
rect 671926 674869 671978 674875
rect 671926 674811 671978 674817
rect 670966 673167 671018 673173
rect 670966 673109 671018 673115
rect 671926 648303 671978 648309
rect 671926 648245 671978 648251
rect 671638 644603 671690 644609
rect 671638 644545 671690 644551
rect 671446 642309 671498 642315
rect 671446 642251 671498 642257
rect 670870 633651 670922 633657
rect 670870 633593 670922 633599
rect 669814 632541 669866 632547
rect 669814 632483 669866 632489
rect 670882 627483 670910 633593
rect 670966 630765 671018 630771
rect 670966 630707 671018 630713
rect 670978 628371 671006 630707
rect 670964 628362 671020 628371
rect 670964 628297 671020 628306
rect 670868 627474 670924 627483
rect 670868 627409 670924 627418
rect 669910 622107 669962 622113
rect 669910 622049 669962 622055
rect 669814 527091 669866 527097
rect 669814 527033 669866 527039
rect 669718 497343 669770 497349
rect 669718 497285 669770 497291
rect 669718 446431 669770 446437
rect 669718 446373 669770 446379
rect 669622 423343 669674 423349
rect 669622 423285 669674 423291
rect 669526 408987 669578 408993
rect 669526 408929 669578 408935
rect 666934 318337 666986 318343
rect 666934 318279 666986 318285
rect 669538 228951 669566 408929
rect 669622 385973 669674 385979
rect 669622 385915 669674 385921
rect 669526 228945 669578 228951
rect 669526 228887 669578 228893
rect 669634 227915 669662 385915
rect 669730 274979 669758 446373
rect 669826 363335 669854 527033
rect 669922 496535 669950 622049
rect 670882 590367 670910 627409
rect 670870 590361 670922 590367
rect 670870 590303 670922 590309
rect 670978 583411 671006 628297
rect 671350 599833 671402 599839
rect 671350 599775 671402 599781
rect 670966 583405 671018 583411
rect 670966 583347 671018 583353
rect 671362 526875 671390 599775
rect 671458 574531 671486 642251
rect 671542 599315 671594 599321
rect 671542 599257 671594 599263
rect 671446 574525 671498 574531
rect 671446 574467 671498 574473
rect 671554 529835 671582 599257
rect 671650 572015 671678 644545
rect 671734 627879 671786 627885
rect 671734 627821 671786 627827
rect 671746 584891 671774 627821
rect 671830 602053 671882 602059
rect 671830 601995 671882 602001
rect 671734 584885 671786 584891
rect 671734 584827 671786 584833
rect 671638 572009 671690 572015
rect 671638 571951 671690 571957
rect 671842 530871 671870 601995
rect 671938 575419 671966 648245
rect 672130 617895 672158 688575
rect 672226 619227 672254 692867
rect 672322 661703 672350 733567
rect 672418 709951 672446 777597
rect 672514 737701 672542 782259
rect 672694 779801 672746 779807
rect 672694 779743 672746 779749
rect 672598 764039 672650 764045
rect 672598 763981 672650 763987
rect 672502 737695 672554 737701
rect 672502 737637 672554 737643
rect 672406 709945 672458 709951
rect 672406 709887 672458 709893
rect 672514 702699 672542 737637
rect 672610 720311 672638 763981
rect 672598 720305 672650 720311
rect 672598 720247 672650 720253
rect 672598 717197 672650 717203
rect 672598 717139 672650 717145
rect 672502 702693 672554 702699
rect 672502 702635 672554 702641
rect 672406 692481 672458 692487
rect 672406 692423 672458 692429
rect 672310 661697 672362 661703
rect 672310 661639 672362 661645
rect 672418 650973 672446 692423
rect 672502 673167 672554 673173
rect 672502 673109 672554 673115
rect 672406 650967 672458 650973
rect 672406 650909 672458 650915
rect 672310 644085 672362 644091
rect 672310 644027 672362 644033
rect 672214 619221 672266 619227
rect 672214 619163 672266 619169
rect 672118 617889 672170 617895
rect 672118 617831 672170 617837
rect 672214 603681 672266 603687
rect 672214 603623 672266 603629
rect 672022 602719 672074 602725
rect 672022 602661 672074 602667
rect 671926 575413 671978 575419
rect 671926 575355 671978 575361
rect 671830 530865 671882 530871
rect 671830 530807 671882 530813
rect 671542 529829 671594 529835
rect 671542 529771 671594 529777
rect 672034 529243 672062 602661
rect 672118 601979 672170 601985
rect 672118 601921 672170 601927
rect 672130 532795 672158 601921
rect 672226 564467 672254 603623
rect 672322 573643 672350 644027
rect 672514 630771 672542 673109
rect 672610 671027 672638 717139
rect 672706 707435 672734 779743
rect 672898 763231 672926 941803
rect 673954 937247 673982 958971
rect 675394 958443 675422 958744
rect 675094 958437 675146 958443
rect 675094 958379 675146 958385
rect 675382 958437 675434 958443
rect 675382 958379 675434 958385
rect 674038 953923 674090 953929
rect 674038 953865 674090 953871
rect 674050 939615 674078 953865
rect 675106 953527 675134 958379
rect 675778 957671 675806 958078
rect 675764 957662 675820 957671
rect 675764 957597 675820 957606
rect 675490 957037 675518 957412
rect 675190 957031 675242 957037
rect 675190 956973 675242 956979
rect 675478 957031 675530 957037
rect 675478 956973 675530 956979
rect 675092 953518 675148 953527
rect 675092 953453 675148 953462
rect 675202 953379 675230 956973
rect 675490 956043 675518 956228
rect 675476 956034 675532 956043
rect 675476 955969 675532 955978
rect 675394 954743 675422 955044
rect 675382 954737 675434 954743
rect 675382 954679 675434 954685
rect 675490 953929 675518 954378
rect 675478 953923 675530 953929
rect 675478 953865 675530 953871
rect 675188 953370 675244 953379
rect 675188 953305 675244 953314
rect 675490 952079 675518 952528
rect 674134 952073 674186 952079
rect 674134 952015 674186 952021
rect 675478 952073 675530 952079
rect 675478 952015 675530 952021
rect 674036 939606 674092 939615
rect 674036 939541 674092 939550
rect 673940 937238 673996 937247
rect 673940 937173 673996 937182
rect 674146 936359 674174 952015
rect 674708 945378 674764 945387
rect 674708 945313 674764 945322
rect 674722 944901 674750 945313
rect 674710 944895 674762 944901
rect 674710 944837 674762 944843
rect 674708 944786 674764 944795
rect 674708 944721 674764 944730
rect 674722 944679 674750 944721
rect 674710 944673 674762 944679
rect 674710 944615 674762 944621
rect 674708 943750 674764 943759
rect 674708 943685 674764 943694
rect 674612 943158 674668 943167
rect 674612 943093 674668 943102
rect 674420 942640 674476 942649
rect 674420 942575 674422 942584
rect 674474 942575 674476 942584
rect 674422 942543 674474 942549
rect 674626 941941 674654 943093
rect 674722 942089 674750 943685
rect 674710 942083 674762 942089
rect 674710 942025 674762 942031
rect 674614 941935 674666 941941
rect 674614 941877 674666 941883
rect 674900 940642 674956 940651
rect 674900 940577 674956 940586
rect 674914 939129 674942 940577
rect 674902 939123 674954 939129
rect 674902 939065 674954 939071
rect 674132 936350 674188 936359
rect 674132 936285 674188 936294
rect 679796 928654 679852 928663
rect 679796 928589 679852 928598
rect 679810 928071 679838 928589
rect 679796 928062 679852 928071
rect 679796 927997 679852 928006
rect 679810 927437 679838 927997
rect 679798 927431 679850 927437
rect 679798 927373 679850 927379
rect 675106 877509 675408 877537
rect 675106 876419 675134 877509
rect 675778 876419 675806 876900
rect 675092 876410 675148 876419
rect 675092 876345 675148 876354
rect 675764 876410 675820 876419
rect 675764 876345 675820 876354
rect 675092 876262 675148 876271
rect 675148 876220 675408 876248
rect 675092 876197 675148 876206
rect 675284 875818 675340 875827
rect 675284 875753 675340 875762
rect 674230 872153 674282 872159
rect 674230 872095 674282 872101
rect 673654 867861 673706 867867
rect 673654 867803 673706 867809
rect 672886 763225 672938 763231
rect 672886 763167 672938 763173
rect 672886 762559 672938 762565
rect 672886 762501 672938 762507
rect 672898 717869 672926 762501
rect 673666 751655 673694 867803
rect 674242 780515 674270 872095
rect 674902 871931 674954 871937
rect 674902 871873 674954 871879
rect 674326 868379 674378 868385
rect 674326 868321 674378 868327
rect 674228 780506 674284 780515
rect 674228 780441 674284 780450
rect 674230 773659 674282 773665
rect 674230 773601 674282 773607
rect 673652 751646 673708 751655
rect 673652 751581 673708 751590
rect 674038 750275 674090 750281
rect 674038 750217 674090 750223
rect 674050 720089 674078 750217
rect 674134 735697 674186 735703
rect 674134 735639 674186 735645
rect 674038 720083 674090 720089
rect 674038 720025 674090 720031
rect 672886 717863 672938 717869
rect 672886 717805 672938 717811
rect 672898 717203 672926 717805
rect 672886 717197 672938 717203
rect 672886 717139 672938 717145
rect 672694 707429 672746 707435
rect 672694 707371 672746 707377
rect 672694 674055 672746 674061
rect 672694 673997 672746 674003
rect 672598 671021 672650 671027
rect 672598 670963 672650 670969
rect 672598 643419 672650 643425
rect 672598 643361 672650 643367
rect 672502 630765 672554 630771
rect 672502 630707 672554 630713
rect 672502 597169 672554 597175
rect 672502 597111 672554 597117
rect 672406 583627 672458 583633
rect 672406 583569 672458 583575
rect 672418 578897 672446 583569
rect 672406 578891 672458 578897
rect 672406 578833 672458 578839
rect 672310 573637 672362 573643
rect 672310 573579 672362 573585
rect 672214 564461 672266 564467
rect 672214 564403 672266 564409
rect 672214 558763 672266 558769
rect 672214 558705 672266 558711
rect 672226 539899 672254 558705
rect 672214 539893 672266 539899
rect 672214 539835 672266 539841
rect 672118 532789 672170 532795
rect 672118 532731 672170 532737
rect 672514 529909 672542 597111
rect 672610 571423 672638 643361
rect 672706 630549 672734 673997
rect 674146 668627 674174 735639
rect 674242 713027 674270 773601
rect 674338 772671 674366 868321
rect 674914 866905 674942 871873
rect 675298 871364 675326 875753
rect 675490 874051 675518 874384
rect 675476 874042 675532 874051
rect 675476 873977 675532 873986
rect 675394 873459 675422 873866
rect 675380 873450 675436 873459
rect 675380 873385 675436 873394
rect 675394 872867 675422 873200
rect 675380 872858 675436 872867
rect 675380 872793 675436 872802
rect 675490 872159 675518 872534
rect 675572 872414 675628 872423
rect 675572 872349 675628 872358
rect 675478 872153 675530 872159
rect 675478 872095 675530 872101
rect 675586 871937 675614 872349
rect 675574 871931 675626 871937
rect 675574 871873 675626 871879
rect 675298 871336 675408 871364
rect 674998 869045 675050 869051
rect 674998 868987 675050 868993
rect 674902 866899 674954 866905
rect 674902 866841 674954 866847
rect 674806 846771 674858 846777
rect 674806 846713 674858 846719
rect 674818 832292 674846 846713
rect 674722 832264 674846 832292
rect 674722 826575 674750 832264
rect 674422 826569 674474 826575
rect 674422 826511 674474 826517
rect 674710 826569 674762 826575
rect 674710 826511 674762 826517
rect 674434 806447 674462 826511
rect 674422 806441 674474 806447
rect 674422 806383 674474 806389
rect 674614 806441 674666 806447
rect 674614 806383 674666 806389
rect 674518 784981 674570 784987
rect 674518 784923 674570 784929
rect 674422 780467 674474 780473
rect 674422 780409 674474 780415
rect 674324 772662 674380 772671
rect 674324 772597 674380 772606
rect 674326 765889 674378 765895
rect 674324 765854 674326 765863
rect 674378 765854 674380 765863
rect 674324 765789 674380 765798
rect 674434 750281 674462 780409
rect 674422 750275 674474 750281
rect 674422 750217 674474 750223
rect 674530 740088 674558 784923
rect 674626 782323 674654 806383
rect 675010 783156 675038 868987
rect 675094 866899 675146 866905
rect 675094 866841 675146 866847
rect 675106 846777 675134 866841
rect 675298 862965 675326 871336
rect 675394 869907 675422 870092
rect 675380 869898 675436 869907
rect 675380 869833 675436 869842
rect 675490 869051 675518 869500
rect 675478 869045 675530 869051
rect 675478 868987 675530 868993
rect 675394 868385 675422 868875
rect 675382 868379 675434 868385
rect 675382 868321 675434 868327
rect 675394 867867 675422 868242
rect 675382 867861 675434 867867
rect 675382 867803 675434 867809
rect 675394 866947 675422 867058
rect 675380 866938 675436 866947
rect 675380 866873 675436 866882
rect 675394 865351 675422 865839
rect 675382 865345 675434 865351
rect 675382 865287 675434 865293
rect 675490 864727 675518 865208
rect 675476 864718 675532 864727
rect 675476 864653 675532 864662
rect 675382 862977 675434 862983
rect 675298 862937 675382 862965
rect 675682 862951 675710 863358
rect 675382 862919 675434 862925
rect 675668 862942 675724 862951
rect 675668 862877 675724 862886
rect 675382 862607 675434 862613
rect 675382 862549 675434 862555
rect 675394 846777 675422 862549
rect 675094 846771 675146 846777
rect 675094 846713 675146 846719
rect 675382 846771 675434 846777
rect 675382 846713 675434 846719
rect 675574 846771 675626 846777
rect 675574 846713 675626 846719
rect 675586 832292 675614 846713
rect 675490 832264 675614 832292
rect 675490 826575 675518 832264
rect 675478 826569 675530 826575
rect 675478 826511 675530 826517
rect 675670 826569 675722 826575
rect 675670 826511 675722 826517
rect 675682 806447 675710 826511
rect 675286 806441 675338 806447
rect 675286 806383 675338 806389
rect 675670 806441 675722 806447
rect 675670 806383 675722 806389
rect 674818 783128 675038 783156
rect 674614 782317 674666 782323
rect 674614 782259 674666 782265
rect 674818 777407 674846 783128
rect 674998 783057 675050 783063
rect 674998 782999 675050 783005
rect 675010 777555 675038 782999
rect 675298 782120 675326 806383
rect 675778 787915 675806 788322
rect 675764 787906 675820 787915
rect 675764 787841 675820 787850
rect 675490 787471 675518 787656
rect 675476 787462 675532 787471
rect 675476 787397 675532 787406
rect 675778 786731 675806 787035
rect 675764 786722 675820 786731
rect 675764 786657 675820 786666
rect 675394 784987 675422 785214
rect 675382 784981 675434 784987
rect 675382 784923 675434 784929
rect 675778 784215 675806 784622
rect 675764 784206 675820 784215
rect 675764 784141 675820 784150
rect 675394 783507 675422 783999
rect 675382 783501 675434 783507
rect 675382 783443 675434 783449
rect 675394 783063 675422 783364
rect 675382 783057 675434 783063
rect 675382 782999 675434 783005
rect 675394 782323 675422 782803
rect 675382 782317 675434 782323
rect 675382 782259 675434 782265
rect 675408 782180 675792 782194
rect 675394 782166 675806 782180
rect 675394 782120 675422 782166
rect 675298 782092 675422 782120
rect 675778 781995 675806 782166
rect 675764 781986 675820 781995
rect 675764 781921 675820 781930
rect 675094 780541 675146 780547
rect 675094 780483 675146 780489
rect 674996 777546 675052 777555
rect 674996 777481 675052 777490
rect 674804 777398 674860 777407
rect 674804 777333 674860 777342
rect 675106 777069 675134 780483
rect 675490 780473 675518 780848
rect 675478 780467 675530 780473
rect 675478 780409 675530 780415
rect 675394 779807 675422 780330
rect 675382 779801 675434 779807
rect 675382 779743 675434 779749
rect 675490 779363 675518 779664
rect 675478 779357 675530 779363
rect 675478 779299 675530 779305
rect 675394 778623 675422 779031
rect 675382 778617 675434 778623
rect 675382 778559 675434 778565
rect 675490 777661 675518 777814
rect 675478 777655 675530 777661
rect 675478 777597 675530 777603
rect 675094 777063 675146 777069
rect 675094 777005 675146 777011
rect 675382 777063 675434 777069
rect 675382 777005 675434 777011
rect 675394 776630 675422 777005
rect 675394 775515 675422 775995
rect 674806 775509 674858 775515
rect 674806 775451 674858 775457
rect 675382 775509 675434 775515
rect 675382 775451 675434 775457
rect 674710 767813 674762 767819
rect 674708 767778 674710 767787
rect 674762 767778 674764 767787
rect 674708 767713 674764 767722
rect 674710 766925 674762 766931
rect 674708 766890 674710 766899
rect 674762 766890 674764 766899
rect 674708 766825 674764 766834
rect 674710 765297 674762 765303
rect 674708 765262 674710 765271
rect 674762 765262 674764 765271
rect 674708 765197 674764 765206
rect 674708 764078 674764 764087
rect 674708 764013 674710 764022
rect 674762 764013 674764 764022
rect 674710 763981 674762 763987
rect 674708 763338 674764 763347
rect 674708 763273 674764 763282
rect 674722 763231 674750 763273
rect 674710 763225 674762 763231
rect 674710 763167 674762 763173
rect 674708 762598 674764 762607
rect 674708 762533 674710 762542
rect 674762 762533 674764 762542
rect 674710 762501 674762 762507
rect 674434 740060 674558 740088
rect 674326 722525 674378 722531
rect 674324 722490 674326 722499
rect 674378 722490 674380 722499
rect 674324 722425 674380 722434
rect 674326 720897 674378 720903
rect 674324 720862 674326 720871
rect 674378 720862 674380 720871
rect 674324 720797 674380 720806
rect 674326 720083 674378 720089
rect 674326 720025 674378 720031
rect 674338 713767 674366 720025
rect 674434 714507 674462 740060
rect 674710 730517 674762 730523
rect 674710 730459 674762 730465
rect 674614 728667 674666 728673
rect 674614 728609 674666 728615
rect 674516 717902 674572 717911
rect 674516 717837 674518 717846
rect 674570 717837 674572 717846
rect 674518 717805 674570 717811
rect 674420 714498 674476 714507
rect 674420 714433 674476 714442
rect 674324 713758 674380 713767
rect 674324 713693 674380 713702
rect 674228 713018 674284 713027
rect 674228 712953 674284 712962
rect 674422 710537 674474 710543
rect 674420 710502 674422 710511
rect 674474 710502 674476 710511
rect 674420 710437 674476 710446
rect 674422 709057 674474 709063
rect 674420 709022 674422 709031
rect 674474 709022 674476 709031
rect 674420 708957 674476 708966
rect 674422 707429 674474 707435
rect 674420 707394 674422 707403
rect 674474 707394 674476 707403
rect 674420 707329 674476 707338
rect 674326 690705 674378 690711
rect 674326 690647 674378 690653
rect 674230 687375 674282 687381
rect 674230 687317 674282 687323
rect 674132 668618 674188 668627
rect 674132 668553 674188 668562
rect 672886 648081 672938 648087
rect 672886 648023 672938 648029
rect 672694 630543 672746 630549
rect 672694 630485 672746 630491
rect 672694 598427 672746 598433
rect 672694 598369 672746 598375
rect 672598 571417 672650 571423
rect 672598 571359 672650 571365
rect 672502 529903 672554 529909
rect 672502 529845 672554 529851
rect 672022 529237 672074 529243
rect 672022 529179 672074 529185
rect 672706 526949 672734 598369
rect 672790 578891 672842 578897
rect 672790 578833 672842 578839
rect 672802 558769 672830 578833
rect 672898 573051 672926 648023
rect 674132 630730 674188 630739
rect 674132 630665 674188 630674
rect 674146 630623 674174 630665
rect 674134 630617 674186 630623
rect 674134 630559 674186 630565
rect 673846 630543 673898 630549
rect 673846 630485 673898 630491
rect 673858 629851 673886 630485
rect 673844 629842 673900 629851
rect 673844 629777 673900 629786
rect 673844 629102 673900 629111
rect 673844 629037 673900 629046
rect 673858 627885 673886 629037
rect 673846 627879 673898 627885
rect 673846 627821 673898 627827
rect 674036 624958 674092 624967
rect 674036 624893 674092 624902
rect 673846 619221 673898 619227
rect 673846 619163 673898 619169
rect 673858 618011 673886 619163
rect 673844 618002 673900 618011
rect 673844 617937 673900 617946
rect 673846 617889 673898 617895
rect 673846 617831 673898 617837
rect 673858 616383 673886 617831
rect 673844 616374 673900 616383
rect 673844 616309 673900 616318
rect 674050 604839 674078 624893
rect 674242 619491 674270 687317
rect 674338 623635 674366 690647
rect 674518 685525 674570 685531
rect 674518 685467 674570 685473
rect 674422 676497 674474 676503
rect 674420 676462 674422 676471
rect 674474 676462 674476 676471
rect 674420 676397 674476 676406
rect 674422 674869 674474 674875
rect 674420 674834 674422 674843
rect 674474 674834 674476 674843
rect 674420 674769 674476 674778
rect 674420 674094 674476 674103
rect 674420 674029 674422 674038
rect 674474 674029 674476 674038
rect 674422 673997 674474 674003
rect 674422 669615 674474 669621
rect 674422 669557 674474 669563
rect 674324 623626 674380 623635
rect 674324 623561 674380 623570
rect 674434 622747 674462 669557
rect 674530 626151 674558 685467
rect 674626 668035 674654 728609
rect 674722 671143 674750 730459
rect 674818 726379 674846 775451
rect 675394 773665 675422 774155
rect 675382 773659 675434 773665
rect 675382 773601 675434 773607
rect 679796 750166 679852 750175
rect 679796 750101 679852 750110
rect 679810 749583 679838 750101
rect 679796 749574 679852 749583
rect 679796 749509 679852 749518
rect 679810 748875 679838 749509
rect 679798 748869 679850 748875
rect 679798 748811 679850 748817
rect 675092 743358 675148 743367
rect 675148 743316 675408 743344
rect 675092 743293 675148 743302
rect 675298 742724 675422 742752
rect 675298 742678 675326 742724
rect 675106 742650 675326 742678
rect 675394 742664 675422 742724
rect 675106 741443 675134 742650
rect 675778 741739 675806 742035
rect 675764 741730 675820 741739
rect 675764 741665 675820 741674
rect 675092 741434 675148 741443
rect 675092 741369 675148 741378
rect 675476 740398 675532 740407
rect 675476 740333 675532 740342
rect 675490 740222 675518 740333
rect 675490 739371 675518 739630
rect 675476 739362 675532 739371
rect 675476 739297 675532 739306
rect 675394 738631 675422 738999
rect 675380 738622 675436 738631
rect 675380 738557 675436 738566
rect 675394 737923 675422 738372
rect 674902 737917 674954 737923
rect 674902 737859 674954 737865
rect 675382 737917 675434 737923
rect 675382 737859 675434 737865
rect 674806 726373 674858 726379
rect 674806 726315 674858 726321
rect 674806 721933 674858 721939
rect 674804 721898 674806 721907
rect 674858 721898 674860 721907
rect 674804 721833 674860 721842
rect 674806 720305 674858 720311
rect 674804 720270 674806 720279
rect 674858 720270 674860 720279
rect 674804 720205 674860 720214
rect 674804 719086 674860 719095
rect 674804 719021 674806 719030
rect 674858 719021 674860 719030
rect 674806 718989 674858 718995
rect 674806 709945 674858 709951
rect 674804 709910 674806 709919
rect 674858 709910 674860 709919
rect 674804 709845 674860 709854
rect 674806 706837 674858 706843
rect 674804 706802 674806 706811
rect 674858 706802 674860 706811
rect 674804 706737 674860 706746
rect 674806 702693 674858 702699
rect 674806 702635 674858 702641
rect 674818 692487 674846 702635
rect 674806 692481 674858 692487
rect 674806 692423 674858 692429
rect 674804 689338 674860 689347
rect 674804 689273 674860 689282
rect 674818 679727 674846 689273
rect 674914 688311 674942 737859
rect 675490 737701 675518 737780
rect 675478 737695 675530 737701
rect 675478 737637 675530 737643
rect 675094 737399 675146 737405
rect 675094 737341 675146 737347
rect 675106 732077 675134 737341
rect 675778 736707 675806 737159
rect 675764 736698 675820 736707
rect 675764 736633 675820 736642
rect 675490 735703 675518 735856
rect 675478 735697 675530 735703
rect 675478 735639 675530 735645
rect 675394 734963 675422 735338
rect 675190 734957 675242 734963
rect 675190 734899 675242 734905
rect 675382 734957 675434 734963
rect 675382 734899 675434 734905
rect 675202 732563 675230 734899
rect 675682 734487 675710 734672
rect 675668 734478 675724 734487
rect 675668 734413 675724 734422
rect 675490 733631 675518 734006
rect 675478 733625 675530 733631
rect 675478 733567 675530 733573
rect 675188 732554 675244 732563
rect 675188 732489 675244 732498
rect 675490 732373 675518 732822
rect 675190 732367 675242 732373
rect 675190 732309 675242 732315
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 675094 732071 675146 732077
rect 675094 732013 675146 732019
rect 675202 726472 675230 732309
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 675490 730523 675518 730972
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 675490 728673 675518 729155
rect 675478 728667 675530 728673
rect 675478 728609 675530 728615
rect 675010 726444 675230 726472
rect 674900 688302 674956 688311
rect 674900 688237 674956 688246
rect 674902 683675 674954 683681
rect 674902 683617 674954 683623
rect 674804 679718 674860 679727
rect 674804 679653 674860 679662
rect 674806 677533 674858 677539
rect 674804 677498 674806 677507
rect 674858 677498 674860 677507
rect 674804 677433 674860 677442
rect 674806 675905 674858 675911
rect 674804 675870 674806 675879
rect 674858 675870 674860 675879
rect 674804 675805 674860 675814
rect 674804 673206 674860 673215
rect 674804 673141 674806 673150
rect 674858 673141 674860 673150
rect 674806 673109 674858 673115
rect 674708 671134 674764 671143
rect 674708 671069 674764 671078
rect 674914 669621 674942 683617
rect 674902 669615 674954 669621
rect 674902 669557 674954 669563
rect 674612 668026 674668 668035
rect 674612 667961 674668 667970
rect 675010 664779 675038 726444
rect 675094 726373 675146 726379
rect 675094 726315 675146 726321
rect 675106 716283 675134 726315
rect 679700 718050 679756 718059
rect 679700 717985 679756 717994
rect 679714 717129 679742 717985
rect 679702 717123 679754 717129
rect 679702 717065 679754 717071
rect 675092 716274 675148 716283
rect 675092 716209 675148 716218
rect 679714 699961 679742 717065
rect 679796 705174 679852 705183
rect 679796 705109 679852 705118
rect 679810 704591 679838 705109
rect 679796 704582 679852 704591
rect 679796 704517 679852 704526
rect 679810 702773 679838 704517
rect 679798 702767 679850 702773
rect 679798 702709 679850 702715
rect 679702 699955 679754 699961
rect 679702 699897 679754 699903
rect 675394 697931 675422 698338
rect 675380 697922 675436 697931
rect 675380 697857 675436 697866
rect 675490 697339 675518 697672
rect 675476 697330 675532 697339
rect 675476 697265 675532 697274
rect 675394 696895 675422 697035
rect 675380 696886 675436 696895
rect 675380 696821 675436 696830
rect 675778 694823 675806 695195
rect 675764 694814 675820 694823
rect 675764 694749 675820 694758
rect 675284 694666 675340 694675
rect 675340 694624 675408 694652
rect 675284 694601 675340 694610
rect 675778 693491 675806 693972
rect 675764 693482 675820 693491
rect 675764 693417 675820 693426
rect 675394 692931 675422 693380
rect 675382 692925 675434 692931
rect 675382 692867 675434 692873
rect 675490 692487 675518 692788
rect 675478 692481 675530 692487
rect 675478 692423 675530 692429
rect 675778 691715 675806 692159
rect 675764 691706 675820 691715
rect 675764 691641 675820 691650
rect 675490 690711 675518 690864
rect 675478 690705 675530 690711
rect 675478 690647 675530 690653
rect 675394 689823 675422 690346
rect 675094 689817 675146 689823
rect 675094 689759 675146 689765
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 675106 685647 675134 689759
rect 675778 689199 675806 689680
rect 675764 689190 675820 689199
rect 675764 689125 675820 689134
rect 675490 688639 675518 689014
rect 675478 688633 675530 688639
rect 675478 688575 675530 688581
rect 675490 687381 675518 687830
rect 675478 687375 675530 687381
rect 675478 687317 675530 687323
rect 675394 686271 675422 686646
rect 675382 686265 675434 686271
rect 675382 686207 675434 686213
rect 675092 685638 675148 685647
rect 675092 685573 675148 685582
rect 675490 685531 675518 685980
rect 675478 685525 675530 685531
rect 675478 685467 675530 685473
rect 675490 683681 675518 684130
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 675092 672318 675148 672327
rect 675092 672253 675148 672262
rect 675106 671027 675134 672253
rect 675094 671021 675146 671027
rect 675094 670963 675146 670969
rect 674996 664770 675052 664779
rect 674996 664705 675052 664714
rect 674710 661697 674762 661703
rect 674708 661662 674710 661671
rect 674762 661662 674764 661671
rect 674708 661597 674764 661606
rect 674996 652782 675052 652791
rect 674996 652717 675052 652726
rect 674806 650967 674858 650973
rect 674806 650909 674858 650915
rect 674614 650893 674666 650899
rect 674614 650835 674666 650841
rect 674626 646459 674654 650835
rect 674818 647643 674846 650909
rect 675010 650899 675038 652717
rect 674998 650893 675050 650899
rect 674998 650835 675050 650841
rect 675106 647736 675134 670963
rect 679796 660034 679852 660043
rect 679796 659969 679852 659978
rect 679810 659303 679838 659969
rect 679796 659294 679852 659303
rect 679796 659229 679852 659238
rect 679810 656745 679838 659229
rect 679798 656739 679850 656745
rect 679798 656681 679850 656687
rect 675490 652643 675518 653124
rect 675476 652634 675532 652643
rect 675476 652569 675532 652578
rect 675490 652199 675518 652458
rect 675476 652190 675532 652199
rect 675476 652125 675532 652134
rect 675298 651821 675408 651849
rect 675298 651015 675326 651821
rect 675284 651006 675340 651015
rect 675284 650941 675340 650950
rect 675778 649683 675806 650016
rect 675764 649674 675820 649683
rect 675764 649609 675820 649618
rect 675298 649484 675422 649512
rect 675298 649438 675326 649484
rect 675202 649410 675326 649438
rect 675394 649424 675422 649484
rect 675202 648351 675230 649410
rect 675298 648785 675408 648813
rect 675188 648342 675244 648351
rect 675298 648309 675326 648785
rect 675188 648277 675244 648286
rect 675286 648303 675338 648309
rect 675286 648245 675338 648251
rect 675202 648152 675408 648180
rect 675202 648087 675230 648152
rect 675190 648081 675242 648087
rect 675190 648023 675242 648029
rect 675010 647708 675134 647736
rect 674806 647637 674858 647643
rect 674806 647579 674858 647585
rect 674614 646453 674666 646459
rect 674614 646395 674666 646401
rect 674516 626142 674572 626151
rect 674516 626077 674572 626086
rect 674420 622738 674476 622747
rect 674420 622673 674476 622682
rect 674228 619482 674284 619491
rect 674228 619417 674284 619426
rect 674036 604830 674092 604839
rect 674036 604765 674092 604774
rect 674626 603687 674654 646395
rect 674806 645121 674858 645127
rect 674806 645063 674858 645069
rect 674710 632541 674762 632547
rect 674708 632506 674710 632515
rect 674762 632506 674764 632515
rect 674708 632441 674764 632450
rect 674710 631801 674762 631807
rect 674708 631766 674710 631775
rect 674762 631766 674764 631775
rect 674708 631701 674764 631710
rect 674818 630864 674846 645063
rect 674900 641978 674956 641987
rect 674900 641913 674956 641922
rect 674722 630836 674846 630864
rect 674722 627164 674750 630836
rect 674722 627136 674846 627164
rect 674614 603681 674666 603687
rect 674614 603623 674666 603629
rect 674818 602873 674846 627136
rect 674914 625707 674942 641913
rect 675010 633657 675038 647708
rect 675094 647637 675146 647643
rect 675146 647589 675408 647617
rect 675094 647579 675146 647585
rect 675106 645127 675134 647579
rect 675394 646459 675422 646982
rect 675382 646453 675434 646459
rect 675382 646395 675434 646401
rect 675490 645539 675518 645650
rect 675476 645530 675532 645539
rect 675476 645465 675532 645474
rect 675190 645269 675242 645275
rect 675190 645211 675242 645217
rect 675094 645121 675146 645127
rect 675094 645063 675146 645069
rect 675202 641871 675230 645211
rect 675490 644609 675518 645132
rect 675478 644603 675530 644609
rect 675478 644545 675530 644551
rect 675490 644091 675518 644466
rect 675478 644085 675530 644091
rect 675478 644027 675530 644033
rect 675394 643425 675422 643831
rect 675382 643419 675434 643425
rect 675382 643361 675434 643367
rect 675490 642315 675518 642616
rect 675478 642309 675530 642315
rect 675478 642251 675530 642257
rect 675190 641865 675242 641871
rect 675190 641807 675242 641813
rect 675382 641865 675434 641871
rect 675382 641807 675434 641813
rect 675394 641432 675422 641807
rect 675092 640498 675148 640507
rect 675092 640433 675148 640442
rect 674998 633651 675050 633657
rect 674998 633593 675050 633599
rect 674900 625698 674956 625707
rect 674900 625633 674956 625642
rect 675106 622155 675134 640433
rect 675778 640359 675806 640795
rect 675764 640350 675820 640359
rect 675764 640285 675820 640294
rect 675394 638583 675422 638955
rect 675380 638574 675436 638583
rect 675380 638509 675436 638518
rect 675188 637834 675244 637843
rect 675188 637769 675244 637778
rect 675202 630147 675230 637769
rect 676724 635022 676780 635031
rect 676724 634957 676780 634966
rect 676052 633246 676108 633255
rect 676052 633181 676108 633190
rect 675188 630138 675244 630147
rect 675188 630073 675244 630082
rect 676066 624819 676094 633181
rect 676738 630147 676766 634957
rect 676724 630138 676780 630147
rect 676724 630073 676780 630082
rect 676052 624810 676108 624819
rect 676052 624745 676108 624754
rect 675092 622146 675148 622155
rect 675092 622081 675148 622090
rect 679700 615042 679756 615051
rect 679700 614977 679756 614986
rect 679714 614459 679742 614977
rect 679700 614450 679756 614459
rect 679700 614385 679756 614394
rect 679714 613529 679742 614385
rect 679702 613523 679754 613529
rect 679702 613465 679754 613471
rect 675106 608118 675408 608146
rect 675106 607799 675134 608118
rect 675092 607790 675148 607799
rect 675092 607725 675148 607734
rect 675092 607494 675148 607503
rect 675148 607452 675408 607480
rect 675092 607429 675148 607438
rect 675682 606467 675710 606835
rect 675668 606458 675724 606467
rect 675668 606393 675724 606402
rect 675106 604987 675408 605009
rect 675092 604981 675408 604987
rect 675092 604978 675148 604981
rect 675092 604913 675148 604922
rect 675106 604418 675408 604446
rect 673750 602867 673802 602873
rect 673750 602809 673802 602815
rect 674806 602867 674858 602873
rect 674806 602809 674858 602815
rect 672886 573045 672938 573051
rect 672886 572987 672938 572993
rect 673762 561655 673790 602809
rect 675106 601985 675134 604418
rect 675202 603785 675408 603813
rect 675202 602059 675230 603785
rect 675286 603681 675338 603687
rect 675286 603623 675338 603629
rect 675190 602053 675242 602059
rect 675190 601995 675242 602001
rect 675094 601979 675146 601985
rect 675298 601973 675326 603623
rect 675394 602725 675422 603174
rect 675478 602867 675530 602873
rect 675478 602809 675530 602815
rect 675382 602719 675434 602725
rect 675382 602661 675434 602667
rect 675490 602582 675518 602809
rect 675298 601945 675408 601973
rect 675094 601921 675146 601927
rect 675190 601905 675242 601911
rect 675190 601847 675242 601853
rect 675202 596879 675230 601847
rect 675778 600251 675806 600658
rect 675764 600242 675820 600251
rect 675764 600177 675820 600186
rect 675394 599839 675422 600140
rect 675382 599833 675434 599839
rect 675382 599775 675434 599781
rect 675394 599321 675422 599474
rect 675382 599315 675434 599321
rect 675382 599257 675434 599263
rect 675490 598433 675518 598808
rect 675478 598427 675530 598433
rect 675478 598369 675530 598375
rect 675490 597175 675518 597624
rect 675478 597169 675530 597175
rect 675478 597111 675530 597117
rect 675190 596873 675242 596879
rect 675190 596815 675242 596821
rect 675382 596873 675434 596879
rect 675382 596815 675434 596821
rect 675394 596440 675422 596815
rect 675778 595367 675806 595774
rect 675764 595358 675820 595367
rect 675764 595293 675820 595302
rect 675778 593443 675806 593955
rect 675764 593434 675820 593443
rect 675764 593369 675820 593378
rect 679702 590361 679754 590367
rect 679702 590303 679754 590309
rect 674708 586478 674764 586487
rect 674708 586413 674764 586422
rect 674422 586365 674474 586371
rect 674420 586330 674422 586339
rect 674474 586330 674476 586339
rect 674420 586265 674476 586274
rect 674422 585477 674474 585483
rect 674420 585442 674422 585451
rect 674474 585442 674476 585451
rect 674420 585377 674476 585386
rect 674614 584885 674666 584891
rect 674612 584850 674614 584859
rect 674666 584850 674668 584859
rect 674722 584817 674750 586413
rect 674612 584785 674668 584794
rect 674710 584811 674762 584817
rect 674710 584753 674762 584759
rect 674228 584554 674284 584563
rect 674228 584489 674284 584498
rect 674242 575979 674270 584489
rect 674708 583666 674764 583675
rect 674708 583601 674710 583610
rect 674762 583601 674764 583610
rect 674710 583569 674762 583575
rect 674710 583405 674762 583411
rect 674708 583370 674710 583379
rect 674762 583370 674764 583379
rect 674708 583305 674764 583314
rect 679714 582935 679742 590303
rect 679990 583405 680042 583411
rect 679990 583347 680042 583353
rect 679700 582926 679756 582935
rect 679700 582861 679756 582870
rect 674228 575970 674284 575979
rect 674228 575905 674284 575914
rect 674710 575413 674762 575419
rect 674708 575378 674710 575387
rect 674762 575378 674764 575387
rect 674708 575313 674764 575322
rect 674710 574525 674762 574531
rect 674708 574490 674710 574499
rect 674762 574490 674764 574499
rect 674708 574425 674764 574434
rect 674422 573637 674474 573643
rect 674420 573602 674422 573611
rect 674474 573602 674476 573611
rect 674420 573537 674476 573546
rect 674710 573045 674762 573051
rect 674708 573010 674710 573019
rect 674762 573010 674764 573019
rect 674708 572945 674764 572954
rect 674422 572009 674474 572015
rect 674420 571974 674422 571983
rect 674474 571974 674476 571983
rect 674420 571909 674476 571918
rect 674710 571417 674762 571423
rect 674708 571382 674710 571391
rect 674762 571382 674764 571391
rect 674708 571317 674764 571326
rect 679796 569754 679852 569763
rect 679796 569689 679852 569698
rect 679810 569171 679838 569689
rect 679796 569162 679852 569171
rect 679796 569097 679852 569106
rect 679810 567427 679838 569097
rect 679798 567421 679850 567427
rect 680002 567395 680030 583347
rect 679798 567363 679850 567369
rect 679988 567386 680044 567395
rect 679988 567321 680044 567330
rect 674998 564461 675050 564467
rect 674998 564403 675050 564409
rect 673750 561649 673802 561655
rect 673750 561591 673802 561597
rect 674230 559577 674282 559583
rect 674230 559519 674282 559525
rect 672790 558763 672842 558769
rect 672790 558705 672842 558711
rect 674134 558097 674186 558103
rect 674134 558039 674186 558045
rect 674038 554545 674090 554551
rect 674038 554487 674090 554493
rect 673846 532789 673898 532795
rect 673846 532731 673898 532737
rect 673858 530987 673886 532731
rect 673844 530978 673900 530987
rect 673844 530913 673900 530922
rect 673846 530865 673898 530871
rect 673846 530807 673898 530813
rect 673858 530099 673886 530807
rect 673844 530090 673900 530099
rect 673844 530025 673900 530034
rect 673846 529903 673898 529909
rect 673846 529845 673898 529851
rect 673750 529829 673802 529835
rect 673750 529771 673802 529777
rect 673762 528619 673790 529771
rect 673858 529359 673886 529845
rect 673844 529350 673900 529359
rect 673844 529285 673900 529294
rect 673846 529237 673898 529243
rect 673846 529179 673898 529185
rect 673748 528610 673804 528619
rect 673748 528545 673804 528554
rect 673858 527879 673886 529179
rect 673844 527870 673900 527879
rect 673844 527805 673900 527814
rect 673748 526982 673804 526991
rect 672694 526943 672746 526949
rect 673748 526917 673804 526926
rect 673846 526943 673898 526949
rect 672694 526885 672746 526891
rect 673762 526875 673790 526917
rect 673846 526885 673898 526891
rect 671350 526869 671402 526875
rect 671350 526811 671402 526817
rect 673750 526869 673802 526875
rect 673750 526811 673802 526817
rect 673858 526251 673886 526885
rect 673844 526242 673900 526251
rect 673844 526177 673900 526186
rect 674050 498089 674078 554487
rect 674038 498083 674090 498089
rect 674038 498025 674090 498031
rect 674146 497960 674174 558039
rect 674050 497932 674174 497960
rect 674242 497941 674270 559519
rect 675010 556790 675038 564403
rect 675092 562946 675148 562955
rect 675148 562904 675408 562932
rect 675092 562881 675148 562890
rect 675298 562312 675422 562340
rect 675298 562266 675326 562312
rect 675106 562238 675326 562266
rect 675394 562252 675422 562312
rect 675106 561771 675134 562238
rect 675092 561762 675148 561771
rect 675092 561697 675148 561706
rect 675094 561649 675146 561655
rect 675094 561591 675146 561597
rect 675284 561614 675340 561623
rect 675106 557417 675134 561591
rect 675394 561600 675422 561660
rect 675340 561572 675422 561600
rect 675284 561549 675340 561558
rect 675394 559583 675422 559810
rect 675382 559577 675434 559583
rect 675382 559519 675434 559525
rect 675490 558959 675518 559218
rect 675476 558950 675532 558959
rect 675476 558885 675532 558894
rect 675394 558103 675422 558626
rect 675382 558097 675434 558103
rect 675382 558039 675434 558045
rect 675778 557775 675806 557960
rect 675764 557766 675820 557775
rect 675764 557701 675820 557710
rect 675106 557389 675408 557417
rect 675010 556762 675326 556790
rect 675298 556716 675326 556762
rect 675394 556716 675422 556776
rect 675298 556688 675422 556716
rect 675190 555877 675242 555883
rect 675190 555819 675242 555825
rect 674326 555063 674378 555069
rect 674326 555005 674378 555011
rect 674338 541176 674366 555005
rect 674998 553953 675050 553959
rect 674998 553895 675050 553901
rect 674902 553213 674954 553219
rect 674902 553155 674954 553161
rect 674518 551955 674570 551961
rect 674518 551897 674570 551903
rect 674422 541373 674474 541379
rect 674420 541338 674422 541347
rect 674474 541338 674476 541347
rect 674420 541273 674476 541282
rect 674338 541148 674462 541176
rect 674326 541077 674378 541083
rect 674326 541019 674378 541025
rect 674230 497935 674282 497941
rect 669910 496529 669962 496535
rect 669910 496471 669962 496477
rect 674050 486143 674078 497932
rect 674230 497877 674282 497883
rect 674338 497812 674366 541019
rect 674146 497784 674366 497812
rect 674036 486134 674092 486143
rect 674036 486069 674092 486078
rect 674146 484663 674174 497784
rect 674230 497713 674282 497719
rect 674230 497655 674282 497661
rect 674242 490139 674270 497655
rect 674326 497639 674378 497645
rect 674326 497581 674378 497587
rect 674228 490130 674284 490139
rect 674228 490065 674284 490074
rect 674338 485329 674366 497581
rect 674434 497516 674462 541148
rect 674530 497645 674558 551897
rect 674614 550105 674666 550111
rect 674614 550047 674666 550053
rect 674518 497639 674570 497645
rect 674518 497581 674570 497587
rect 674434 497488 674558 497516
rect 674422 497343 674474 497349
rect 674420 497308 674422 497317
rect 674474 497308 674476 497317
rect 674420 497243 674476 497252
rect 674422 496529 674474 496535
rect 674420 496494 674422 496503
rect 674474 496494 674476 496503
rect 674420 496429 674476 496438
rect 674530 489695 674558 497488
rect 674626 491915 674654 550047
rect 674806 548255 674858 548261
rect 674806 548197 674858 548203
rect 674708 541634 674764 541643
rect 674708 541569 674764 541578
rect 674722 541527 674750 541569
rect 674710 541521 674762 541527
rect 674710 541463 674762 541469
rect 674710 540781 674762 540787
rect 674708 540746 674710 540755
rect 674762 540746 674764 540755
rect 674708 540681 674764 540690
rect 674710 539893 674762 539899
rect 674708 539858 674710 539867
rect 674762 539858 674764 539867
rect 674708 539793 674764 539802
rect 674818 539696 674846 548197
rect 674722 539668 674846 539696
rect 674722 497941 674750 539668
rect 674804 537638 674860 537647
rect 674804 537573 674860 537582
rect 674710 497935 674762 497941
rect 674710 497877 674762 497883
rect 674708 497826 674764 497835
rect 674708 497761 674764 497770
rect 674722 495573 674750 497761
rect 674710 495567 674762 495573
rect 674710 495509 674762 495515
rect 674818 494315 674846 537573
rect 674914 518384 674942 553155
rect 675010 541083 675038 553895
rect 675202 551591 675230 555819
rect 675490 555069 675518 555444
rect 675478 555063 675530 555069
rect 675478 555005 675530 555011
rect 675394 554551 675422 554926
rect 675382 554545 675434 554551
rect 675382 554487 675434 554493
rect 675490 553959 675518 554260
rect 675478 553953 675530 553959
rect 675478 553895 675530 553901
rect 675394 553219 675422 553631
rect 675382 553213 675434 553219
rect 675382 553155 675434 553161
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 675190 551585 675242 551591
rect 675190 551527 675242 551533
rect 675382 551585 675434 551591
rect 675382 551527 675434 551533
rect 675394 551226 675422 551527
rect 675490 550111 675518 550595
rect 675478 550105 675530 550111
rect 675478 550047 675530 550053
rect 675394 548261 675422 548755
rect 675382 548255 675434 548261
rect 675382 548197 675434 548203
rect 679796 547110 679852 547119
rect 679796 547045 679852 547054
rect 674998 541077 675050 541083
rect 674998 541019 675050 541025
rect 676724 538674 676780 538683
rect 676724 538609 676780 538618
rect 676630 535749 676682 535755
rect 676630 535691 676682 535697
rect 674914 518356 675038 518384
rect 675010 498256 675038 518356
rect 675010 498228 675134 498256
rect 674998 498083 675050 498089
rect 674998 498025 675050 498031
rect 674902 497935 674954 497941
rect 674902 497877 674954 497883
rect 674806 494309 674858 494315
rect 674806 494251 674858 494257
rect 674612 491906 674668 491915
rect 674612 491841 674668 491850
rect 674516 489686 674572 489695
rect 674516 489621 674572 489630
rect 674914 488807 674942 497877
rect 674900 488798 674956 488807
rect 674900 488733 674956 488742
rect 674324 485320 674380 485329
rect 674324 485255 674380 485264
rect 674132 484654 674188 484663
rect 674132 484589 674188 484598
rect 675010 483183 675038 498025
rect 674996 483174 675052 483183
rect 674996 483109 675052 483118
rect 675106 482443 675134 498228
rect 676642 493099 676670 535691
rect 676738 495911 676766 538609
rect 679810 537647 679838 547045
rect 679796 537638 679852 537647
rect 679796 537573 679852 537582
rect 679810 535755 679838 537573
rect 679798 535749 679850 535755
rect 679798 535691 679850 535697
rect 679796 524762 679852 524771
rect 679796 524697 679852 524706
rect 679810 524179 679838 524697
rect 679796 524170 679852 524179
rect 679796 524105 679852 524114
rect 679810 521325 679838 524105
rect 679798 521319 679850 521325
rect 679798 521261 679850 521267
rect 676724 495902 676780 495911
rect 676724 495837 676780 495846
rect 676724 494570 676780 494579
rect 676724 494505 676780 494514
rect 676628 493090 676684 493099
rect 676628 493025 676684 493034
rect 675092 482434 675148 482443
rect 675092 482369 675148 482378
rect 676642 411995 676670 493025
rect 676628 411986 676684 411995
rect 676628 411921 676684 411930
rect 674422 409949 674474 409955
rect 674420 409914 674422 409923
rect 674474 409914 674476 409923
rect 674420 409849 674476 409858
rect 674710 409357 674762 409363
rect 674708 409322 674710 409331
rect 674762 409322 674764 409331
rect 674708 409257 674764 409266
rect 674710 408469 674762 408475
rect 674708 408434 674710 408443
rect 674762 408434 674764 408443
rect 674708 408369 674764 408378
rect 676738 407703 676766 494505
rect 679700 494422 679756 494431
rect 679700 494357 679756 494366
rect 679714 494315 679742 494357
rect 679702 494309 679754 494315
rect 679702 494251 679754 494257
rect 679892 493534 679948 493543
rect 679892 493469 679948 493478
rect 679796 480806 679852 480815
rect 679796 480741 679852 480750
rect 679810 480075 679838 480741
rect 679796 480066 679852 480075
rect 679796 480001 679852 480010
rect 679810 478183 679838 480001
rect 679798 478177 679850 478183
rect 679798 478119 679850 478125
rect 679906 475339 679934 493469
rect 679892 475330 679948 475339
rect 679892 475265 679948 475274
rect 676724 407694 676780 407703
rect 676724 407629 676780 407638
rect 673844 406658 673900 406667
rect 673844 406593 673900 406602
rect 669814 363329 669866 363335
rect 669814 363271 669866 363277
rect 673858 362267 673886 406593
rect 674900 404142 674956 404151
rect 674900 404077 674956 404086
rect 674132 401922 674188 401931
rect 674132 401857 674188 401866
rect 674036 397186 674092 397195
rect 674036 397121 674092 397130
rect 674050 375767 674078 397121
rect 674146 383167 674174 401857
rect 674612 398518 674668 398527
rect 674612 398453 674668 398462
rect 674324 397926 674380 397935
rect 674324 397861 674380 397870
rect 674338 384351 674366 397861
rect 674420 396446 674476 396455
rect 674420 396381 674476 396390
rect 674326 384345 674378 384351
rect 674326 384287 674378 384293
rect 674134 383161 674186 383167
rect 674134 383103 674186 383109
rect 674434 377617 674462 396381
rect 674516 393782 674572 393791
rect 674516 393717 674572 393726
rect 674422 377611 674474 377617
rect 674422 377553 674474 377559
rect 674530 376877 674558 393717
rect 674626 382501 674654 398453
rect 674804 395410 674860 395419
rect 674804 395345 674860 395354
rect 674708 394522 674764 394531
rect 674708 394457 674764 394466
rect 674614 382495 674666 382501
rect 674614 382437 674666 382443
rect 674722 378209 674750 394457
rect 674818 381336 674846 395345
rect 674914 384444 674942 404077
rect 675380 402514 675436 402523
rect 675380 402449 675436 402458
rect 675284 399406 675340 399415
rect 675284 399341 675340 399350
rect 675298 391696 675326 399341
rect 675202 391668 675326 391696
rect 675202 385110 675230 391668
rect 675394 391548 675422 402449
rect 679796 392598 679852 392607
rect 679796 392533 679852 392542
rect 679810 392163 679838 392533
rect 679796 392154 679852 392163
rect 679796 392089 679852 392098
rect 679810 391751 679838 392089
rect 679798 391745 679850 391751
rect 679798 391687 679850 391693
rect 675298 391520 675422 391548
rect 675298 385737 675326 391520
rect 675298 385709 675408 385737
rect 675202 385082 675326 385110
rect 675298 385036 675326 385082
rect 675394 385036 675422 385096
rect 675298 385008 675422 385036
rect 674914 384416 675408 384444
rect 675094 384345 675146 384351
rect 675094 384287 675146 384293
rect 675106 381410 675134 384287
rect 675382 383161 675434 383167
rect 675382 383103 675434 383109
rect 675394 382580 675422 383103
rect 675478 382495 675530 382501
rect 675478 382437 675530 382443
rect 675490 382062 675518 382437
rect 675106 381382 675408 381410
rect 674818 381308 675422 381336
rect 675394 380730 675422 381308
rect 675106 380198 675408 380226
rect 674710 378203 674762 378209
rect 674710 378145 674762 378151
rect 674518 376871 674570 376877
rect 674518 376813 674570 376819
rect 674038 375761 674090 375767
rect 674038 375703 674090 375709
rect 675106 374551 675134 380198
rect 675202 379532 675408 379560
rect 675092 374542 675148 374551
rect 675092 374477 675148 374486
rect 675202 371591 675230 379532
rect 675476 378834 675532 378843
rect 675476 378769 675532 378778
rect 675490 378288 675518 378769
rect 675382 378203 675434 378209
rect 675382 378145 675434 378151
rect 675394 377696 675422 378145
rect 675382 377611 675434 377617
rect 675382 377553 675434 377559
rect 675394 377075 675422 377553
rect 675478 376871 675530 376877
rect 675478 376813 675530 376819
rect 675490 376438 675518 376813
rect 675478 375761 675530 375767
rect 675478 375703 675530 375709
rect 675490 375254 675518 375703
rect 675476 373950 675532 373959
rect 675476 373885 675532 373894
rect 675490 373404 675518 373885
rect 675380 372026 675436 372035
rect 675380 371961 675436 371970
rect 675188 371582 675244 371591
rect 675394 371554 675422 371961
rect 675188 371517 675244 371526
rect 674708 364478 674764 364487
rect 674708 364413 674764 364422
rect 674422 363921 674474 363927
rect 674420 363886 674422 363895
rect 674474 363886 674476 363895
rect 674420 363821 674476 363830
rect 674614 363329 674666 363335
rect 674612 363294 674614 363303
rect 674666 363294 674668 363303
rect 674612 363229 674668 363238
rect 674722 363113 674750 364413
rect 674710 363107 674762 363113
rect 674710 363049 674762 363055
rect 673844 362258 673900 362267
rect 673844 362193 673900 362202
rect 679892 360186 679948 360195
rect 679892 360121 679948 360130
rect 674036 359150 674092 359159
rect 674036 359085 674092 359094
rect 674050 339581 674078 359085
rect 674516 357226 674572 357235
rect 674516 357161 674572 357170
rect 674324 352786 674380 352795
rect 674324 352721 674380 352730
rect 674228 351306 674284 351315
rect 674228 351241 674284 351250
rect 674038 339575 674090 339581
rect 674038 339517 674090 339523
rect 674242 332255 674270 351241
rect 674338 336621 674366 352721
rect 674530 340987 674558 357161
rect 675188 356486 675244 356495
rect 675188 356421 675244 356430
rect 675092 353378 675148 353387
rect 675092 353313 675148 353322
rect 674900 350270 674956 350279
rect 674900 350205 674956 350214
rect 674708 349382 674764 349391
rect 674708 349317 674764 349326
rect 674518 340981 674570 340987
rect 674518 340923 674570 340929
rect 674326 336615 674378 336621
rect 674326 336557 674378 336563
rect 674722 332773 674750 349317
rect 674914 336325 674942 350205
rect 674996 348642 675052 348651
rect 674996 348577 675052 348586
rect 674902 336319 674954 336325
rect 674902 336261 674954 336267
rect 674710 332767 674762 332773
rect 674710 332709 674762 332715
rect 674230 332249 674282 332255
rect 674230 332191 674282 332197
rect 675010 331811 675038 348577
rect 675106 336862 675134 353313
rect 675202 337409 675230 356421
rect 675284 354118 675340 354127
rect 675284 354053 675340 354062
rect 675298 339896 675326 354053
rect 679796 347458 679852 347467
rect 679796 347393 679852 347402
rect 679810 346727 679838 347393
rect 679796 346718 679852 346727
rect 679796 346653 679852 346662
rect 679810 345649 679838 346653
rect 679798 345643 679850 345649
rect 679798 345585 679850 345591
rect 679906 345543 679934 360121
rect 679892 345534 679948 345543
rect 679892 345469 679948 345478
rect 675478 340981 675530 340987
rect 675478 340923 675530 340929
rect 675490 340548 675518 340923
rect 675298 339868 675408 339896
rect 675382 339575 675434 339581
rect 675382 339517 675434 339523
rect 675394 339216 675422 339517
rect 675202 337381 675408 337409
rect 675106 336834 675408 336862
rect 675382 336615 675434 336621
rect 675382 336557 675434 336563
rect 675094 336319 675146 336325
rect 675094 336261 675146 336267
rect 675106 335569 675134 336261
rect 675394 336182 675422 336557
rect 675106 335541 675408 335569
rect 675476 335174 675532 335183
rect 675476 335109 675532 335118
rect 675490 335012 675518 335109
rect 675202 334998 675518 335012
rect 675202 334984 675504 334998
rect 674998 331805 675050 331811
rect 674998 331747 675050 331753
rect 675202 329559 675230 334984
rect 675490 333851 675518 334332
rect 675476 333842 675532 333851
rect 675476 333777 675532 333786
rect 675380 333546 675436 333555
rect 675380 333481 675436 333490
rect 675394 333074 675422 333481
rect 675382 332767 675434 332773
rect 675382 332709 675434 332715
rect 675394 332519 675422 332709
rect 675478 332249 675530 332255
rect 675478 332191 675530 332197
rect 675490 331890 675518 332191
rect 675382 331805 675434 331811
rect 675382 331747 675434 331753
rect 675394 331224 675422 331747
rect 675476 330586 675532 330595
rect 675476 330521 675532 330530
rect 675490 330040 675518 330521
rect 675188 329550 675244 329559
rect 675188 329485 675244 329494
rect 675380 328366 675436 328375
rect 675380 328301 675436 328310
rect 675394 328190 675422 328301
rect 675380 326886 675436 326895
rect 675380 326821 675436 326830
rect 675394 326340 675422 326821
rect 674710 319965 674762 319971
rect 674708 319930 674710 319939
rect 674762 319930 674764 319939
rect 674708 319865 674764 319874
rect 674422 318929 674474 318935
rect 674420 318894 674422 318903
rect 674474 318894 674476 318903
rect 674420 318829 674476 318838
rect 674710 318337 674762 318343
rect 674708 318302 674710 318311
rect 674762 318302 674764 318311
rect 674708 318237 674764 318246
rect 677012 313862 677068 313871
rect 677012 313797 677068 313806
rect 674324 312530 674380 312539
rect 674324 312465 674380 312474
rect 673940 306166 673996 306175
rect 673940 306101 673996 306110
rect 673954 287263 673982 306101
rect 674036 304538 674092 304547
rect 674036 304473 674092 304482
rect 674050 287781 674078 304473
rect 674228 303798 674284 303807
rect 674228 303733 674284 303742
rect 674038 287775 674090 287781
rect 674038 287717 674090 287723
rect 673942 287257 673994 287263
rect 673942 287199 673994 287205
rect 674242 286819 674270 303733
rect 674338 295995 674366 312465
rect 676916 311494 676972 311503
rect 676916 311429 676972 311438
rect 676820 310754 676876 310763
rect 676820 310689 676876 310698
rect 674612 309126 674668 309135
rect 674612 309061 674668 309070
rect 674420 308534 674476 308543
rect 674420 308469 674476 308478
rect 674326 295989 674378 295995
rect 674326 295931 674378 295937
rect 674434 292739 674462 308469
rect 674626 295403 674654 309061
rect 675092 307498 675148 307507
rect 675092 307433 675148 307442
rect 674996 305278 675052 305287
rect 674996 305213 675052 305222
rect 674902 299541 674954 299547
rect 674902 299483 674954 299489
rect 674614 295397 674666 295403
rect 674614 295339 674666 295345
rect 674422 292733 674474 292739
rect 674422 292675 674474 292681
rect 674914 288595 674942 299483
rect 675010 290569 675038 305213
rect 675106 291204 675134 307433
rect 676834 299547 676862 310689
rect 676822 299541 676874 299547
rect 676822 299483 676874 299489
rect 676930 299473 676958 311429
rect 675190 299467 675242 299473
rect 675190 299409 675242 299415
rect 676918 299467 676970 299473
rect 676918 299409 676970 299415
rect 675202 292832 675230 299409
rect 677026 299399 677054 313797
rect 679796 302466 679852 302475
rect 679796 302401 679852 302410
rect 679810 301735 679838 302401
rect 679796 301726 679852 301735
rect 679796 301661 679852 301670
rect 679810 299621 679838 301661
rect 679798 299615 679850 299621
rect 679798 299557 679850 299563
rect 675286 299393 675338 299399
rect 675286 299335 675338 299341
rect 677014 299393 677066 299399
rect 677014 299335 677066 299341
rect 675298 294238 675326 299335
rect 675382 295989 675434 295995
rect 675382 295931 675434 295937
rect 675394 295523 675422 295931
rect 675478 295397 675530 295403
rect 675478 295339 675530 295345
rect 675490 294890 675518 295339
rect 675298 294210 675408 294238
rect 675202 292804 675422 292832
rect 675190 292733 675242 292739
rect 675190 292675 675242 292681
rect 675202 291870 675230 292675
rect 675394 292374 675422 292804
rect 675202 291842 675408 291870
rect 675106 291176 675408 291204
rect 675010 290541 675408 290569
rect 675476 290182 675532 290191
rect 675476 290117 675532 290126
rect 675490 290020 675518 290117
rect 675010 290006 675518 290020
rect 675010 289992 675504 290006
rect 674902 288589 674954 288595
rect 674902 288531 674954 288537
rect 674230 286813 674282 286819
rect 674230 286755 674282 286761
rect 675010 282347 675038 289992
rect 675380 289590 675436 289599
rect 675380 289525 675436 289534
rect 675394 289354 675422 289525
rect 675394 289340 675504 289354
rect 675408 289326 675518 289340
rect 675490 288836 675518 289326
rect 675202 288808 675518 288836
rect 674996 282338 675052 282347
rect 674996 282273 675052 282282
rect 669718 274973 669770 274979
rect 674710 274973 674762 274979
rect 669718 274915 669770 274921
rect 674708 274938 674710 274947
rect 674762 274938 674764 274947
rect 674708 274873 674764 274882
rect 675202 274355 675230 288808
rect 675478 288589 675530 288595
rect 675478 288531 675530 288537
rect 675490 288082 675518 288531
rect 675382 287775 675434 287781
rect 675382 287717 675434 287723
rect 675394 287519 675422 287717
rect 675478 287257 675530 287263
rect 675478 287199 675530 287205
rect 675490 286898 675518 287199
rect 675382 286813 675434 286819
rect 675382 286755 675434 286761
rect 675394 286232 675422 286755
rect 675476 285298 675532 285307
rect 675476 285233 675532 285242
rect 675490 285048 675518 285233
rect 675380 283670 675436 283679
rect 675380 283605 675436 283614
rect 675394 283198 675422 283605
rect 675380 281894 675436 281903
rect 675380 281829 675436 281838
rect 675394 281348 675422 281829
rect 675188 274346 675244 274355
rect 675188 274281 675244 274290
rect 674710 274085 674762 274091
rect 674708 274050 674710 274059
rect 674762 274050 674764 274059
rect 674708 273985 674764 273994
rect 675202 273615 675230 274281
rect 675188 273606 675244 273615
rect 675188 273541 675244 273550
rect 674710 273345 674762 273351
rect 674708 273310 674710 273319
rect 674762 273310 674764 273319
rect 674708 273245 674764 273254
rect 674804 272718 674860 272727
rect 674804 272653 674860 272662
rect 674420 262802 674476 262811
rect 674420 262737 674476 262746
rect 674132 261174 674188 261183
rect 674132 261109 674188 261118
rect 671062 255733 671114 255739
rect 671060 255698 671062 255707
rect 671114 255698 671116 255707
rect 671060 255633 671116 255642
rect 674146 242419 674174 261109
rect 674324 258806 674380 258815
rect 674324 258741 674380 258750
rect 674134 242413 674186 242419
rect 674134 242355 674186 242361
rect 674338 241753 674366 258741
rect 674434 246785 674462 262737
rect 674818 262219 674846 272653
rect 680084 270942 680140 270951
rect 680084 270877 680140 270886
rect 675380 267242 675436 267251
rect 675380 267177 675436 267186
rect 675284 264134 675340 264143
rect 675284 264069 675340 264078
rect 675188 263394 675244 263403
rect 675188 263329 675244 263338
rect 674804 262210 674860 262219
rect 674804 262145 674860 262154
rect 674900 261766 674956 261775
rect 674900 261701 674956 261710
rect 674806 253439 674858 253445
rect 674806 253381 674858 253387
rect 674818 250263 674846 253381
rect 674806 250257 674858 250263
rect 674806 250199 674858 250205
rect 674422 246779 674474 246785
rect 674422 246721 674474 246727
rect 674326 241747 674378 241753
rect 674326 241689 674378 241695
rect 674914 240569 674942 261701
rect 675092 260138 675148 260147
rect 675092 260073 675148 260082
rect 674996 259398 675052 259407
rect 674996 259333 675052 259342
rect 675010 243011 675038 259333
rect 675106 245546 675134 260073
rect 675202 246878 675230 263329
rect 675298 250356 675326 264069
rect 675394 251225 675422 267177
rect 676820 266502 676876 266511
rect 676820 266437 676876 266446
rect 676834 253445 676862 266437
rect 679700 257474 679756 257483
rect 679700 257409 679756 257418
rect 679714 256891 679742 257409
rect 679700 256882 679756 256891
rect 679700 256817 679756 256826
rect 679714 256405 679742 256817
rect 679702 256399 679754 256405
rect 679702 256341 679754 256347
rect 680098 256299 680126 270877
rect 680084 256290 680140 256299
rect 680084 256225 680140 256234
rect 676822 253439 676874 253445
rect 676822 253381 676874 253387
rect 675382 251219 675434 251225
rect 675382 251161 675434 251167
rect 675382 250997 675434 251003
rect 675382 250939 675434 250945
rect 675394 250523 675422 250939
rect 675298 250328 675518 250356
rect 675286 250257 675338 250263
rect 675286 250199 675338 250205
rect 675298 247396 675326 250199
rect 675490 249898 675518 250328
rect 675380 249630 675436 249639
rect 675380 249565 675436 249574
rect 675394 249232 675422 249565
rect 675298 247368 675408 247396
rect 675202 246850 675326 246878
rect 675298 246804 675326 246850
rect 675394 246804 675422 246864
rect 675190 246779 675242 246785
rect 675298 246776 675422 246804
rect 675190 246721 675242 246727
rect 675202 246212 675230 246721
rect 675202 246184 675408 246212
rect 675298 245592 675422 245620
rect 675298 245546 675326 245592
rect 675106 245518 675326 245546
rect 675394 245532 675422 245592
rect 675284 245042 675340 245051
rect 675340 245000 675408 245028
rect 675284 244977 675340 244986
rect 675476 244746 675532 244755
rect 675476 244681 675532 244690
rect 675490 244362 675518 244681
rect 675106 244348 675518 244362
rect 675106 244334 675504 244348
rect 674998 243005 675050 243011
rect 674998 242947 675050 242953
rect 674902 240563 674954 240569
rect 674902 240505 674954 240511
rect 675106 238983 675134 244334
rect 675476 243562 675532 243571
rect 675476 243497 675532 243506
rect 675490 243090 675518 243497
rect 675382 243005 675434 243011
rect 675382 242947 675434 242953
rect 675394 242498 675422 242947
rect 675382 242413 675434 242419
rect 675382 242355 675434 242361
rect 675394 241875 675422 242355
rect 675478 241747 675530 241753
rect 675478 241689 675530 241695
rect 675490 241240 675518 241689
rect 675478 240563 675530 240569
rect 675478 240505 675530 240511
rect 675490 240056 675518 240505
rect 675092 238974 675148 238983
rect 675092 238909 675148 238918
rect 675668 238678 675724 238687
rect 675668 238613 675724 238622
rect 675682 238206 675710 238613
rect 675380 236902 675436 236911
rect 675380 236837 675436 236846
rect 675394 236356 675422 236837
rect 674422 229537 674474 229543
rect 674420 229502 674422 229511
rect 674474 229502 674476 229511
rect 674420 229437 674476 229446
rect 674710 228945 674762 228951
rect 674708 228910 674710 228919
rect 674762 228910 674764 228919
rect 674708 228845 674764 228854
rect 669622 227909 669674 227915
rect 674422 227909 674474 227915
rect 669622 227851 669674 227857
rect 674420 227874 674422 227883
rect 674474 227874 674476 227883
rect 674420 227809 674476 227818
rect 679796 225062 679852 225071
rect 679796 224997 679852 225006
rect 676820 223730 676876 223739
rect 676820 223665 676876 223674
rect 674516 222102 674572 222111
rect 674516 222037 674572 222046
rect 674420 217514 674476 217523
rect 674420 217449 674476 217458
rect 674132 216034 674188 216043
rect 674132 215969 674188 215978
rect 674146 197057 674174 215969
rect 674434 201349 674462 217449
rect 674530 205789 674558 222037
rect 674996 221214 675052 221223
rect 674996 221149 675052 221158
rect 674612 221066 674668 221075
rect 674612 221001 674668 221010
rect 674518 205783 674570 205789
rect 674518 205725 674570 205731
rect 674626 201687 674654 221001
rect 674900 214998 674956 215007
rect 674900 214933 674956 214942
rect 674804 214258 674860 214267
rect 674804 214193 674860 214202
rect 674708 213370 674764 213379
rect 674708 213305 674764 213314
rect 674612 201678 674668 201687
rect 674612 201613 674668 201622
rect 674422 201343 674474 201349
rect 674422 201285 674474 201291
rect 674134 197051 674186 197057
rect 674134 196993 674186 196999
rect 674722 196613 674750 213305
rect 674818 197649 674846 214193
rect 674914 200369 674942 214933
rect 675010 204920 675038 221149
rect 675188 218994 675244 219003
rect 675188 218929 675244 218938
rect 675092 218106 675148 218115
rect 675092 218041 675148 218050
rect 675106 205049 675134 218041
rect 675202 205049 675230 218929
rect 676834 206275 676862 223665
rect 679700 212186 679756 212195
rect 679700 212121 679756 212130
rect 679714 211455 679742 212121
rect 679700 211446 679756 211455
rect 679700 211381 679756 211390
rect 679714 210303 679742 211381
rect 679702 210297 679754 210303
rect 679702 210239 679754 210245
rect 679810 210123 679838 224997
rect 679796 210114 679852 210123
rect 679796 210049 679852 210058
rect 676820 206266 676876 206275
rect 676820 206201 676876 206210
rect 675478 205783 675530 205789
rect 675478 205725 675530 205731
rect 675490 205350 675518 205725
rect 675094 205043 675146 205049
rect 675094 204985 675146 204991
rect 675190 205043 675242 205049
rect 675190 204985 675242 204991
rect 675478 205043 675530 205049
rect 675478 204985 675530 204991
rect 675010 204892 675230 204920
rect 674998 204821 675050 204827
rect 674998 204763 675050 204769
rect 675010 201664 675038 204763
rect 675202 202182 675230 204892
rect 675490 204684 675518 204985
rect 675764 204490 675820 204499
rect 675764 204425 675820 204434
rect 675778 204018 675806 204425
rect 675298 202228 675422 202256
rect 675298 202182 675326 202228
rect 675202 202154 675326 202182
rect 675394 202168 675422 202228
rect 675010 201636 675408 201664
rect 675382 201343 675434 201349
rect 675382 201285 675434 201291
rect 675394 200984 675422 201285
rect 674914 200341 675408 200369
rect 675476 200050 675532 200059
rect 675476 199985 675532 199994
rect 675490 199814 675518 199985
rect 675106 199800 675518 199814
rect 675106 199786 675504 199800
rect 674806 197643 674858 197649
rect 674806 197585 674858 197591
rect 674710 196607 674762 196613
rect 674710 196549 674762 196555
rect 675106 193251 675134 199786
rect 675380 199458 675436 199467
rect 675380 199393 675436 199402
rect 675394 199296 675422 199393
rect 675298 199268 675422 199296
rect 675298 199148 675326 199268
rect 675202 199120 675326 199148
rect 675394 199134 675422 199268
rect 675092 193242 675148 193251
rect 675092 193177 675148 193186
rect 675202 193103 675230 199120
rect 675476 198422 675532 198431
rect 675476 198357 675532 198366
rect 675490 197876 675518 198357
rect 675382 197643 675434 197649
rect 675382 197585 675434 197591
rect 675394 197319 675422 197585
rect 675478 197051 675530 197057
rect 675478 196993 675530 196999
rect 675490 196692 675518 196993
rect 675382 196607 675434 196613
rect 675382 196549 675434 196555
rect 675394 196026 675422 196549
rect 675476 195314 675532 195323
rect 675476 195249 675532 195258
rect 675490 194842 675518 195249
rect 675380 193538 675436 193547
rect 675380 193473 675436 193482
rect 675188 193094 675244 193103
rect 675188 193029 675244 193038
rect 675394 192992 675422 193473
rect 675380 191614 675436 191623
rect 675380 191549 675436 191558
rect 675394 191142 675422 191549
rect 674420 184510 674476 184519
rect 674420 184445 674476 184454
rect 674434 184403 674462 184445
rect 674422 184397 674474 184403
rect 674422 184339 674474 184345
rect 674710 183953 674762 183959
rect 674708 183918 674710 183927
rect 674762 183918 674764 183927
rect 674708 183853 674764 183862
rect 666742 182917 666794 182923
rect 674422 182917 674474 182923
rect 666742 182859 666794 182865
rect 674420 182882 674422 182891
rect 674474 182882 674476 182891
rect 674420 182817 674476 182826
rect 676916 178738 676972 178747
rect 676916 178673 676972 178682
rect 674516 177110 674572 177119
rect 674516 177045 674572 177054
rect 674036 171042 674092 171051
rect 674036 170977 674092 170986
rect 674050 152065 674078 170977
rect 674228 169414 674284 169423
rect 674228 169349 674284 169358
rect 674242 152657 674270 169349
rect 674530 168512 674558 177045
rect 676820 176222 676876 176231
rect 676820 176157 676876 176166
rect 675668 174002 675724 174011
rect 675668 173937 675724 173946
rect 674900 173114 674956 173123
rect 674900 173049 674956 173058
rect 674434 168484 674558 168512
rect 674434 160797 674462 168484
rect 674516 168378 674572 168387
rect 674516 168313 674572 168322
rect 674422 160791 674474 160797
rect 674422 160733 674474 160739
rect 674230 152651 674282 152657
rect 674230 152593 674282 152599
rect 674038 152059 674090 152065
rect 674038 152001 674090 152007
rect 674530 151547 674558 168313
rect 674708 167342 674764 167351
rect 674708 167277 674764 167286
rect 674722 167235 674750 167277
rect 674710 167229 674762 167235
rect 674710 167171 674762 167177
rect 674612 166750 674668 166759
rect 674612 166685 674668 166694
rect 674626 164201 674654 166685
rect 674708 165714 674764 165723
rect 674708 165649 674764 165658
rect 674722 164275 674750 165649
rect 674710 164269 674762 164275
rect 674710 164211 674762 164217
rect 674614 164195 674666 164201
rect 674614 164137 674666 164143
rect 674914 162592 674942 173049
rect 674996 172374 675052 172383
rect 674996 172309 675052 172318
rect 674818 162564 674942 162592
rect 674818 156949 674846 162564
rect 675010 162444 675038 172309
rect 675092 170006 675148 170015
rect 675092 169941 675148 169950
rect 674914 162416 675038 162444
rect 674914 157097 674942 162416
rect 675106 162296 675134 169941
rect 675190 163085 675242 163091
rect 675190 163027 675242 163033
rect 675010 162268 675134 162296
rect 674902 157091 674954 157097
rect 674902 157033 674954 157039
rect 674806 156943 674858 156949
rect 674806 156885 674858 156891
rect 675010 155369 675038 162268
rect 675094 162123 675146 162129
rect 675094 162065 675146 162071
rect 675106 157190 675134 162065
rect 675202 159040 675230 163027
rect 675682 161019 675710 173937
rect 676834 162129 676862 176157
rect 676930 163091 676958 178673
rect 677012 175630 677068 175639
rect 677012 175565 677068 175574
rect 676918 163085 676970 163091
rect 676918 163027 676970 163033
rect 676822 162123 676874 162129
rect 676822 162065 676874 162071
rect 677026 161431 677054 175565
rect 677012 161422 677068 161431
rect 677012 161357 677068 161366
rect 675670 161013 675722 161019
rect 675670 160955 675722 160961
rect 675382 160791 675434 160797
rect 675382 160733 675434 160739
rect 675394 160323 675422 160733
rect 675670 160051 675722 160057
rect 675670 159993 675722 159999
rect 675682 159692 675710 159993
rect 675202 159012 675408 159040
rect 675106 157162 675326 157190
rect 675298 157116 675326 157162
rect 675490 157116 675518 157176
rect 675094 157091 675146 157097
rect 675298 157088 675518 157116
rect 675094 157033 675146 157039
rect 675106 156006 675134 157033
rect 675478 156943 675530 156949
rect 675478 156885 675530 156891
rect 675490 156658 675518 156885
rect 675106 155978 675408 156006
rect 675010 155341 675408 155369
rect 675284 155206 675340 155215
rect 675284 155141 675340 155150
rect 675298 154452 675326 155141
rect 675476 155058 675532 155067
rect 675476 154993 675532 155002
rect 675490 154808 675518 154993
rect 675298 154424 675422 154452
rect 675394 154142 675422 154424
rect 675764 153430 675820 153439
rect 675764 153365 675820 153374
rect 675778 152884 675806 153365
rect 675382 152651 675434 152657
rect 675382 152593 675434 152599
rect 675394 152292 675422 152593
rect 675478 152059 675530 152065
rect 675478 152001 675530 152007
rect 675490 151700 675518 152001
rect 674518 151541 674570 151547
rect 674518 151483 674570 151489
rect 675382 151541 675434 151547
rect 675382 151483 675434 151489
rect 675394 151034 675422 151483
rect 675476 150322 675532 150331
rect 675476 150257 675532 150266
rect 675490 149850 675518 150257
rect 675476 148546 675532 148555
rect 675476 148481 675532 148490
rect 675490 148000 675518 148481
rect 675380 146474 675436 146483
rect 675380 146409 675436 146418
rect 675394 146150 675422 146409
rect 674324 142774 674380 142783
rect 674324 142709 674380 142718
rect 674338 142667 674366 142709
rect 674326 142661 674378 142667
rect 674326 142603 674378 142609
rect 679702 142661 679754 142667
rect 679702 142603 679754 142609
rect 674708 138778 674764 138787
rect 674708 138713 674764 138722
rect 674722 138597 674750 138713
rect 674710 138591 674762 138597
rect 674710 138533 674762 138539
rect 674420 138482 674476 138491
rect 674420 138417 674422 138426
rect 674474 138417 674476 138426
rect 674422 138385 674474 138391
rect 674708 137150 674764 137159
rect 674708 137085 674764 137094
rect 674722 135637 674750 137085
rect 655414 135631 655466 135637
rect 655414 135573 655466 135579
rect 674710 135631 674762 135637
rect 674710 135573 674762 135579
rect 679714 135531 679742 142603
rect 674708 135522 674764 135531
rect 674708 135457 674764 135466
rect 679700 135522 679756 135531
rect 679700 135457 679756 135466
rect 674722 135415 674750 135457
rect 674710 135409 674762 135415
rect 674710 135351 674762 135357
rect 674420 134560 674476 134569
rect 674420 134495 674476 134504
rect 674434 132529 674462 134495
rect 675284 133450 675340 133459
rect 675284 133385 675340 133394
rect 643606 132523 643658 132529
rect 643606 132465 643658 132471
rect 674422 132523 674474 132529
rect 674422 132465 674474 132471
rect 675188 131822 675244 131831
rect 675188 131757 675244 131766
rect 674132 131230 674188 131239
rect 674132 131165 674188 131174
rect 673364 126790 673420 126799
rect 673420 126748 673486 126776
rect 673364 126725 673420 126734
rect 674036 125902 674092 125911
rect 674036 125837 674092 125846
rect 642068 121758 642124 121767
rect 642068 121693 642124 121702
rect 642082 121281 642110 121693
rect 642070 121275 642122 121281
rect 642070 121217 642122 121223
rect 642166 121201 642218 121207
rect 642164 121166 642166 121175
rect 642218 121166 642220 121175
rect 641398 121127 641450 121133
rect 642164 121101 642220 121110
rect 641398 121069 641450 121075
rect 641410 120731 641438 121069
rect 641396 120722 641452 120731
rect 641396 120657 641452 120666
rect 640724 120130 640780 120139
rect 640724 120065 640780 120074
rect 665204 112286 665260 112295
rect 665204 112221 665260 112230
rect 652534 100851 652586 100857
rect 652534 100793 652586 100799
rect 641014 92711 641066 92717
rect 641014 92653 641066 92659
rect 640726 92267 640778 92273
rect 640726 92209 640778 92215
rect 640630 81093 640682 81099
rect 640630 81035 640682 81041
rect 640642 80729 640670 81035
rect 640630 80723 640682 80729
rect 640630 80665 640682 80671
rect 640150 60447 640202 60453
rect 640150 60389 640202 60395
rect 640162 60347 640190 60389
rect 640148 60338 640204 60347
rect 640148 60273 640204 60282
rect 640738 55463 640766 92209
rect 640822 92193 640874 92199
rect 640822 92135 640874 92141
rect 640834 58719 640862 92135
rect 640918 86495 640970 86501
rect 640918 86437 640970 86443
rect 640820 58710 640876 58719
rect 640820 58645 640876 58654
rect 640930 57535 640958 86437
rect 641026 61383 641054 92653
rect 652546 87833 652574 100793
rect 665218 96491 665246 112221
rect 668180 111250 668236 111259
rect 668180 111185 668236 111194
rect 668194 100857 668222 111185
rect 674050 106925 674078 125837
rect 674146 118636 674174 131165
rect 675092 128714 675148 128723
rect 675092 128649 675148 128658
rect 674420 128122 674476 128131
rect 674420 128057 674476 128066
rect 674324 127382 674380 127391
rect 674324 127317 674380 127326
rect 674228 126494 674284 126503
rect 674228 126429 674284 126438
rect 674242 118784 674270 126429
rect 674338 118932 674366 127317
rect 674434 119080 674462 128057
rect 674996 124866 675052 124875
rect 674996 124801 675052 124810
rect 674900 123978 674956 123987
rect 674900 123913 674956 123922
rect 674516 123238 674572 123247
rect 674516 123173 674572 123182
rect 674530 119228 674558 123173
rect 674804 122202 674860 122211
rect 674804 122137 674860 122146
rect 674612 121610 674668 121619
rect 674612 121545 674668 121554
rect 674626 121133 674654 121545
rect 674708 121314 674764 121323
rect 674708 121249 674710 121258
rect 674762 121249 674764 121258
rect 674710 121217 674762 121223
rect 674818 121207 674846 122137
rect 674806 121201 674858 121207
rect 674806 121143 674858 121149
rect 674614 121127 674666 121133
rect 674614 121069 674666 121075
rect 674914 119672 674942 123913
rect 674818 119644 674942 119672
rect 674530 119200 674654 119228
rect 674434 119052 674558 119080
rect 674338 118904 674462 118932
rect 674242 118756 674366 118784
rect 674146 118608 674270 118636
rect 674134 118537 674186 118543
rect 674134 118479 674186 118485
rect 674146 114177 674174 118479
rect 674134 114171 674186 114177
rect 674134 114113 674186 114119
rect 674242 113659 674270 118608
rect 674230 113653 674282 113659
rect 674230 113595 674282 113601
rect 674038 106919 674090 106925
rect 674038 106861 674090 106867
rect 674338 105223 674366 118756
rect 674434 111217 674462 118904
rect 674530 113363 674558 119052
rect 674518 113357 674570 113363
rect 674518 113299 674570 113305
rect 674422 111211 674474 111217
rect 674422 111153 674474 111159
rect 674626 106407 674654 119200
rect 674818 107591 674846 119644
rect 674902 119573 674954 119579
rect 674902 119515 674954 119521
rect 674914 114843 674942 119515
rect 674902 114837 674954 114843
rect 674902 114779 674954 114785
rect 674900 110806 674956 110815
rect 674900 110741 674956 110750
rect 674914 109016 674942 110741
rect 675010 110169 675038 124801
rect 675106 119579 675134 128649
rect 675094 119573 675146 119579
rect 675094 119515 675146 119521
rect 675202 119376 675230 131757
rect 675106 119348 675230 119376
rect 675106 115158 675134 119348
rect 675298 118543 675326 133385
rect 675286 118537 675338 118543
rect 675286 118479 675338 118485
rect 675106 115130 675326 115158
rect 675298 115084 675326 115130
rect 675394 115084 675422 115144
rect 675298 115056 675422 115084
rect 675094 114837 675146 114843
rect 675094 114779 675146 114785
rect 675106 114492 675134 114779
rect 675106 114464 675408 114492
rect 675382 114171 675434 114177
rect 675382 114113 675434 114119
rect 675394 113812 675422 114113
rect 675190 113653 675242 113659
rect 675190 113595 675242 113601
rect 675094 113357 675146 113363
rect 675094 113299 675146 113305
rect 675106 111458 675134 113299
rect 675202 112009 675230 113595
rect 675202 111981 675408 112009
rect 675106 111430 675408 111458
rect 675382 111211 675434 111217
rect 675382 111153 675434 111159
rect 675394 110778 675422 111153
rect 675010 110141 675408 110169
rect 675572 110066 675628 110075
rect 675572 110001 675628 110010
rect 675586 109594 675614 110001
rect 674914 108988 675038 109016
rect 675010 108973 675038 108988
rect 675010 108945 675408 108973
rect 675380 108142 675436 108151
rect 675380 108077 675436 108086
rect 675394 107670 675422 108077
rect 674806 107585 674858 107591
rect 674806 107527 674858 107533
rect 675382 107585 675434 107591
rect 675382 107527 675434 107533
rect 675394 107119 675422 107527
rect 675478 106919 675530 106925
rect 675478 106861 675530 106867
rect 675490 106486 675518 106861
rect 674614 106401 674666 106407
rect 674614 106343 674666 106349
rect 675382 106401 675434 106407
rect 675382 106343 675434 106349
rect 675394 105820 675422 106343
rect 674326 105217 674378 105223
rect 674326 105159 674378 105165
rect 675382 105217 675434 105223
rect 675382 105159 675434 105165
rect 675394 104636 675422 105159
rect 675380 103258 675436 103267
rect 675380 103193 675436 103202
rect 675394 102786 675422 103193
rect 675380 101482 675436 101491
rect 675380 101417 675436 101426
rect 675394 100936 675422 101417
rect 668182 100851 668234 100857
rect 668182 100793 668234 100799
rect 663286 96485 663338 96491
rect 663286 96427 663338 96433
rect 665206 96485 665258 96491
rect 665206 96427 665258 96433
rect 662518 92859 662570 92865
rect 662518 92801 662570 92807
rect 659830 92711 659882 92717
rect 659830 92653 659882 92659
rect 658870 92637 658922 92643
rect 658870 92579 658922 92585
rect 658294 92563 658346 92569
rect 658294 92505 658346 92511
rect 657526 92193 657578 92199
rect 657526 92135 657578 92141
rect 657538 88000 657566 92135
rect 657538 87972 657792 88000
rect 658306 87986 658334 92505
rect 658882 87986 658910 92579
rect 659350 92489 659402 92495
rect 659350 92431 659402 92437
rect 659362 88000 659390 92431
rect 659842 88000 659870 92653
rect 661174 92415 661226 92421
rect 661174 92357 661226 92363
rect 660694 92341 660746 92347
rect 660694 92283 660746 92289
rect 659362 87972 659616 88000
rect 659842 87972 660144 88000
rect 660706 87986 660734 92283
rect 661186 88000 661214 92357
rect 661750 92267 661802 92273
rect 661750 92209 661802 92215
rect 661762 88000 661790 92209
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 92801
rect 663094 92785 663146 92791
rect 663094 92727 663146 92733
rect 663106 87986 663134 92727
rect 652534 87827 652586 87833
rect 652534 87769 652586 87775
rect 652628 86978 652684 86987
rect 652628 86913 652684 86922
rect 652642 86501 652670 86913
rect 652630 86495 652682 86501
rect 652630 86437 652682 86443
rect 653588 86238 653644 86247
rect 653588 86173 653644 86182
rect 653492 85350 653548 85359
rect 653492 85285 653548 85294
rect 641110 83757 641162 83763
rect 641110 83699 641162 83705
rect 641012 61374 641068 61383
rect 641012 61309 641068 61318
rect 640916 57526 640972 57535
rect 640916 57461 640972 57470
rect 641122 56499 641150 83699
rect 653506 83615 653534 85285
rect 653602 83763 653630 86173
rect 663298 85780 663326 96427
rect 663298 85752 663806 85780
rect 663380 85646 663436 85655
rect 663380 85581 663436 85590
rect 653684 84314 653740 84323
rect 653684 84249 653740 84258
rect 653590 83757 653642 83763
rect 653590 83699 653642 83705
rect 653698 83689 653726 84249
rect 663284 84018 663340 84027
rect 663202 83976 663284 84004
rect 653686 83683 653738 83689
rect 653686 83625 653738 83631
rect 653494 83609 653546 83615
rect 653494 83551 653546 83557
rect 653588 83426 653644 83435
rect 653588 83361 653644 83370
rect 641302 80945 641354 80951
rect 641302 80887 641354 80893
rect 641206 80797 641258 80803
rect 641206 80739 641258 80745
rect 641218 58127 641246 80739
rect 641204 58118 641260 58127
rect 641204 58053 641260 58062
rect 641314 57091 641342 80887
rect 653602 80729 653630 83361
rect 653684 82686 653740 82695
rect 653684 82621 653740 82630
rect 653698 80803 653726 82621
rect 662420 81206 662476 81215
rect 662420 81141 662476 81150
rect 656962 81016 657216 81044
rect 657538 81016 657792 81044
rect 653686 80797 653738 80803
rect 653686 80739 653738 80745
rect 641398 80723 641450 80729
rect 641398 80665 641450 80671
rect 653590 80723 653642 80729
rect 653590 80665 653642 80671
rect 641410 59607 641438 80665
rect 641494 77763 641546 77769
rect 641494 77705 641546 77711
rect 641396 59598 641452 59607
rect 641396 59533 641452 59542
rect 641300 57082 641356 57091
rect 641300 57017 641356 57026
rect 641108 56490 641164 56499
rect 641108 56425 641164 56434
rect 640724 55454 640780 55463
rect 640724 55389 640780 55398
rect 641506 54871 641534 77705
rect 642166 77689 642218 77695
rect 642166 77631 642218 77637
rect 641590 76949 641642 76955
rect 641590 76891 641642 76897
rect 641602 59755 641630 76891
rect 641686 76801 641738 76807
rect 641686 76743 641738 76749
rect 641588 59746 641644 59755
rect 641588 59681 641644 59690
rect 641698 56351 641726 76743
rect 642178 75591 642206 77631
rect 656962 76733 656990 81016
rect 657538 77769 657566 81016
rect 657526 77763 657578 77769
rect 657526 77705 657578 77711
rect 658306 76881 658334 81030
rect 658294 76875 658346 76881
rect 658294 76817 658346 76823
rect 658882 76807 658910 81030
rect 659602 80859 659630 81030
rect 659602 80831 659678 80859
rect 659650 76955 659678 80831
rect 659638 76949 659690 76955
rect 659638 76891 659690 76897
rect 658870 76801 658922 76807
rect 658870 76743 658922 76749
rect 656950 76727 657002 76733
rect 656950 76669 657002 76675
rect 660130 76437 660158 81030
rect 660706 76659 660734 81030
rect 661186 81016 661440 81044
rect 661762 81016 662016 81044
rect 660694 76653 660746 76659
rect 660694 76595 660746 76601
rect 661186 76585 661214 81016
rect 661174 76579 661226 76585
rect 661174 76521 661226 76527
rect 661762 76511 661790 81016
rect 662434 80877 662462 81141
rect 662422 80871 662474 80877
rect 662422 80813 662474 80819
rect 661750 76505 661802 76511
rect 661750 76447 661802 76453
rect 660118 76431 660170 76437
rect 660118 76373 660170 76379
rect 662530 76363 662558 81030
rect 662518 76357 662570 76363
rect 662518 76299 662570 76305
rect 642164 75582 642220 75591
rect 642164 75517 642220 75526
rect 641684 56342 641740 56351
rect 641684 56277 641740 56286
rect 641492 54862 641548 54871
rect 641492 54797 641548 54806
rect 639958 54675 640010 54681
rect 639958 54617 640010 54623
rect 639970 46911 639998 54617
rect 663202 47725 663230 83976
rect 663284 83953 663340 83962
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81099 663326 82029
rect 663286 81093 663338 81099
rect 663286 81035 663338 81041
rect 663394 48317 663422 85581
rect 663572 84758 663628 84767
rect 663572 84693 663628 84702
rect 663476 82834 663532 82843
rect 663476 82769 663532 82778
rect 663490 80951 663518 82769
rect 663478 80945 663530 80951
rect 663478 80887 663530 80893
rect 663586 60453 663614 84693
rect 663778 77695 663806 85752
rect 663766 77689 663818 77695
rect 663766 77631 663818 77637
rect 663574 60447 663626 60453
rect 663574 60389 663626 60395
rect 663382 48311 663434 48317
rect 663382 48253 663434 48259
rect 663190 47719 663242 47725
rect 663190 47661 663242 47667
rect 639958 46905 640010 46911
rect 639958 46847 640010 46853
rect 639862 46609 639914 46615
rect 639862 46551 639914 46557
rect 613462 44685 613514 44691
rect 613462 44627 613514 44633
rect 635542 44685 635594 44691
rect 635542 44627 635594 44633
rect 523892 43170 523948 43179
rect 523892 43105 523948 43114
rect 529268 43170 529324 43179
rect 529268 43105 529324 43114
rect 525908 42134 525964 42143
rect 521602 42092 521856 42120
rect 521204 42069 521260 42078
rect 525964 42092 526176 42120
rect 529282 42106 529310 43105
rect 525908 42069 525964 42078
rect 518516 41838 518572 41847
rect 514882 41805 515136 41824
rect 514870 41799 515136 41805
rect 514922 41796 515136 41799
rect 518572 41796 518832 41824
rect 518516 41773 518572 41782
rect 514870 41741 514922 41747
rect 512564 40802 512620 40811
rect 512564 40737 512620 40746
rect 499990 40393 500042 40399
rect 499990 40335 500042 40341
rect 512578 40325 512606 40737
rect 613474 40663 613502 44627
rect 613460 40654 613516 40663
rect 613460 40589 613516 40598
rect 512566 40319 512618 40325
rect 512566 40261 512618 40267
rect 446518 37433 446570 37439
rect 446518 37375 446570 37381
rect 459190 37433 459242 37439
rect 459190 37375 459242 37381
<< via2 >>
rect 41780 968706 41836 968762
rect 41780 967078 41836 967134
rect 41780 965006 41836 965062
rect 41780 963970 41836 964026
rect 41780 963378 41836 963434
rect 41780 962786 41836 962842
rect 41876 962194 41932 962250
rect 42356 962194 42412 962250
rect 42068 961750 42124 961806
rect 41780 959678 41836 959734
rect 41876 959086 41932 959142
rect 42068 958346 42124 958402
rect 42164 957754 42220 957810
rect 42164 956126 42220 956182
rect 42260 907473 42262 907490
rect 42262 907473 42314 907490
rect 42314 907473 42316 907490
rect 42260 907434 42316 907473
rect 42644 908065 42646 908082
rect 42646 908065 42698 908082
rect 42698 908065 42700 908082
rect 42644 908026 42700 908065
rect 42356 906694 42412 906750
rect 40340 905362 40396 905418
rect 40052 901366 40108 901422
rect 40148 842610 40204 842666
rect 39956 827514 40012 827570
rect 42644 904809 42646 904826
rect 42646 904809 42698 904826
rect 42698 904809 42700 904826
rect 42644 904770 42700 904809
rect 43124 907138 43180 907194
rect 43028 901070 43084 901126
rect 42932 897666 42988 897722
rect 42356 891154 42412 891210
rect 42356 889691 42412 889730
rect 42356 889674 42358 889691
rect 42358 889674 42410 889691
rect 42410 889674 42412 889691
rect 43220 904178 43276 904234
rect 44756 904178 44812 904234
rect 44564 903290 44620 903346
rect 43220 901514 43276 901570
rect 43124 887306 43180 887362
rect 40820 852674 40876 852730
rect 40340 820706 40396 820762
rect 42356 823853 42358 823870
rect 42358 823853 42410 823870
rect 42410 823853 42412 823870
rect 42356 823814 42412 823853
rect 42452 822630 42508 822686
rect 42356 822225 42358 822242
rect 42358 822225 42410 822242
rect 42410 822225 42412 822242
rect 42356 822186 42412 822225
rect 43220 821150 43276 821206
rect 40820 819522 40876 819578
rect 40148 819374 40204 819430
rect 42356 817894 42412 817950
rect 40244 816710 40300 816766
rect 37268 815822 37324 815878
rect 37364 812714 37420 812770
rect 37268 802058 37324 802114
rect 41972 814342 42028 814398
rect 41876 813602 41932 813658
rect 41684 811086 41740 811142
rect 37364 801910 37420 801966
rect 41780 809606 41836 809662
rect 41684 800430 41740 800486
rect 41780 800282 41836 800338
rect 42068 809162 42124 809218
rect 42164 808274 42220 808330
rect 42068 800282 42124 800338
rect 42260 805183 42316 805222
rect 42260 805166 42262 805183
rect 42262 805166 42314 805183
rect 42314 805166 42316 805183
rect 42452 815230 42508 815286
rect 43124 812270 43180 812326
rect 42932 807238 42988 807294
rect 42260 799986 42316 800042
rect 42452 797914 42508 797970
rect 41780 794214 41836 794270
rect 43124 810346 43180 810402
rect 42740 794806 42796 794862
rect 42260 792142 42316 792198
rect 41780 791106 41836 791162
rect 42164 790958 42220 791014
rect 42740 791994 42796 792050
rect 42452 791846 42508 791902
rect 42740 791698 42796 791754
rect 43124 791994 43180 792050
rect 42740 780467 42796 780506
rect 42740 780450 42742 780467
rect 42742 780450 42794 780467
rect 42794 780450 42796 780467
rect 42452 779897 42454 779914
rect 42454 779897 42506 779914
rect 42506 779897 42508 779914
rect 42452 779858 42508 779897
rect 42740 778861 42742 778878
rect 42742 778861 42794 778878
rect 42794 778861 42796 778878
rect 42740 778822 42796 778861
rect 43220 777194 43276 777250
rect 43220 776454 43276 776510
rect 43412 777934 43468 777990
rect 42836 774826 42892 774882
rect 38804 773494 38860 773550
rect 35924 772606 35980 772662
rect 37364 769498 37420 769554
rect 35924 760174 35980 760230
rect 37364 759582 37420 759638
rect 41972 771126 42028 771182
rect 41780 770386 41836 770442
rect 38804 758546 38860 758602
rect 41876 767870 41932 767926
rect 42452 769054 42508 769110
rect 42164 765946 42220 766002
rect 42068 765206 42124 765262
rect 42740 764540 42796 764596
rect 42164 757066 42220 757122
rect 41876 754846 41932 754902
rect 42452 754254 42508 754310
rect 41780 748630 41836 748686
rect 41972 747298 42028 747354
rect 42932 772458 42988 772514
rect 43124 767722 43180 767778
rect 42932 766982 42988 767038
rect 42836 751886 42892 751942
rect 42740 751590 42796 751646
rect 42836 747150 42892 747206
rect 42932 746854 42988 746910
rect 43220 761802 43276 761858
rect 42644 737251 42700 737290
rect 42644 737234 42646 737251
rect 42646 737234 42698 737251
rect 42698 737234 42700 737251
rect 42356 736681 42358 736698
rect 42358 736681 42410 736698
rect 42410 736681 42412 736698
rect 42356 736642 42412 736681
rect 42356 735475 42412 735514
rect 42356 735458 42358 735475
rect 42358 735458 42410 735475
rect 42410 735458 42412 735475
rect 43220 734866 43276 734922
rect 42932 731610 42988 731666
rect 40244 730278 40300 730334
rect 41588 728798 41644 728854
rect 41492 727170 41548 727226
rect 41780 727910 41836 727966
rect 41684 725838 41740 725894
rect 42068 724654 42124 724710
rect 41972 723174 42028 723230
rect 41780 716070 41836 716126
rect 41876 713998 41932 714054
rect 42164 724062 42220 724118
rect 42260 719918 42316 719974
rect 42260 718751 42316 718790
rect 42260 718734 42262 718751
rect 42262 718734 42314 718751
rect 42314 718734 42316 718751
rect 42068 713850 42124 713906
rect 42068 711630 42124 711686
rect 43028 723026 43084 723082
rect 42932 711778 42988 711834
rect 43028 711630 43084 711686
rect 43124 711186 43180 711242
rect 42836 711038 42892 711094
rect 42068 708522 42124 708578
rect 42164 707338 42220 707394
rect 41972 706450 42028 706506
rect 41780 704674 41836 704730
rect 42068 704082 42124 704138
rect 42260 703638 42316 703694
rect 43028 707782 43084 707838
rect 42836 703490 42892 703546
rect 42260 700826 42316 700882
rect 42260 700530 42316 700586
rect 42644 694035 42700 694074
rect 42644 694018 42646 694035
rect 42646 694018 42698 694035
rect 42698 694018 42700 694035
rect 42356 693426 42412 693482
rect 41396 692686 41452 692742
rect 40244 687062 40300 687118
rect 42644 692429 42646 692446
rect 42646 692429 42698 692446
rect 42698 692429 42700 692446
rect 42644 692390 42700 692429
rect 43412 733978 43468 734034
rect 43412 691650 43468 691706
rect 43220 690762 43276 690818
rect 41588 688246 41644 688302
rect 41396 674778 41452 674834
rect 41684 685582 41740 685638
rect 41780 683954 41836 684010
rect 41012 670930 41068 670986
rect 41876 681438 41932 681494
rect 41972 680846 42028 680902
rect 42260 679958 42316 680014
rect 43124 678182 43180 678238
rect 42356 677146 42412 677202
rect 42356 675683 42412 675722
rect 42356 675666 42358 675683
rect 42358 675666 42410 675683
rect 42410 675666 42412 675683
rect 42644 670930 42700 670986
rect 43028 670930 43084 670986
rect 42548 668858 42604 668914
rect 41780 668414 41836 668470
rect 42164 665306 42220 665362
rect 42932 666490 42988 666546
rect 42548 663382 42604 663438
rect 41780 661310 41836 661366
rect 41876 661014 41932 661070
rect 42836 660866 42892 660922
rect 43124 668266 43180 668322
rect 41780 656130 41836 656186
rect 42836 650802 42892 650858
rect 42452 649783 42508 649822
rect 42452 649766 42454 649783
rect 42454 649766 42506 649783
rect 42506 649766 42508 649783
rect 42452 649509 42454 649526
rect 42454 649509 42506 649526
rect 42506 649509 42508 649526
rect 42452 649470 42508 649509
rect 43220 648434 43276 648490
rect 42548 645474 42604 645530
rect 40052 643846 40108 643902
rect 41684 642366 41740 642422
rect 41492 641626 41548 641682
rect 41204 627714 41260 627770
rect 41780 640738 41836 640794
rect 41876 639406 41932 639462
rect 42068 636742 42124 636798
rect 41972 636298 42028 636354
rect 41972 627566 42028 627622
rect 41876 627418 41932 627474
rect 42932 638370 42988 638426
rect 42644 635854 42700 635910
rect 42164 633486 42220 633542
rect 42260 632467 42316 632506
rect 42260 632450 42262 632467
rect 42262 632450 42314 632467
rect 42314 632450 42316 632467
rect 43124 638074 43180 638130
rect 42164 625198 42220 625254
rect 42452 624458 42508 624514
rect 42164 622090 42220 622146
rect 42068 620906 42124 620962
rect 42452 620758 42508 620814
rect 41780 619130 41836 619186
rect 41876 618242 41932 618298
rect 42836 618242 42892 618298
rect 42740 618094 42796 618150
rect 42452 617650 42508 617706
rect 42740 607699 42742 607716
rect 42742 607699 42794 607716
rect 42794 607699 42796 607716
rect 42740 607660 42796 607699
rect 42740 606863 42796 606902
rect 42740 606846 42742 606863
rect 42742 606846 42794 606863
rect 42794 606846 42796 606863
rect 42452 606254 42508 606310
rect 43604 679810 43660 679866
rect 43412 647546 43468 647602
rect 43316 646066 43372 646122
rect 43220 604626 43276 604682
rect 43508 605218 43564 605274
rect 43316 602850 43372 602906
rect 42932 602110 42988 602166
rect 40052 600630 40108 600686
rect 41876 598410 41932 598466
rect 41780 597522 41836 597578
rect 41972 596190 42028 596246
rect 41876 584350 41932 584406
rect 42068 595154 42124 595210
rect 42836 594858 42892 594914
rect 42164 593674 42220 593730
rect 42068 584498 42124 584554
rect 41972 584202 42028 584258
rect 42452 592342 42508 592398
rect 42548 591898 42604 591954
rect 42548 590714 42604 590770
rect 42548 589251 42604 589290
rect 42548 589234 42550 589251
rect 42550 589234 42602 589251
rect 42602 589234 42604 589251
rect 42548 584942 42604 584998
rect 43028 599594 43084 599650
rect 42932 586570 42988 586626
rect 43124 593378 43180 593434
rect 42452 584498 42508 584554
rect 42452 584202 42508 584258
rect 42932 584350 42988 584406
rect 42836 581242 42892 581298
rect 41780 577098 41836 577154
rect 42452 576950 42508 577006
rect 41876 575026 41932 575082
rect 41780 574878 41836 574934
rect 42260 573990 42316 574046
rect 41780 573842 41836 573898
rect 42932 578282 42988 578338
rect 43028 577542 43084 577598
rect 42836 573250 42892 573306
rect 34484 564666 34540 564722
rect 43316 564518 43372 564574
rect 42452 563499 42508 563538
rect 42452 563482 42454 563499
rect 42454 563482 42506 563499
rect 42506 563482 42508 563499
rect 42356 563038 42412 563094
rect 43220 562002 43276 562058
rect 41972 558598 42028 558654
rect 40148 557414 40204 557470
rect 41684 555934 41740 555990
rect 41876 555194 41932 555250
rect 41780 554306 41836 554362
rect 42068 552974 42124 553030
rect 41876 541282 41932 541338
rect 41972 541134 42028 541190
rect 42356 551938 42412 551994
rect 42164 550014 42220 550070
rect 42068 540986 42124 541042
rect 42932 551642 42988 551698
rect 42836 551050 42892 551106
rect 42644 546257 42700 546296
rect 42644 546240 42646 546257
rect 42646 546240 42698 546257
rect 42698 546240 42700 546257
rect 42068 538914 42124 538970
rect 43028 549274 43084 549330
rect 42932 538618 42988 538674
rect 42836 536842 42892 536898
rect 41780 531662 41836 531718
rect 41876 531218 41932 531274
rect 42644 532550 42700 532606
rect 42740 532254 42796 532310
rect 43124 548534 43180 548590
rect 43604 564518 43660 564574
rect 43508 561558 43564 561614
rect 43796 560522 43852 560578
rect 43604 559782 43660 559838
rect 42644 436907 42646 436924
rect 42646 436907 42698 436924
rect 42698 436907 42700 436924
rect 42644 436868 42700 436907
rect 42644 436093 42646 436110
rect 42646 436093 42698 436110
rect 42698 436093 42700 436110
rect 42644 436054 42700 436093
rect 42356 435462 42412 435518
rect 43412 434426 43468 434482
rect 43220 433538 43276 433594
rect 41876 429838 41932 429894
rect 41780 426730 41836 426786
rect 43796 432946 43852 433002
rect 43604 432058 43660 432114
rect 43124 424362 43180 424418
rect 42740 424066 42796 424122
rect 42164 423178 42220 423234
rect 42644 420070 42700 420126
rect 42644 418607 42700 418646
rect 42644 418590 42646 418607
rect 42646 418590 42698 418607
rect 42698 418590 42700 418607
rect 41780 406010 41836 406066
rect 41780 404234 41836 404290
rect 42068 403790 42124 403846
rect 42932 422586 42988 422642
rect 42836 420958 42892 421014
rect 43028 421254 43084 421310
rect 41780 402458 41836 402514
rect 41780 402014 41836 402070
rect 41780 400090 41836 400146
rect 41780 399498 41836 399554
rect 41780 398758 41836 398814
rect 42356 393913 42358 393930
rect 42358 393913 42410 393930
rect 42410 393913 42412 393930
rect 42356 393874 42412 393913
rect 42356 393173 42358 393190
rect 42358 393173 42410 393190
rect 42410 393173 42412 393190
rect 42356 393134 42412 393173
rect 42356 392285 42358 392302
rect 42358 392285 42410 392302
rect 42410 392285 42412 392302
rect 42356 392246 42412 392285
rect 43220 391210 43276 391266
rect 42068 386622 42124 386678
rect 37364 379962 37420 380018
rect 42356 383514 42412 383570
rect 42260 378778 42316 378834
rect 42164 376558 42220 376614
rect 42164 375243 42220 375282
rect 42164 375226 42166 375243
rect 42166 375226 42218 375243
rect 42218 375226 42220 375243
rect 42836 381738 42892 381794
rect 42740 377742 42796 377798
rect 43028 380850 43084 380906
rect 43124 378482 43180 378538
rect 41780 362794 41836 362850
rect 42068 360870 42124 360926
rect 41780 360574 41836 360630
rect 42068 359390 42124 359446
rect 41780 358650 41836 358706
rect 41876 356874 41932 356930
rect 41780 356430 41836 356486
rect 41780 355542 41836 355598
rect 42356 350697 42358 350714
rect 42358 350697 42410 350714
rect 42410 350697 42412 350714
rect 42356 350658 42412 350697
rect 42644 349661 42646 349678
rect 42646 349661 42698 349678
rect 42698 349661 42700 349678
rect 42644 349622 42700 349661
rect 42356 349069 42358 349086
rect 42358 349069 42410 349086
rect 42410 349069 42412 349086
rect 42356 349030 42412 349069
rect 43316 390914 43372 390970
rect 43316 347994 43372 348050
rect 43220 347698 43276 347754
rect 42740 344072 42796 344128
rect 37268 340298 37324 340354
rect 37172 337190 37228 337246
rect 37364 337190 37420 337246
rect 42356 333342 42412 333398
rect 42356 332027 42412 332066
rect 42356 332010 42358 332027
rect 42358 332010 42410 332027
rect 42410 332010 42412 332027
rect 43124 335414 43180 335470
rect 43028 334526 43084 334582
rect 43412 338522 43468 338578
rect 41780 319726 41836 319782
rect 42164 318690 42220 318746
rect 41780 317950 41836 318006
rect 41876 317358 41932 317414
rect 41780 316026 41836 316082
rect 41780 315582 41836 315638
rect 41780 313658 41836 313714
rect 41780 313214 41836 313270
rect 41780 312326 41836 312382
rect 42260 307481 42262 307498
rect 42262 307481 42314 307498
rect 42314 307481 42316 307498
rect 42260 307442 42316 307481
rect 42260 306741 42262 306758
rect 42262 306741 42314 306758
rect 42314 306741 42316 306758
rect 42260 306702 42316 306741
rect 42836 305666 42892 305722
rect 43412 304778 43468 304834
rect 43220 304038 43276 304094
rect 39956 300338 40012 300394
rect 37364 293974 37420 294030
rect 41780 297230 41836 297286
rect 42164 294714 42220 294770
rect 43124 293826 43180 293882
rect 42260 292346 42316 292402
rect 42836 292198 42892 292254
rect 42548 290866 42604 290922
rect 42260 283614 42316 283670
rect 42644 289107 42700 289146
rect 42644 289090 42646 289107
rect 42646 289090 42698 289107
rect 42698 289090 42700 289107
rect 42644 281542 42700 281598
rect 41780 276510 41836 276566
rect 41972 274734 42028 274790
rect 43220 290570 43276 290626
rect 41972 273994 42028 274050
rect 41780 272810 41836 272866
rect 41780 272366 41836 272422
rect 41780 270590 41836 270646
rect 41780 269998 41836 270054
rect 41780 269110 41836 269166
rect 42260 264265 42262 264282
rect 42262 264265 42314 264282
rect 42314 264265 42316 264282
rect 42260 264226 42316 264265
rect 42260 263525 42262 263542
rect 42262 263525 42314 263542
rect 42314 263525 42316 263542
rect 42260 263486 42316 263525
rect 42836 262450 42892 262506
rect 43316 264818 43372 264874
rect 43220 260822 43276 260878
rect 43796 261562 43852 261618
rect 43316 260082 43372 260138
rect 42260 257122 42316 257178
rect 37268 254014 37324 254070
rect 37172 250758 37228 250814
rect 34580 247058 34636 247114
rect 34580 246022 34636 246078
rect 41972 251498 42028 251554
rect 37364 250758 37420 250814
rect 42068 248390 42124 248446
rect 43124 249722 43180 249778
rect 43028 248094 43084 248150
rect 42644 240694 42700 240750
rect 42164 234774 42220 234830
rect 41780 233294 41836 233350
rect 41780 231666 41836 231722
rect 41876 231518 41932 231574
rect 41780 229742 41836 229798
rect 41780 229002 41836 229058
rect 41780 227226 41836 227282
rect 41780 226782 41836 226838
rect 41780 225894 41836 225950
rect 42356 221049 42358 221066
rect 42358 221049 42410 221066
rect 42410 221049 42412 221066
rect 42356 221010 42412 221049
rect 42356 220309 42358 220326
rect 42358 220309 42410 220326
rect 42410 220309 42412 220326
rect 42356 220270 42412 220309
rect 42356 219421 42358 219438
rect 42358 219421 42410 219438
rect 42410 219421 42412 219438
rect 42356 219382 42412 219421
rect 43604 259342 43660 259398
rect 44852 762246 44908 762302
rect 43316 216866 43372 216922
rect 43604 217606 43660 217662
rect 43412 216126 43468 216182
rect 41876 213906 41932 213962
rect 37364 210798 37420 210854
rect 41684 206062 41740 206118
rect 41684 197626 41740 197682
rect 41972 209170 42028 209226
rect 42068 208282 42124 208338
rect 42740 208060 42796 208116
rect 42356 204325 42358 204342
rect 42358 204325 42410 204342
rect 42410 204325 42412 204342
rect 42356 204286 42412 204325
rect 42356 202806 42412 202862
rect 43028 207394 43084 207450
rect 43124 205766 43180 205822
rect 43028 204582 43084 204638
rect 41780 190078 41836 190134
rect 41972 189042 42028 189098
rect 41780 188302 41836 188358
rect 42644 195702 42700 195758
rect 45620 251942 45676 251998
rect 46484 274734 46540 274790
rect 46292 273994 46348 274050
rect 46484 273994 46540 274050
rect 46292 273254 46348 273310
rect 45908 252090 45964 252146
rect 59540 972998 59596 973054
rect 74708 997270 74764 997326
rect 74900 997270 74956 997326
rect 92564 996086 92620 996142
rect 78644 995790 78700 995846
rect 89684 995642 89740 995698
rect 80180 993718 80236 993774
rect 86516 995346 86572 995402
rect 87860 995198 87916 995254
rect 88724 993866 88780 993922
rect 62036 993570 62092 993626
rect 83444 993570 83500 993626
rect 92948 993570 93004 993626
rect 61844 962194 61900 962250
rect 62036 962046 62092 962102
rect 59348 958642 59404 958698
rect 59540 944286 59596 944342
rect 59540 929930 59596 929986
rect 59540 915426 59596 915482
rect 59540 901218 59596 901274
rect 59540 886714 59596 886770
rect 58964 872358 59020 872414
rect 58196 829477 58198 829494
rect 58198 829477 58250 829494
rect 58250 829477 58252 829494
rect 58196 829438 58252 829477
rect 59540 858002 59596 858058
rect 59540 843646 59596 843702
rect 59540 814934 59596 814990
rect 59540 800578 59596 800634
rect 58964 786222 59020 786278
rect 58196 757527 58252 757566
rect 58196 757510 58198 757527
rect 58198 757510 58250 757527
rect 58250 757510 58252 757527
rect 58580 743154 58636 743210
rect 59540 771883 59596 771922
rect 59540 771866 59542 771883
rect 59542 771866 59594 771883
rect 59594 771866 59596 771883
rect 59540 728798 59596 728854
rect 59540 714311 59596 714350
rect 59540 714294 59542 714311
rect 59542 714294 59594 714311
rect 59594 714294 59596 714311
rect 59540 700086 59596 700142
rect 58676 685582 58732 685638
rect 58388 671374 58444 671430
rect 59540 656870 59596 656926
rect 59540 642662 59596 642718
rect 58388 628158 58444 628214
rect 58388 613802 58444 613858
rect 59540 599446 59596 599502
rect 59540 585238 59596 585294
rect 59540 570734 59596 570790
rect 59540 556526 59596 556582
rect 59540 542170 59596 542226
rect 59444 527518 59500 527574
rect 59540 513310 59596 513366
rect 58100 498954 58156 499010
rect 59540 484450 59596 484506
rect 59540 470242 59596 470298
rect 59540 455738 59596 455794
rect 59540 441382 59596 441438
rect 59348 427026 59404 427082
rect 57812 412670 57868 412726
rect 59060 398314 59116 398370
rect 58964 355246 59020 355302
rect 57620 283466 57676 283522
rect 59540 383958 59596 384014
rect 59540 369602 59596 369658
rect 59540 340890 59596 340946
rect 59540 326386 59596 326442
rect 59540 312178 59596 312234
rect 59540 297674 59596 297730
rect 65012 254902 65068 254958
rect 108692 1005449 108694 1005466
rect 108694 1005449 108746 1005466
rect 108746 1005449 108748 1005466
rect 108692 1005410 108748 1005449
rect 115220 1005427 115276 1005466
rect 115220 1005410 115222 1005427
rect 115222 1005410 115274 1005427
rect 115274 1005410 115276 1005427
rect 321044 1005410 321100 1005466
rect 321428 1005410 321484 1005466
rect 325460 1005410 325516 1005466
rect 358676 1005427 358732 1005466
rect 358676 1005410 358678 1005427
rect 358678 1005410 358730 1005427
rect 358730 1005410 358732 1005427
rect 106580 1005279 106636 1005318
rect 106580 1005262 106582 1005279
rect 106582 1005262 106634 1005279
rect 106634 1005262 106636 1005279
rect 109460 1005301 109462 1005318
rect 109462 1005301 109514 1005318
rect 109514 1005301 109516 1005318
rect 109460 1005262 109516 1005301
rect 217268 1005279 217324 1005318
rect 217268 1005262 217270 1005279
rect 217270 1005262 217322 1005279
rect 217322 1005262 217324 1005279
rect 218900 1005279 218956 1005318
rect 218900 1005262 218902 1005279
rect 218902 1005262 218954 1005279
rect 218954 1005262 218956 1005279
rect 223124 1005262 223180 1005318
rect 308756 1005301 308758 1005318
rect 308758 1005301 308810 1005318
rect 308810 1005301 308812 1005318
rect 114164 1005114 114220 1005170
rect 207284 1005153 207286 1005170
rect 207286 1005153 207338 1005170
rect 207338 1005153 207340 1005170
rect 151508 1002615 151564 1002654
rect 151508 1002598 151510 1002615
rect 151510 1002598 151562 1002615
rect 151562 1002598 151564 1002615
rect 101492 995955 101548 995994
rect 101492 995938 101494 995955
rect 101494 995938 101546 995955
rect 101546 995938 101548 995955
rect 103892 995977 103894 995994
rect 103894 995977 103946 995994
rect 103946 995977 103948 995994
rect 103892 995938 103948 995977
rect 106964 995938 107020 995994
rect 113396 995955 113452 995994
rect 113396 995938 113398 995955
rect 113398 995938 113450 995955
rect 113450 995938 113452 995955
rect 95060 995790 95116 995846
rect 99764 995790 99820 995846
rect 105428 995807 105484 995846
rect 105428 995790 105430 995807
rect 105430 995790 105482 995807
rect 105482 995790 105484 995807
rect 94964 995642 95020 995698
rect 98900 995642 98956 995698
rect 99668 995642 99724 995698
rect 103124 995642 103180 995698
rect 98900 995346 98956 995402
rect 100724 995050 100780 995106
rect 113396 995807 113452 995846
rect 113396 995790 113398 995807
rect 113398 995790 113450 995807
rect 113450 995790 113452 995807
rect 123860 995790 123916 995846
rect 134516 995790 134572 995846
rect 115220 995642 115276 995698
rect 108212 995494 108268 995550
rect 115316 995494 115372 995550
rect 106964 993718 107020 993774
rect 115220 995346 115276 995402
rect 129716 994162 129772 994218
rect 136724 995790 136780 995846
rect 137972 995790 138028 995846
rect 137396 995642 137452 995698
rect 143636 995642 143692 995698
rect 152852 1002489 152854 1002506
rect 152854 1002489 152906 1002506
rect 152906 1002489 152908 1002506
rect 152852 1002450 152908 1002489
rect 153620 1002467 153676 1002506
rect 153620 1002450 153622 1002467
rect 153622 1002450 153674 1002467
rect 153674 1002450 153676 1002467
rect 150356 1002341 150358 1002358
rect 150358 1002341 150410 1002358
rect 150410 1002341 150412 1002358
rect 150356 1002302 150412 1002341
rect 144212 995938 144268 995994
rect 144020 995790 144076 995846
rect 136148 994310 136204 994366
rect 134612 994014 134668 994070
rect 160244 1000839 160300 1000878
rect 160244 1000822 160246 1000839
rect 160246 1000822 160298 1000839
rect 160298 1000822 160300 1000839
rect 155156 999507 155212 999546
rect 155156 999490 155158 999507
rect 155158 999490 155210 999507
rect 155210 999490 155212 999507
rect 156884 999381 156886 999398
rect 156886 999381 156938 999398
rect 156938 999381 156940 999398
rect 156884 999342 156940 999381
rect 145268 995938 145324 995994
rect 149108 995938 149164 995994
rect 149492 995938 149548 995994
rect 151988 995955 152044 995994
rect 151988 995938 151990 995955
rect 151990 995938 152042 995955
rect 152042 995938 152044 995955
rect 140372 993718 140428 993774
rect 159476 995938 159532 995994
rect 158612 995790 158668 995846
rect 146804 995659 146860 995698
rect 146804 995642 146806 995659
rect 146806 995642 146858 995659
rect 146858 995642 146860 995659
rect 158324 995642 158380 995698
rect 146804 995494 146860 995550
rect 158324 994162 158380 994218
rect 164084 996103 164140 996142
rect 164084 996086 164086 996103
rect 164086 996086 164138 996103
rect 164138 996086 164140 996103
rect 164180 995977 164182 995994
rect 164182 995977 164234 995994
rect 164234 995977 164236 995994
rect 164180 995938 164236 995977
rect 165620 995807 165676 995846
rect 165620 995790 165622 995807
rect 165622 995790 165674 995807
rect 165674 995790 165676 995807
rect 166196 995790 166252 995846
rect 178484 995790 178540 995846
rect 185204 995790 185260 995846
rect 162932 995642 162988 995698
rect 162644 995494 162700 995550
rect 170228 995642 170284 995698
rect 185108 995494 185164 995550
rect 187604 995790 187660 995846
rect 192500 995790 192556 995846
rect 189428 995642 189484 995698
rect 195380 995938 195436 995994
rect 195284 995790 195340 995846
rect 185396 994162 185452 994218
rect 190580 995494 190636 995550
rect 185972 994014 186028 994070
rect 181460 985469 181462 985486
rect 181462 985469 181514 985486
rect 181514 985469 181516 985486
rect 181460 985430 181516 985469
rect 187316 985430 187372 985486
rect 207284 1005114 207340 1005153
rect 221876 1005114 221932 1005170
rect 211700 1003673 211702 1003690
rect 211702 1003673 211754 1003690
rect 211754 1003673 211756 1003690
rect 211700 1003634 211756 1003673
rect 208148 1000861 208150 1000878
rect 208150 1000861 208202 1000878
rect 208202 1000861 208204 1000878
rect 208148 1000822 208204 1000861
rect 209396 997901 209398 997918
rect 209398 997901 209450 997918
rect 209450 997901 209452 997918
rect 209396 997862 209452 997901
rect 213332 996125 213334 996142
rect 213334 996125 213386 996142
rect 213386 996125 213388 996142
rect 213332 996086 213388 996125
rect 215636 996103 215692 996142
rect 215636 996086 215638 996103
rect 215638 996086 215690 996103
rect 215690 996086 215692 996103
rect 200276 995955 200332 995994
rect 200276 995938 200278 995955
rect 200278 995938 200330 995955
rect 200330 995938 200332 995955
rect 200948 995955 201004 995994
rect 200948 995938 200950 995955
rect 200950 995938 201002 995955
rect 201002 995938 201004 995955
rect 204212 995938 204268 995994
rect 206612 995938 206668 995994
rect 202868 995807 202924 995846
rect 202868 995790 202870 995807
rect 202870 995790 202922 995807
rect 202922 995790 202924 995807
rect 203348 995790 203404 995846
rect 216788 995955 216844 995994
rect 216788 995938 216790 995955
rect 216790 995938 216842 995955
rect 216842 995938 216844 995955
rect 203348 995346 203404 995402
rect 212660 995346 212716 995402
rect 201524 995198 201580 995254
rect 210164 995198 210220 995254
rect 211028 995198 211084 995254
rect 218900 995642 218956 995698
rect 214388 995346 214444 995402
rect 238868 995790 238924 995846
rect 239540 995790 239596 995846
rect 240212 995642 240268 995698
rect 231476 994310 231532 994366
rect 227540 994162 227596 994218
rect 234356 994458 234412 994514
rect 240788 995494 240844 995550
rect 241844 995346 241900 995402
rect 237428 994014 237484 994070
rect 243572 994606 243628 994662
rect 243188 994014 243244 994070
rect 258836 999507 258892 999546
rect 258836 999490 258838 999507
rect 258838 999490 258890 999507
rect 258890 999490 258892 999507
rect 260756 999529 260758 999546
rect 260758 999529 260810 999546
rect 260810 999529 260812 999546
rect 260756 999490 260812 999529
rect 246644 995938 246700 995994
rect 247604 995938 247660 995994
rect 259604 999381 259606 999398
rect 259606 999381 259658 999398
rect 259658 999381 259660 999398
rect 259604 999342 259660 999381
rect 263924 996547 263980 996586
rect 263924 996530 263926 996547
rect 263926 996530 263978 996547
rect 263978 996530 263980 996547
rect 250484 995807 250540 995846
rect 250484 995790 250486 995807
rect 250486 995790 250538 995807
rect 250538 995790 250540 995807
rect 254036 995807 254092 995846
rect 254036 995790 254038 995807
rect 254038 995790 254090 995807
rect 254090 995790 254092 995807
rect 254900 995829 254902 995846
rect 254902 995829 254954 995846
rect 254954 995829 254956 995846
rect 254900 995790 254956 995829
rect 255668 995790 255724 995846
rect 257300 995829 257302 995846
rect 257302 995829 257354 995846
rect 257354 995829 257356 995846
rect 257300 995790 257356 995829
rect 250388 995681 250390 995698
rect 250390 995681 250442 995698
rect 250442 995681 250444 995698
rect 250388 995642 250444 995681
rect 250484 995050 250540 995106
rect 265076 996125 265078 996142
rect 265078 996125 265130 996142
rect 265130 996125 265132 996142
rect 265076 996086 265132 996125
rect 266996 996103 267052 996142
rect 266996 996086 266998 996103
rect 266998 996086 267050 996103
rect 267050 996086 267052 996103
rect 266900 995938 266956 995994
rect 262676 995790 262732 995846
rect 268532 995807 268588 995846
rect 268532 995790 268534 995807
rect 268534 995790 268586 995807
rect 268586 995790 268588 995807
rect 273620 995790 273676 995846
rect 265748 995642 265804 995698
rect 268052 995642 268108 995698
rect 262676 994606 262732 994662
rect 292532 995790 292588 995846
rect 295412 995642 295468 995698
rect 308756 1005262 308812 1005301
rect 309620 1005279 309676 1005318
rect 309620 1005262 309622 1005279
rect 309622 1005262 309674 1005279
rect 309674 1005262 309676 1005279
rect 299444 995829 299446 995846
rect 299446 995829 299498 995846
rect 299498 995829 299500 995846
rect 299444 995790 299500 995829
rect 298196 995642 298252 995698
rect 298484 995642 298540 995698
rect 286772 995494 286828 995550
rect 286292 994606 286348 994662
rect 284372 994458 284428 994514
rect 279284 993609 279286 993626
rect 279286 993609 279338 993626
rect 279338 993609 279340 993626
rect 279284 993570 279340 993609
rect 293588 995346 293644 995402
rect 290324 994754 290380 994810
rect 288980 994162 289036 994218
rect 294548 994162 294604 994218
rect 288404 993570 288460 993626
rect 431636 1005427 431692 1005466
rect 431636 1005410 431638 1005427
rect 431638 1005410 431690 1005427
rect 431690 1005410 431692 1005427
rect 433268 1005449 433270 1005466
rect 433270 1005449 433322 1005466
rect 433322 1005449 433324 1005466
rect 433268 1005410 433324 1005449
rect 365012 1005301 365014 1005318
rect 365014 1005301 365066 1005318
rect 365066 1005301 365068 1005318
rect 365012 1005262 365068 1005301
rect 314228 1005153 314230 1005170
rect 314230 1005153 314282 1005170
rect 314282 1005153 314284 1005170
rect 314228 1005114 314284 1005153
rect 358004 1005153 358006 1005170
rect 358006 1005153 358058 1005170
rect 358058 1005153 358060 1005170
rect 311252 999381 311254 999398
rect 311254 999381 311306 999398
rect 311306 999381 311308 999398
rect 311252 999342 311308 999381
rect 318452 997753 318454 997770
rect 318454 997753 318506 997770
rect 318506 997753 318508 997770
rect 318452 997714 318508 997753
rect 316340 996125 316342 996142
rect 316342 996125 316394 996142
rect 316394 996125 316396 996142
rect 316340 996086 316396 996125
rect 318644 996103 318700 996142
rect 318644 996086 318646 996103
rect 318646 996086 318698 996103
rect 318698 996086 318700 996103
rect 305684 995938 305740 995994
rect 313844 995938 313900 995994
rect 304724 995829 304726 995846
rect 304726 995829 304778 995846
rect 304778 995829 304780 995846
rect 304724 995790 304780 995829
rect 307316 995790 307372 995846
rect 310292 995807 310348 995846
rect 310292 995790 310294 995807
rect 310294 995790 310346 995807
rect 310346 995790 310348 995807
rect 299540 995494 299596 995550
rect 302324 995533 302326 995550
rect 302326 995533 302378 995550
rect 302378 995533 302380 995550
rect 302324 995494 302380 995533
rect 309236 995642 309292 995698
rect 313364 995642 313420 995698
rect 309236 994754 309292 994810
rect 313364 994458 313420 994514
rect 317492 995790 317548 995846
rect 323924 995642 323980 995698
rect 326804 995938 326860 995994
rect 358004 1005114 358060 1005153
rect 356756 1003947 356812 1003986
rect 356756 1003930 356758 1003947
rect 356758 1003930 356810 1003947
rect 356810 1003930 356812 1003947
rect 355988 1003799 356044 1003838
rect 355988 1003782 355990 1003799
rect 355990 1003782 356042 1003799
rect 356042 1003782 356044 1003799
rect 359060 1003821 359062 1003838
rect 359062 1003821 359114 1003838
rect 359114 1003821 359116 1003838
rect 359060 1003782 359116 1003821
rect 359924 1003673 359926 1003690
rect 359926 1003673 359978 1003690
rect 359978 1003673 359980 1003690
rect 359924 1003634 359980 1003673
rect 361556 1000839 361612 1000878
rect 361556 1000822 361558 1000839
rect 361558 1000822 361610 1000839
rect 361610 1000822 361612 1000839
rect 367892 997901 367894 997918
rect 367894 997901 367946 997918
rect 367946 997901 367948 997918
rect 367892 997862 367948 997901
rect 369044 997753 369046 997770
rect 369046 997753 369098 997770
rect 369098 997753 369100 997770
rect 369044 997714 369100 997753
rect 367124 996103 367180 996142
rect 367124 996086 367126 996103
rect 367126 996086 367178 996103
rect 367178 996086 367180 996103
rect 362324 995938 362380 995994
rect 370196 995955 370252 995994
rect 370196 995938 370198 995955
rect 370198 995938 370250 995955
rect 370250 995938 370252 995955
rect 350132 995790 350188 995846
rect 360980 995807 361036 995846
rect 360980 995790 360982 995807
rect 360982 995790 361034 995807
rect 361034 995790 361036 995807
rect 365876 995790 365932 995846
rect 377492 995938 377548 995994
rect 368852 995642 368908 995698
rect 374420 995642 374476 995698
rect 365780 994458 365836 994514
rect 377300 995790 377356 995846
rect 380276 996086 380332 996142
rect 380180 995790 380236 995846
rect 381428 995642 381484 995698
rect 424532 1005279 424588 1005318
rect 424532 1005262 424534 1005279
rect 424534 1005262 424586 1005279
rect 424586 1005262 424588 1005279
rect 425300 1005301 425302 1005318
rect 425302 1005301 425354 1005318
rect 425354 1005301 425356 1005318
rect 425300 1005262 425356 1005301
rect 434804 1005301 434806 1005318
rect 434806 1005301 434858 1005318
rect 434858 1005301 434860 1005318
rect 426068 1005153 426070 1005170
rect 426070 1005153 426122 1005170
rect 426122 1005153 426124 1005170
rect 426068 1005114 426124 1005153
rect 434804 1005262 434860 1005301
rect 435572 1005131 435628 1005170
rect 435572 1005114 435574 1005131
rect 435574 1005114 435626 1005131
rect 435626 1005114 435628 1005131
rect 423380 1003799 423436 1003838
rect 423380 1003782 423382 1003799
rect 423382 1003782 423434 1003799
rect 423434 1003782 423436 1003799
rect 428084 1003821 428086 1003838
rect 428086 1003821 428138 1003838
rect 428138 1003821 428140 1003838
rect 428084 1003782 428140 1003821
rect 426452 1003673 426454 1003690
rect 426454 1003673 426506 1003690
rect 426506 1003673 426508 1003690
rect 426452 1003634 426508 1003673
rect 434036 1001135 434092 1001174
rect 434036 1001118 434038 1001135
rect 434038 1001118 434090 1001135
rect 434090 1001118 434092 1001135
rect 430868 1000987 430924 1001026
rect 430868 1000970 430870 1000987
rect 430870 1000970 430922 1000987
rect 430922 1000970 430924 1000987
rect 432500 1001009 432502 1001026
rect 432502 1001009 432554 1001026
rect 432554 1001009 432556 1001026
rect 432500 1000970 432556 1001009
rect 427316 1000839 427372 1000878
rect 427316 1000822 427318 1000839
rect 427318 1000822 427370 1000839
rect 427370 1000822 427372 1000839
rect 428948 1000861 428950 1000878
rect 428950 1000861 429002 1000878
rect 429002 1000861 429004 1000878
rect 428948 1000822 429004 1000861
rect 436436 996125 436438 996142
rect 436438 996125 436490 996142
rect 436490 996125 436492 996142
rect 436436 996086 436492 996125
rect 438740 1005262 438796 1005318
rect 439700 1005262 439756 1005318
rect 444884 1005262 444940 1005318
rect 429716 995938 429772 995994
rect 436436 995977 436438 995994
rect 436438 995977 436490 995994
rect 436490 995977 436492 995994
rect 436436 995938 436492 995977
rect 388820 995790 388876 995846
rect 396692 995790 396748 995846
rect 393044 995642 393100 995698
rect 410324 995642 410380 995698
rect 385844 995494 385900 995550
rect 387476 995346 387532 995402
rect 382004 995050 382060 995106
rect 379028 994902 379084 994958
rect 388340 994458 388396 994514
rect 392084 995198 392140 995254
rect 392660 995050 392716 995106
rect 394868 995494 394924 995550
rect 393716 994902 393772 994958
rect 391124 994458 391180 994514
rect 396308 994310 396364 994366
rect 390164 993570 390220 993626
rect 390164 992090 390220 992146
rect 440660 995642 440716 995698
rect 445076 1005114 445132 1005170
rect 504596 1005449 504598 1005466
rect 504598 1005449 504650 1005466
rect 504650 1005449 504652 1005466
rect 466484 995790 466540 995846
rect 469556 994606 469612 994662
rect 504596 1005410 504652 1005449
rect 502292 1005279 502348 1005318
rect 502292 1005262 502294 1005279
rect 502294 1005262 502346 1005279
rect 502346 1005262 502348 1005279
rect 498356 1005114 498412 1005170
rect 498740 1005114 498796 1005170
rect 508628 1005153 508630 1005170
rect 508630 1005153 508682 1005170
rect 508682 1005153 508684 1005170
rect 508628 1005114 508684 1005153
rect 554516 1005279 554572 1005318
rect 554516 1005262 554518 1005279
rect 554518 1005262 554570 1005279
rect 554570 1005262 554572 1005279
rect 501140 1003821 501142 1003838
rect 501142 1003821 501194 1003838
rect 501194 1003821 501196 1003838
rect 501140 1003782 501196 1003821
rect 500372 1003673 500374 1003690
rect 500374 1003673 500426 1003690
rect 500426 1003673 500428 1003690
rect 500372 1003634 500428 1003673
rect 502772 1002489 502774 1002506
rect 502774 1002489 502826 1002506
rect 502826 1002489 502828 1002506
rect 502772 1002450 502828 1002489
rect 503444 1002467 503500 1002506
rect 503444 1002450 503446 1002467
rect 503446 1002450 503498 1002467
rect 503498 1002450 503500 1002467
rect 472052 995938 472108 995994
rect 488852 999342 488908 999398
rect 477044 995790 477100 995846
rect 481460 995790 481516 995846
rect 469460 993587 469516 993626
rect 480116 995642 480172 995698
rect 488852 995642 488908 995698
rect 479828 994458 479884 994514
rect 485972 994606 486028 994662
rect 505076 1002319 505132 1002358
rect 505076 1002302 505078 1002319
rect 505078 1002302 505130 1002319
rect 505130 1002302 505132 1002319
rect 510932 1000987 510988 1001026
rect 510932 1000970 510934 1000987
rect 510934 1000970 510986 1000987
rect 510986 1000970 510988 1000987
rect 509300 1000839 509356 1000878
rect 509300 1000822 509302 1000839
rect 509302 1000822 509354 1000839
rect 509354 1000822 509356 1000839
rect 497588 999342 497644 999398
rect 506324 999359 506380 999398
rect 506324 999342 506326 999359
rect 506326 999342 506378 999359
rect 506378 999342 506380 999359
rect 507860 996547 507916 996586
rect 507860 996530 507862 996547
rect 507862 996530 507914 996547
rect 507914 996530 507916 996547
rect 510260 996569 510262 996586
rect 510262 996569 510314 996586
rect 510314 996569 510316 996586
rect 510260 996530 510316 996569
rect 511124 996103 511180 996142
rect 511124 996086 511126 996103
rect 511126 996086 511178 996103
rect 511178 996086 511180 996103
rect 513428 996125 513430 996142
rect 513430 996125 513482 996142
rect 513482 996125 513484 996142
rect 513428 996086 513484 996125
rect 511892 995977 511894 995994
rect 511894 995977 511946 995994
rect 511946 995977 511948 995994
rect 511892 995938 511948 995977
rect 513428 995977 513430 995994
rect 513430 995977 513482 995994
rect 513482 995977 513484 995994
rect 513428 995938 513484 995977
rect 506612 995346 506668 995402
rect 515540 994606 515596 994662
rect 516692 1000987 516748 1001026
rect 516692 1000970 516694 1000987
rect 516694 1000970 516746 1000987
rect 516746 1000970 516748 1000987
rect 516692 1000839 516748 1000878
rect 516692 1000822 516694 1000839
rect 516694 1000822 516746 1000839
rect 516746 1000822 516748 1000839
rect 516788 1000674 516844 1000730
rect 516692 999507 516748 999546
rect 516692 999490 516694 999507
rect 516694 999490 516746 999507
rect 516746 999490 516748 999507
rect 516692 999359 516748 999398
rect 516692 999342 516694 999359
rect 516694 999342 516746 999359
rect 516746 999342 516748 999359
rect 518420 995642 518476 995698
rect 469460 993570 469462 993587
rect 469462 993570 469514 993587
rect 469514 993570 469516 993587
rect 518516 995494 518572 995550
rect 519476 995790 519532 995846
rect 521396 999638 521452 999694
rect 523604 1000970 523660 1001026
rect 523508 1000674 523564 1000730
rect 523412 999934 523468 999990
rect 521492 999490 521548 999546
rect 521012 995494 521068 995550
rect 521204 995642 521260 995698
rect 521396 995938 521452 995994
rect 523700 1000822 523756 1000878
rect 523892 999638 523948 999694
rect 523796 999342 523852 999398
rect 547124 1005114 547180 1005170
rect 553748 1005153 553750 1005170
rect 553750 1005153 553802 1005170
rect 553802 1005153 553804 1005170
rect 553748 1005114 553804 1005153
rect 562484 1005153 562486 1005170
rect 562486 1005153 562538 1005170
rect 562538 1005153 562540 1005170
rect 562484 1005114 562540 1005153
rect 524084 999490 524140 999546
rect 532820 995790 532876 995846
rect 532244 995642 532300 995698
rect 523412 995346 523468 995402
rect 530900 995346 530956 995402
rect 534068 995494 534124 995550
rect 533684 994606 533740 994662
rect 531188 994458 531244 994514
rect 551732 1003821 551734 1003838
rect 551734 1003821 551786 1003838
rect 551786 1003821 551788 1003838
rect 551732 1003782 551788 1003821
rect 556532 1003799 556588 1003838
rect 556532 1003782 556534 1003799
rect 556534 1003782 556586 1003799
rect 556586 1003782 556588 1003799
rect 552596 1003673 552598 1003690
rect 552598 1003673 552650 1003690
rect 552650 1003673 552652 1003690
rect 552596 1003634 552652 1003673
rect 559124 1002489 559126 1002506
rect 559126 1002489 559178 1002506
rect 559178 1002489 559180 1002506
rect 559124 1002450 559180 1002489
rect 559892 1002467 559948 1002506
rect 559892 1002450 559894 1002467
rect 559894 1002450 559946 1002467
rect 559946 1002450 559948 1002467
rect 560564 1002341 560566 1002358
rect 560566 1002341 560618 1002358
rect 560618 1002341 560620 1002358
rect 560564 1002302 560620 1002341
rect 561524 1002319 561580 1002358
rect 561524 1002302 561526 1002319
rect 561526 1002302 561578 1002319
rect 561578 1002302 561580 1002319
rect 564788 1002341 564790 1002358
rect 564790 1002341 564842 1002358
rect 564842 1002341 564844 1002358
rect 555188 997901 555190 997918
rect 555190 997901 555242 997918
rect 555242 997901 555244 997918
rect 555188 997862 555244 997901
rect 557300 997879 557356 997918
rect 557300 997862 557302 997879
rect 557302 997862 557354 997879
rect 557354 997862 557356 997879
rect 556148 997753 556150 997770
rect 556150 997753 556202 997770
rect 556202 997753 556204 997770
rect 556148 997714 556204 997753
rect 564788 1002302 564844 1002341
rect 564788 995977 564790 995994
rect 564790 995977 564842 995994
rect 564842 995977 564844 995994
rect 564788 995938 564844 995977
rect 563732 995807 563788 995846
rect 563732 995790 563734 995807
rect 563734 995790 563786 995807
rect 563786 995790 563788 995807
rect 562772 995659 562828 995698
rect 562772 995642 562774 995659
rect 562774 995642 562826 995659
rect 562826 995642 562828 995659
rect 557972 995346 558028 995402
rect 570260 995642 570316 995698
rect 570452 995494 570508 995550
rect 570356 994754 570412 994810
rect 570836 994902 570892 994958
rect 573140 995790 573196 995846
rect 571028 994606 571084 994662
rect 576020 993866 576076 993922
rect 629972 994902 630028 994958
rect 630740 994458 630796 994514
rect 632756 994458 632812 994514
rect 633620 993718 633676 993774
rect 634292 994754 634348 994810
rect 638516 994310 638572 994366
rect 639188 994606 639244 994662
rect 640724 994162 640780 994218
rect 650036 994014 650092 994070
rect 66164 273271 66220 273310
rect 66164 273254 66166 273271
rect 66166 273254 66218 273271
rect 66218 273254 66220 273271
rect 66932 269258 66988 269314
rect 65876 259046 65932 259102
rect 65108 254754 65164 254810
rect 69332 269702 69388 269758
rect 71732 269406 71788 269462
rect 72980 263486 73036 263542
rect 70580 258898 70636 258954
rect 74132 258750 74188 258806
rect 77684 269850 77740 269906
rect 76532 258602 76588 258658
rect 80564 273271 80620 273310
rect 80564 273254 80566 273271
rect 80566 273254 80618 273271
rect 80618 273254 80620 273271
rect 81332 269554 81388 269610
rect 83636 269998 83692 270054
rect 78932 258454 78988 258510
rect 80660 255681 80662 255698
rect 80662 255681 80714 255698
rect 80714 255681 80716 255698
rect 80660 255642 80716 255681
rect 86228 273254 86284 273310
rect 86420 273254 86476 273310
rect 86036 258306 86092 258362
rect 87188 258010 87244 258066
rect 90740 270146 90796 270202
rect 93140 270294 93196 270350
rect 95540 270442 95596 270498
rect 91988 258158 92044 258214
rect 88436 257714 88492 257770
rect 86708 255659 86764 255698
rect 86708 255642 86710 255659
rect 86710 255642 86762 255659
rect 86762 255642 86764 255659
rect 100916 273419 100972 273458
rect 100916 273402 100918 273419
rect 100918 273402 100970 273419
rect 100970 273402 100972 273419
rect 100244 270590 100300 270646
rect 96788 257862 96844 257918
rect 107444 269110 107500 269166
rect 116948 263782 117004 263838
rect 113396 263634 113452 263690
rect 120788 273419 120844 273458
rect 120788 273402 120790 273419
rect 120790 273402 120842 273419
rect 120842 273402 120844 273419
rect 120500 263930 120556 263986
rect 138164 255790 138220 255846
rect 118100 255681 118102 255698
rect 118102 255681 118154 255698
rect 118154 255681 118156 255698
rect 118100 255642 118156 255681
rect 144020 248094 144076 248150
rect 144116 246318 144172 246374
rect 144020 245282 144076 245338
rect 144020 242766 144076 242822
rect 144020 239083 144076 239122
rect 144020 239066 144022 239083
rect 144022 239066 144074 239083
rect 144074 239066 144076 239083
rect 144020 237882 144076 237938
rect 144116 234330 144172 234386
rect 144020 233442 144076 233498
rect 144020 231222 144076 231278
rect 144116 229446 144172 229502
rect 144020 228854 144076 228910
rect 145460 249278 145516 249334
rect 145748 242026 145804 242082
rect 145364 236106 145420 236162
rect 144020 225006 144076 225062
rect 144020 223970 144076 224026
rect 144116 221306 144172 221362
rect 144020 219974 144076 220030
rect 144020 218067 144076 218106
rect 144020 218050 144022 218067
rect 144022 218050 144074 218067
rect 144074 218050 144076 218067
rect 144020 214350 144076 214406
rect 144020 210798 144076 210854
rect 144020 209022 144076 209078
rect 144980 203398 145036 203454
rect 144980 200586 145036 200642
rect 144404 199402 144460 199458
rect 145268 197626 145324 197682
rect 144980 196146 145036 196202
rect 144596 193926 144652 193982
rect 144308 192150 144364 192206
rect 144884 190966 144940 191022
rect 41780 185934 41836 185990
rect 41780 184158 41836 184214
rect 41780 183566 41836 183622
rect 41780 182826 41836 182882
rect 144692 182678 144748 182734
rect 145172 187414 145228 187470
rect 145076 184306 145132 184362
rect 144884 180754 144940 180810
rect 144020 179126 144076 179182
rect 144692 177794 144748 177850
rect 42740 177054 42796 177110
rect 144500 177054 144556 177110
rect 144404 172318 144460 172374
rect 144020 164622 144076 164678
rect 144308 163882 144364 163938
rect 144212 162106 144268 162162
rect 144308 160330 144364 160386
rect 144116 158554 144172 158610
rect 144308 156186 144364 156242
rect 144212 155446 144268 155502
rect 144308 153670 144364 153726
rect 144308 150710 144364 150766
rect 144212 148934 144268 148990
rect 144308 147750 144364 147806
rect 144308 145234 144364 145290
rect 144308 143458 144364 143514
rect 144308 140498 144364 140554
rect 144212 139314 144268 139370
rect 144596 169950 144652 170006
rect 144500 157370 144556 157426
rect 144500 153078 144556 153134
rect 144500 151894 144556 151950
rect 144500 147010 144556 147066
rect 144500 144346 144556 144402
rect 144500 142291 144556 142330
rect 144500 142274 144502 142291
rect 144502 142274 144554 142291
rect 144554 142274 144556 142291
rect 144500 138574 144556 138630
rect 144212 136946 144268 137002
rect 144116 135910 144172 135966
rect 144116 135022 144172 135078
rect 144020 132671 144076 132710
rect 144020 132654 144022 132671
rect 144022 132654 144074 132671
rect 144074 132654 144076 132671
rect 144212 133838 144268 133894
rect 144116 130878 144172 130934
rect 144212 130138 144268 130194
rect 144116 128510 144172 128566
rect 144212 127326 144268 127382
rect 144020 126586 144076 126642
rect 144212 125402 144268 125458
rect 144116 124218 144172 124274
rect 144212 121850 144268 121906
rect 144116 120074 144172 120130
rect 144020 118890 144076 118946
rect 144212 118150 144268 118206
rect 144116 116966 144172 117022
rect 144212 115486 144268 115542
rect 144116 114154 144172 114210
rect 144212 113414 144268 113470
rect 144020 111638 144076 111694
rect 144116 110454 144172 110510
rect 144212 109714 144268 109770
rect 144212 106902 144268 106958
rect 144020 105718 144076 105774
rect 144116 104978 144172 105034
rect 144212 103811 144268 103850
rect 144212 103794 144214 103811
rect 144214 103794 144266 103811
rect 144266 103794 144268 103811
rect 144212 102018 144268 102074
rect 144212 100094 144268 100150
rect 144116 97282 144172 97338
rect 144020 95358 144076 95414
rect 143924 92250 143980 92306
rect 144212 96542 144268 96598
rect 144212 93599 144268 93638
rect 144212 93582 144214 93599
rect 144214 93582 144266 93599
rect 144266 93582 144268 93599
rect 144116 91806 144172 91862
rect 144212 90639 144268 90678
rect 144212 90622 144214 90639
rect 144214 90622 144266 90639
rect 144266 90622 144268 90639
rect 144212 89307 144268 89346
rect 144212 89290 144214 89307
rect 144214 89290 144266 89307
rect 144266 89290 144268 89307
rect 144116 88106 144172 88162
rect 144212 86922 144268 86978
rect 144116 85146 144172 85202
rect 144116 83370 144172 83426
rect 144116 79670 144172 79726
rect 144212 78486 144268 78542
rect 144212 77319 144268 77358
rect 144212 77302 144214 77319
rect 144214 77302 144266 77319
rect 144266 77302 144268 77319
rect 144212 75822 144268 75878
rect 143924 73767 143980 73806
rect 143924 73750 143926 73767
rect 143926 73750 143978 73767
rect 143978 73750 143980 73767
rect 143924 72122 143980 72178
rect 143828 68274 143884 68330
rect 143924 67090 143980 67146
rect 143924 66811 143980 66850
rect 143924 66794 143926 66811
rect 143926 66794 143978 66811
rect 143978 66794 143980 66811
rect 143924 64722 143980 64778
rect 143924 54658 143980 54714
rect 144212 54658 144268 54714
rect 144788 173502 144844 173558
rect 144980 175870 145036 175926
rect 144980 174242 145036 174298
rect 144980 170542 145036 170598
rect 144980 168618 145036 168674
rect 144980 167138 145036 167194
rect 144980 165806 145036 165862
rect 144980 161514 145036 161570
rect 145460 232406 145516 232462
rect 145556 227670 145612 227726
rect 145652 225894 145708 225950
rect 145748 222786 145804 222842
rect 145844 219234 145900 219290
rect 145940 216274 145996 216330
rect 146516 215534 146572 215590
rect 146036 213314 146092 213370
rect 146132 211538 146188 211594
rect 146228 207838 146284 207894
rect 146804 207098 146860 207154
rect 146324 206062 146380 206118
rect 146804 204878 146860 204934
rect 146420 202362 146476 202418
rect 146708 198662 146764 198718
rect 146516 190374 146572 190430
rect 146612 186230 146668 186286
rect 146804 194666 146860 194722
rect 146804 189190 146860 189246
rect 146804 185490 146860 185546
rect 146804 181938 146860 181994
rect 147476 122442 147532 122498
rect 147380 100834 147436 100890
rect 147284 98466 147340 98522
rect 146900 83831 146956 83870
rect 146900 83814 146902 83831
rect 146902 83814 146954 83831
rect 146954 83814 146956 83831
rect 146996 82203 147052 82242
rect 146996 82186 146998 82203
rect 146998 82186 147050 82203
rect 147050 82186 147052 82203
rect 146900 81002 146956 81058
rect 146900 74951 146956 74990
rect 146900 74934 146902 74951
rect 146902 74934 146954 74951
rect 146954 74934 146956 74951
rect 146996 71234 147052 71290
rect 146900 70067 146956 70106
rect 146900 70050 146902 70067
rect 146902 70050 146954 70067
rect 146954 70050 146956 70067
rect 146900 64147 146956 64186
rect 146900 64130 146902 64147
rect 146902 64130 146954 64147
rect 146954 64130 146956 64147
rect 147572 108530 147628 108586
rect 146996 62206 147052 62262
rect 146900 61170 146956 61226
rect 148244 48590 148300 48646
rect 148052 47702 148108 47758
rect 148436 48442 148492 48498
rect 148628 48294 148684 48350
rect 149204 48146 149260 48202
rect 148820 47554 148876 47610
rect 149396 47998 149452 48054
rect 149588 47850 149644 47906
rect 156884 228558 156940 228614
rect 181556 273402 181612 273458
rect 181556 273106 181612 273162
rect 197876 264670 197932 264726
rect 198740 260691 198796 260730
rect 198740 260674 198742 260691
rect 198742 260674 198794 260691
rect 198794 260674 198796 260691
rect 199796 222046 199852 222102
rect 199700 221750 199756 221806
rect 198740 219086 198796 219142
rect 198740 218642 198796 218698
rect 198836 217458 198892 217514
rect 199028 218050 199084 218106
rect 198932 217310 198988 217366
rect 198740 216422 198796 216478
rect 198740 215847 198796 215886
rect 198740 215830 198742 215847
rect 198742 215830 198794 215847
rect 198794 215830 198796 215847
rect 198836 215721 198838 215738
rect 198838 215721 198890 215738
rect 198890 215721 198892 215738
rect 198836 215682 198892 215721
rect 198740 214794 198796 214850
rect 198836 214202 198892 214258
rect 198932 214054 198988 214110
rect 199028 213166 199084 213222
rect 198740 212574 198796 212630
rect 198836 93434 198892 93490
rect 198740 92398 198796 92454
rect 198932 93286 198988 93342
rect 198740 91806 198796 91862
rect 198836 91066 198892 91122
rect 199124 91658 199180 91714
rect 199028 90178 199084 90234
rect 198932 90030 198988 90086
rect 198740 89011 198796 89050
rect 198740 88994 198742 89011
rect 198742 88994 198794 89011
rect 198794 88994 198796 89011
rect 198932 88550 198988 88606
rect 198836 87810 198892 87866
rect 199220 88402 199276 88458
rect 199028 86922 199084 86978
rect 198836 86182 198892 86238
rect 198740 86073 198742 86090
rect 198742 86073 198794 86090
rect 198794 86073 198796 86090
rect 198740 86034 198796 86073
rect 198932 85294 198988 85350
rect 199124 84998 199180 85054
rect 199028 84554 199084 84610
rect 199220 83666 199276 83722
rect 198740 83239 198796 83278
rect 198740 83222 198742 83239
rect 198742 83222 198794 83239
rect 198794 83222 198796 83239
rect 198836 81742 198892 81798
rect 199508 82038 199564 82094
rect 198932 81298 198988 81354
rect 198740 80427 198796 80466
rect 198740 80410 198742 80427
rect 198742 80410 198794 80427
rect 198794 80410 198796 80427
rect 198740 79818 198796 79874
rect 198836 79670 198892 79726
rect 198932 78782 198988 78838
rect 199028 78190 199084 78246
rect 198740 77637 198742 77654
rect 198742 77637 198794 77654
rect 198794 77637 198796 77654
rect 198740 77598 198796 77637
rect 198740 77154 198796 77210
rect 198932 76562 198988 76618
rect 198836 76414 198892 76470
rect 199028 75526 199084 75582
rect 199124 74934 199180 74990
rect 198740 74490 198796 74546
rect 198932 73898 198988 73954
rect 198836 73306 198892 73362
rect 199028 73158 199084 73214
rect 199124 72270 199180 72326
rect 198740 71695 198796 71734
rect 198740 71678 198742 71695
rect 198742 71678 198794 71695
rect 198794 71678 198796 71695
rect 198836 70050 198892 70106
rect 199604 70938 199660 70994
rect 198932 69902 198988 69958
rect 198836 68883 198892 68922
rect 198836 68866 198838 68883
rect 198838 68866 198890 68883
rect 198890 68866 198892 68883
rect 198740 68274 198796 68330
rect 199028 68422 199084 68478
rect 198932 67682 198988 67738
rect 199124 66794 199180 66850
rect 198932 66054 198988 66110
rect 198740 65923 198796 65962
rect 198740 65906 198742 65923
rect 198742 65906 198794 65923
rect 198794 65906 198796 65923
rect 198836 65166 198892 65222
rect 199028 64870 199084 64926
rect 199124 64426 199180 64482
rect 199220 63538 199276 63594
rect 198740 63094 198796 63150
rect 198836 62798 198892 62854
rect 198932 61910 198988 61966
rect 199028 61614 199084 61670
rect 199124 61170 199180 61226
rect 198740 60299 198796 60338
rect 198740 60282 198742 60299
rect 198742 60282 198794 60299
rect 198794 60282 198796 60299
rect 198836 59690 198892 59746
rect 198932 59542 198988 59598
rect 200276 222046 200332 222102
rect 200180 221306 200236 221362
rect 200468 221750 200524 221806
rect 200372 220714 200428 220770
rect 200564 219826 200620 219882
rect 207284 273419 207340 273458
rect 207284 273402 207286 273419
rect 207286 273402 207338 273419
rect 207338 273402 207340 273419
rect 208436 273254 208492 273310
rect 202580 228706 202636 228762
rect 202580 227670 202636 227726
rect 201236 221306 201292 221362
rect 201140 219826 201196 219882
rect 200756 219678 200812 219734
rect 200372 202806 200428 202862
rect 200948 202806 201004 202862
rect 200852 181346 200908 181402
rect 200948 166842 201004 166898
rect 200756 126734 200812 126790
rect 200948 126734 201004 126790
rect 200756 82926 200812 82982
rect 200756 71530 200812 71586
rect 201332 220714 201388 220770
rect 201332 55546 201388 55602
rect 161300 46683 161356 46722
rect 161300 46666 161302 46683
rect 161302 46666 161354 46683
rect 161354 46666 161356 46683
rect 181364 46683 181420 46722
rect 181364 46666 181366 46683
rect 181366 46666 181418 46683
rect 181418 46666 181420 46683
rect 202868 53326 202924 53382
rect 203060 52734 203116 52790
rect 203156 52586 203212 52642
rect 204020 62206 204076 62262
rect 203540 53474 203596 53530
rect 204500 230038 204556 230094
rect 203924 52882 203980 52938
rect 204404 58062 204460 58118
rect 204884 230334 204940 230390
rect 204980 230038 205036 230094
rect 205460 230186 205516 230242
rect 205460 223970 205516 224026
rect 205844 223822 205900 223878
rect 212948 238770 213004 238826
rect 218804 260565 218806 260582
rect 218806 260565 218858 260582
rect 218858 260565 218860 260582
rect 218804 260526 218860 260565
rect 221492 238474 221548 238530
rect 237044 263190 237100 263246
rect 247892 273550 247948 273606
rect 247892 273254 247948 273310
rect 256340 273293 256342 273310
rect 256342 273293 256394 273310
rect 256394 273293 256396 273310
rect 256340 273254 256396 273293
rect 276404 273698 276460 273754
rect 282164 273737 282166 273754
rect 282166 273737 282218 273754
rect 282218 273737 282220 273754
rect 282164 273698 282220 273737
rect 282356 245282 282412 245338
rect 282260 244729 282262 244746
rect 282262 244729 282314 244746
rect 282314 244729 282316 244746
rect 282260 244690 282316 244729
rect 282260 243654 282316 243710
rect 227444 238326 227500 238382
rect 213044 234922 213100 234978
rect 208052 230334 208108 230390
rect 208436 230334 208492 230390
rect 207860 226782 207916 226838
rect 207764 226634 207820 226690
rect 208148 226486 208204 226542
rect 208052 223822 208108 223878
rect 208436 223822 208492 223878
rect 282548 257566 282604 257622
rect 282452 242470 282508 242526
rect 282356 242322 282412 242378
rect 282836 253274 282892 253330
rect 282740 249574 282796 249630
rect 283124 248834 283180 248890
rect 283028 243062 283084 243118
rect 283700 266742 283756 266798
rect 283796 266446 283852 266502
rect 283700 251202 283756 251258
rect 283892 266298 283948 266354
rect 283796 250166 283852 250222
rect 283892 248982 283948 249038
rect 284276 244098 284332 244154
rect 284948 241434 285004 241490
rect 285908 248094 285964 248150
rect 285812 247206 285868 247262
rect 287828 252978 287884 253034
rect 288020 249278 288076 249334
rect 288212 253866 288268 253922
rect 288212 248686 288268 248742
rect 288500 251054 288556 251110
rect 288404 249278 288460 249334
rect 288212 248242 288268 248298
rect 288020 242174 288076 242230
rect 288500 248834 288556 248890
rect 288500 248242 288556 248298
rect 288404 242174 288460 242230
rect 288404 240250 288460 240306
rect 289172 254754 289228 254810
rect 288884 252978 288940 253034
rect 289172 252978 289228 253034
rect 289556 267038 289612 267094
rect 289460 252978 289516 253034
rect 289940 266890 289996 266946
rect 290324 266594 290380 266650
rect 290708 265854 290764 265910
rect 291092 265706 291148 265762
rect 299444 273737 299446 273754
rect 299446 273737 299498 273754
rect 299498 273737 299500 273754
rect 299444 273698 299500 273737
rect 291476 262006 291532 262062
rect 291764 261858 291820 261914
rect 292148 261710 292204 261766
rect 292532 261562 292588 261618
rect 292916 261414 292972 261470
rect 293300 261266 293356 261322
rect 293204 253274 293260 253330
rect 293972 261118 294028 261174
rect 294356 260970 294412 261026
rect 294740 260822 294796 260878
rect 295124 260674 295180 260730
rect 295508 260526 295564 260582
rect 295316 252978 295372 253034
rect 299636 260378 299692 260434
rect 300788 256678 300844 256734
rect 302324 273698 302380 273754
rect 302324 273402 302380 273458
rect 312404 264374 312460 264430
rect 318644 264374 318700 264430
rect 319700 273737 319702 273754
rect 319702 273737 319754 273754
rect 319754 273737 319756 273754
rect 319700 273698 319756 273737
rect 309140 260378 309196 260434
rect 310868 256678 310924 256734
rect 310964 256530 311020 256586
rect 314996 260082 315052 260138
rect 319028 256826 319084 256882
rect 317972 256678 318028 256734
rect 317204 256530 317260 256586
rect 315668 254014 315724 254070
rect 316724 254014 316780 254070
rect 316436 253718 316492 253774
rect 318644 253422 318700 253478
rect 319700 256086 319756 256142
rect 322676 267926 322732 267982
rect 322004 256974 322060 257030
rect 320180 256826 320236 256882
rect 319700 254162 319756 254218
rect 319412 253718 319468 253774
rect 320468 256086 320524 256142
rect 321236 254162 321292 254218
rect 322580 254606 322636 254662
rect 322580 254014 322636 254070
rect 322676 253866 322732 253922
rect 323828 254162 323884 254218
rect 323444 254014 323500 254070
rect 324884 254606 324940 254662
rect 324500 254310 324556 254366
rect 325268 254310 325324 254366
rect 327092 260230 327148 260286
rect 327476 260378 327532 260434
rect 329204 264966 329260 265022
rect 330740 263930 330796 263986
rect 330452 262598 330508 262654
rect 330932 263634 330988 263690
rect 330836 262746 330892 262802
rect 332660 264522 332716 264578
rect 331124 263782 331180 263838
rect 332276 262450 332332 262506
rect 333044 264374 333100 264430
rect 333428 264226 333484 264282
rect 333716 264078 333772 264134
rect 334004 263486 334060 263542
rect 334004 257418 334060 257474
rect 335636 263930 335692 263986
rect 334484 259934 334540 259990
rect 335924 263782 335980 263838
rect 336308 263634 336364 263690
rect 336692 263486 336748 263542
rect 339764 273550 339820 273606
rect 339764 267965 339766 267982
rect 339766 267965 339818 267982
rect 339818 267965 339820 267982
rect 339764 267926 339820 267965
rect 338708 264966 338764 265022
rect 337460 255938 337516 255994
rect 337460 254606 337516 254662
rect 344564 268074 344620 268130
rect 345044 254606 345100 254662
rect 348404 273402 348460 273458
rect 348596 273402 348652 273458
rect 348212 268091 348268 268130
rect 348212 268074 348214 268091
rect 348214 268074 348266 268091
rect 348266 268074 348268 268091
rect 351476 257122 351532 257178
rect 359348 255642 359404 255698
rect 364436 255494 364492 255550
rect 364340 255346 364396 255402
rect 367124 258750 367180 258806
rect 367796 258602 367852 258658
rect 367604 258454 367660 258510
rect 370292 258306 370348 258362
rect 371444 258898 371500 258954
rect 377780 255198 377836 255254
rect 380180 268113 380182 268130
rect 380182 268113 380234 268130
rect 380234 268113 380236 268130
rect 380180 268074 380236 268113
rect 378452 257270 378508 257326
rect 382196 265410 382252 265466
rect 383444 265558 383500 265614
rect 383156 257122 383212 257178
rect 383444 255050 383500 255106
rect 385652 265410 385708 265466
rect 384500 263190 384556 263246
rect 387476 264670 387532 264726
rect 387284 254754 387340 254810
rect 388436 257270 388492 257326
rect 389780 265558 389836 265614
rect 389972 254902 390028 254958
rect 391604 259046 391660 259102
rect 398900 268518 398956 268574
rect 398132 268074 398188 268130
rect 397076 257122 397132 257178
rect 401204 268518 401260 268574
rect 403124 273567 403180 273606
rect 403124 273550 403126 273567
rect 403126 273550 403178 273567
rect 403178 273550 403180 273567
rect 410708 273846 410764 273902
rect 410420 273254 410476 273310
rect 409556 268666 409612 268722
rect 416660 268814 416716 268870
rect 417812 268222 417868 268278
rect 419348 268814 419404 268870
rect 423572 269850 423628 269906
rect 420980 259046 421036 259102
rect 414740 258898 414796 258954
rect 411764 258750 411820 258806
rect 409556 257270 409612 257326
rect 408980 256086 409036 256142
rect 408980 255790 409036 255846
rect 410708 255642 410764 255698
rect 409940 255198 409996 255254
rect 410324 254902 410380 254958
rect 410996 253422 411052 253478
rect 413204 258454 413260 258510
rect 412532 258306 412588 258362
rect 412916 257122 412972 257178
rect 413588 253126 413644 253182
rect 415124 258602 415180 258658
rect 419156 255494 419212 255550
rect 418772 255050 418828 255106
rect 417620 254754 417676 254810
rect 416180 253718 416236 253774
rect 415412 252978 415468 253034
rect 415796 252978 415852 253034
rect 418388 253866 418444 253922
rect 419828 255346 419884 255402
rect 419540 253570 419596 253626
rect 423764 268962 423820 269018
rect 425012 268370 425068 268426
rect 424628 256382 424684 256438
rect 424244 256234 424300 256290
rect 424436 256234 424492 256290
rect 421556 255790 421612 255846
rect 421748 255790 421804 255846
rect 425396 254458 425452 254514
rect 425876 269702 425932 269758
rect 426356 270442 426412 270498
rect 426164 268962 426220 269018
rect 426836 259934 426892 259990
rect 427220 262746 427276 262802
rect 427124 262598 427180 262654
rect 426068 257418 426124 257474
rect 425684 254458 425740 254514
rect 425684 253422 425740 253478
rect 428468 269998 428524 270054
rect 429236 273402 429292 273458
rect 429044 273254 429100 273310
rect 429140 266002 429196 266058
rect 430292 270590 430348 270646
rect 430100 270294 430156 270350
rect 429716 262450 429772 262506
rect 431156 269258 431212 269314
rect 430964 262894 431020 262950
rect 432020 266150 432076 266206
rect 432212 270146 432268 270202
rect 432308 265854 432364 265910
rect 432116 265706 432172 265762
rect 432788 269998 432844 270054
rect 433268 269702 433324 269758
rect 433460 269406 433516 269462
rect 434228 257566 434284 257622
rect 434900 267778 434956 267834
rect 435956 269110 436012 269166
rect 435668 258158 435724 258214
rect 435284 258010 435340 258066
rect 437780 273441 437782 273458
rect 437782 273441 437834 273458
rect 437834 273441 437836 273458
rect 437780 273402 437836 273441
rect 437204 269554 437260 269610
rect 437876 268370 437932 268426
rect 437876 268074 437932 268130
rect 439316 270294 439372 270350
rect 438068 263042 438124 263098
rect 437012 254310 437068 254366
rect 437012 253422 437068 253478
rect 439028 255198 439084 255254
rect 439508 254902 439564 254958
rect 440468 268370 440524 268426
rect 443540 273698 443596 273754
rect 444020 270590 444076 270646
rect 442868 270442 442924 270498
rect 441620 263338 441676 263394
rect 440276 252978 440332 253034
rect 440660 254458 440716 254514
rect 440756 254310 440812 254366
rect 449972 270590 450028 270646
rect 451124 270442 451180 270498
rect 448820 267630 448876 267686
rect 443540 254458 443596 254514
rect 443636 254310 443692 254366
rect 444308 254014 444364 254070
rect 444980 253274 445036 253330
rect 445364 253422 445420 253478
rect 445364 252995 445420 253034
rect 445364 252978 445366 252995
rect 445366 252978 445418 252995
rect 445418 252978 445420 252995
rect 446228 252978 446284 253034
rect 446420 254310 446476 254366
rect 446420 254201 446422 254218
rect 446422 254201 446474 254218
rect 446474 254201 446476 254218
rect 446420 254162 446476 254201
rect 446420 252978 446476 253034
rect 447476 257714 447532 257770
rect 448148 257862 448204 257918
rect 455924 264818 455980 264874
rect 288980 239510 289036 239566
rect 289748 239510 289804 239566
rect 289556 239362 289612 239418
rect 290900 239510 290956 239566
rect 291188 239527 291244 239566
rect 291188 239510 291190 239527
rect 291190 239510 291242 239527
rect 291242 239510 291244 239527
rect 291380 239510 291436 239566
rect 291572 239510 291628 239566
rect 291956 239510 292012 239566
rect 292340 239510 292396 239566
rect 292724 239510 292780 239566
rect 293108 239510 293164 239566
rect 293108 239362 293164 239418
rect 293396 239362 293452 239418
rect 293780 239066 293836 239122
rect 294932 239510 294988 239566
rect 295316 236106 295372 236162
rect 294548 235958 294604 236014
rect 295988 238918 296044 238974
rect 295604 235810 295660 235866
rect 296564 236402 296620 236458
rect 296756 235662 296812 235718
rect 296372 235514 296428 235570
rect 297812 239214 297868 239270
rect 298004 238918 298060 238974
rect 298004 238622 298060 238678
rect 297524 235810 297580 235866
rect 298964 236402 299020 236458
rect 300500 237142 300556 237198
rect 301556 237882 301612 237938
rect 301172 237438 301228 237494
rect 301940 236994 301996 237050
rect 300788 236846 300844 236902
rect 300116 236698 300172 236754
rect 299732 236550 299788 236606
rect 299348 236254 299404 236310
rect 298580 235366 298636 235422
rect 297140 235070 297196 235126
rect 302708 234182 302764 234238
rect 302996 233442 303052 233498
rect 303764 227374 303820 227430
rect 303380 227078 303436 227134
rect 304532 226930 304588 226986
rect 305108 238178 305164 238234
rect 305204 227226 305260 227282
rect 306740 226634 306796 226690
rect 307412 226782 307468 226838
rect 310388 234774 310444 234830
rect 309620 234626 309676 234682
rect 313364 235218 313420 235274
rect 312596 235070 312652 235126
rect 314804 235662 314860 235718
rect 315572 235366 315628 235422
rect 316244 235514 316300 235570
rect 308180 226190 308236 226246
rect 305972 226042 306028 226098
rect 325556 237734 325612 237790
rect 325940 237734 325996 237790
rect 326900 226338 326956 226394
rect 331028 232702 331084 232758
rect 330644 232406 330700 232462
rect 332852 232850 332908 232906
rect 331700 232258 331756 232314
rect 337940 231370 337996 231426
rect 338516 235958 338572 236014
rect 341300 234922 341356 234978
rect 341684 238918 341740 238974
rect 342452 238622 342508 238678
rect 342740 235810 342796 235866
rect 343124 232554 343180 232610
rect 342836 230926 342892 230982
rect 342068 230778 342124 230834
rect 345620 238195 345676 238234
rect 345620 238178 345622 238195
rect 345622 238178 345674 238195
rect 345674 238178 345676 238195
rect 345908 238178 345964 238234
rect 343892 237734 343948 237790
rect 343796 227670 343852 227726
rect 343508 224266 343564 224322
rect 347540 238178 347596 238234
rect 347156 238030 347212 238086
rect 344948 228262 345004 228318
rect 345332 228114 345388 228170
rect 345716 227522 345772 227578
rect 348020 224562 348076 224618
rect 348404 226486 348460 226542
rect 348788 234774 348844 234830
rect 348788 225894 348844 225950
rect 349172 223822 349228 223878
rect 351764 234626 351820 234682
rect 351764 225746 351820 225802
rect 353684 237290 353740 237346
rect 353012 229002 353068 229058
rect 354548 237142 354604 237198
rect 354068 229485 354070 229502
rect 354070 229485 354122 229502
rect 354122 229485 354124 229502
rect 354068 229446 354124 229485
rect 354164 229150 354220 229206
rect 354836 236846 354892 236902
rect 355124 234774 355180 234830
rect 356180 231074 356236 231130
rect 357044 236994 357100 237050
rect 357044 235958 357100 236014
rect 356756 234922 356812 234978
rect 357524 234626 357580 234682
rect 358196 236106 358252 236162
rect 358292 235662 358348 235718
rect 358868 235070 358924 235126
rect 358772 229446 358828 229502
rect 358484 228410 358540 228466
rect 358388 227818 358444 227874
rect 359156 236698 359212 236754
rect 358964 233590 359020 233646
rect 359156 227818 359212 227874
rect 358868 225450 358924 225506
rect 359444 235218 359500 235274
rect 359444 225598 359500 225654
rect 359540 223822 359596 223878
rect 360500 236550 360556 236606
rect 360308 235810 360364 235866
rect 360116 235662 360172 235718
rect 360500 235662 360556 235718
rect 359732 233886 359788 233942
rect 360020 230334 360076 230390
rect 360692 235810 360748 235866
rect 360500 223970 360556 224026
rect 361076 228410 361132 228466
rect 362228 235514 362284 235570
rect 362420 235366 362476 235422
rect 362612 235218 362668 235274
rect 363380 234034 363436 234090
rect 362708 223822 362764 223878
rect 364148 235070 364204 235126
rect 364244 223839 364300 223878
rect 364244 223822 364246 223839
rect 364246 223822 364298 223839
rect 364298 223822 364300 223839
rect 365396 235366 365452 235422
rect 367028 235514 367084 235570
rect 367124 224118 367180 224174
rect 367796 229150 367852 229206
rect 368084 229611 368140 229650
rect 368564 235958 368620 236014
rect 368084 229594 368086 229611
rect 368086 229594 368138 229611
rect 368138 229594 368140 229611
rect 369236 229298 369292 229354
rect 370004 235662 370060 235718
rect 371348 235810 371404 235866
rect 370676 229002 370732 229058
rect 372212 230482 372268 230538
rect 373364 229611 373420 229650
rect 373364 229594 373366 229611
rect 373366 229594 373418 229611
rect 373418 229594 373420 229611
rect 374324 228410 374380 228466
rect 377396 231518 377452 231574
rect 378164 229890 378220 229946
rect 378932 228706 378988 228762
rect 379412 223839 379468 223878
rect 379412 223822 379414 223839
rect 379414 223822 379466 223839
rect 379466 223822 379468 223839
rect 379604 230038 379660 230094
rect 380276 233146 380332 233202
rect 383348 236994 383404 237050
rect 383252 231666 383308 231722
rect 381812 229742 381868 229798
rect 381140 227670 381196 227726
rect 382580 228558 382636 228614
rect 383636 232998 383692 233054
rect 384404 233294 384460 233350
rect 383924 230186 383980 230242
rect 385172 237290 385228 237346
rect 385076 234478 385132 234534
rect 384692 229446 384748 229502
rect 385556 239510 385612 239566
rect 385460 229594 385516 229650
rect 385844 234330 385900 234386
rect 387956 236698 388012 236754
rect 386228 225006 386284 225062
rect 385844 224858 385900 224914
rect 388340 238770 388396 238826
rect 389876 239066 389932 239122
rect 389492 236846 389548 236902
rect 389684 232110 389740 232166
rect 389684 231222 389740 231278
rect 388724 224710 388780 224766
rect 388724 223822 388780 223878
rect 390644 238918 390700 238974
rect 390356 223822 390412 223878
rect 392084 238770 392140 238826
rect 392468 238474 392524 238530
rect 392660 238474 392716 238530
rect 391028 225154 391084 225210
rect 391700 224710 391756 224766
rect 391892 224118 391948 224174
rect 391700 223822 391756 223878
rect 392756 224118 392812 224174
rect 393044 228114 393100 228170
rect 393140 227966 393196 228022
rect 393236 225302 393292 225358
rect 394388 224414 394444 224470
rect 394964 224710 395020 224766
rect 396500 238326 396556 238382
rect 396308 237586 396364 237642
rect 396500 237586 396556 237642
rect 396308 236550 396364 236606
rect 395444 228114 395500 228170
rect 395924 223970 395980 224026
rect 397364 231814 397420 231870
rect 398132 230630 398188 230686
rect 398516 239214 398572 239270
rect 398804 237290 398860 237346
rect 398804 236994 398860 237050
rect 398996 233442 399052 233498
rect 399188 236994 399244 237050
rect 399380 236994 399436 237050
rect 398900 227818 398956 227874
rect 398900 223970 398956 224026
rect 399668 234182 399724 234238
rect 399668 223822 399724 223878
rect 400244 234182 400300 234238
rect 400244 225006 400300 225062
rect 400244 223822 400300 223878
rect 401204 233442 401260 233498
rect 401876 233755 401932 233794
rect 401876 233738 401878 233755
rect 401878 233738 401930 233755
rect 401930 233738 401932 233755
rect 403220 237438 403276 237494
rect 402260 230351 402316 230390
rect 402260 230334 402262 230351
rect 402262 230334 402314 230351
rect 402314 230334 402316 230351
rect 403028 225006 403084 225062
rect 403316 233590 403372 233646
rect 403316 228114 403372 228170
rect 404468 236846 404524 236902
rect 404468 233886 404524 233942
rect 404372 230334 404428 230390
rect 405236 236106 405292 236162
rect 405428 236106 405484 236162
rect 406100 237882 406156 237938
rect 406100 234182 406156 234238
rect 406676 236550 406732 236606
rect 406292 234182 406348 234238
rect 406580 231814 406636 231870
rect 406868 236550 406924 236606
rect 406388 231222 406444 231278
rect 406580 231222 406636 231278
rect 407252 233738 407308 233794
rect 406964 231814 407020 231870
rect 408212 237438 408268 237494
rect 408884 239527 408940 239566
rect 408404 233886 408460 233942
rect 408884 239510 408886 239527
rect 408886 239510 408938 239527
rect 408938 239510 408940 239527
rect 408884 239362 408940 239418
rect 408788 236846 408844 236902
rect 408692 233442 408748 233498
rect 408980 233442 409036 233498
rect 408884 228114 408940 228170
rect 409076 230334 409132 230390
rect 409460 233886 409516 233942
rect 409364 228114 409420 228170
rect 409652 228114 409708 228170
rect 410708 239510 410764 239566
rect 410900 233590 410956 233646
rect 411764 239510 411820 239566
rect 411764 237882 411820 237938
rect 411284 237586 411340 237642
rect 411764 236106 411820 236162
rect 411764 234182 411820 234238
rect 412340 234182 412396 234238
rect 413492 233442 413548 233498
rect 412628 232110 412684 232166
rect 413396 231962 413452 232018
rect 413108 230334 413164 230390
rect 413972 237586 414028 237642
rect 414356 233886 414412 233942
rect 413972 228114 414028 228170
rect 413972 227818 414028 227874
rect 414164 227818 414220 227874
rect 414452 233590 414508 233646
rect 415508 239362 415564 239418
rect 414548 232110 414604 232166
rect 414644 231962 414700 232018
rect 416756 233738 416812 233794
rect 415220 230334 415276 230390
rect 416372 228854 416428 228910
rect 416564 228854 416620 228910
rect 418292 233442 418348 233498
rect 420116 236106 420172 236162
rect 419348 226930 419404 226986
rect 418964 225746 419020 225802
rect 419252 226042 419308 226098
rect 419540 225894 419596 225950
rect 420884 236106 420940 236162
rect 421940 239362 421996 239418
rect 421940 237882 421996 237938
rect 423380 233442 423436 233498
rect 424244 236106 424300 236162
rect 422324 228854 422380 228910
rect 420596 226042 420652 226098
rect 420788 226042 420844 226098
rect 420500 225598 420556 225654
rect 420692 225598 420748 225654
rect 420980 225615 421036 225654
rect 420980 225598 420982 225615
rect 420982 225598 421034 225615
rect 421034 225598 421036 225615
rect 421940 225450 421996 225506
rect 423380 227391 423436 227430
rect 423380 227374 423382 227391
rect 423382 227374 423434 227391
rect 423434 227374 423436 227391
rect 423476 227265 423478 227282
rect 423478 227265 423530 227282
rect 423530 227265 423532 227282
rect 423476 227226 423532 227265
rect 423380 227095 423436 227134
rect 423380 227078 423382 227095
rect 423382 227078 423434 227095
rect 423434 227078 423436 227095
rect 423188 225746 423244 225802
rect 423572 226634 423628 226690
rect 423668 226042 423724 226098
rect 423956 225450 424012 225506
rect 425876 228854 425932 228910
rect 426068 227078 426124 227134
rect 427988 231814 428044 231870
rect 426164 226634 426220 226690
rect 426260 226525 426262 226542
rect 426262 226525 426314 226542
rect 426314 226525 426316 226542
rect 426260 226486 426316 226525
rect 426164 225598 426220 225654
rect 426260 225341 426262 225358
rect 426262 225341 426314 225358
rect 426314 225341 426316 225358
rect 426260 225302 426316 225341
rect 426356 224710 426412 224766
rect 426548 224727 426604 224766
rect 426548 224710 426550 224727
rect 426550 224710 426602 224727
rect 426602 224710 426604 224727
rect 427604 226930 427660 226986
rect 427508 226782 427564 226838
rect 427796 226782 427852 226838
rect 427316 225598 427372 225654
rect 428084 226486 428140 226542
rect 429044 232110 429100 232166
rect 428852 230778 428908 230834
rect 428276 226042 428332 226098
rect 428180 225302 428236 225358
rect 429236 225746 429292 225802
rect 429428 225746 429484 225802
rect 429620 223822 429676 223878
rect 430388 224710 430444 224766
rect 430772 226338 430828 226394
rect 431156 226190 431212 226246
rect 430772 224858 430828 224914
rect 432596 227522 432652 227578
rect 432308 227078 432364 227134
rect 432500 227078 432556 227134
rect 432116 226634 432172 226690
rect 432308 226634 432364 226690
rect 431924 226338 431980 226394
rect 431828 225894 431884 225950
rect 431732 225598 431788 225654
rect 431540 224710 431596 224766
rect 431732 224710 431788 224766
rect 432116 226338 432172 226394
rect 432020 225598 432076 225654
rect 435284 237882 435340 237938
rect 435380 234034 435436 234090
rect 435284 232554 435340 232610
rect 435092 231814 435148 231870
rect 432884 227226 432940 227282
rect 433076 227226 433132 227282
rect 432884 225746 432940 225802
rect 432884 225598 432940 225654
rect 433076 225598 433132 225654
rect 433268 224858 433324 224914
rect 433460 224858 433516 224914
rect 435188 227374 435244 227430
rect 435572 234034 435628 234090
rect 435476 232554 435532 232610
rect 435860 231814 435916 231870
rect 436820 231962 436876 232018
rect 436916 230926 436972 230982
rect 437780 239601 437836 239603
rect 437780 239549 437782 239601
rect 437782 239549 437834 239601
rect 437834 239549 437836 239601
rect 437780 239547 437836 239549
rect 437588 228854 437644 228910
rect 438452 231962 438508 232018
rect 440084 231370 440140 231426
rect 439988 230926 440044 230982
rect 440564 231370 440620 231426
rect 440564 228854 440620 228910
rect 441044 230926 441100 230982
rect 441428 236106 441484 236162
rect 441524 234182 441580 234238
rect 442676 239362 442732 239418
rect 442676 237290 442732 237346
rect 442772 230778 442828 230834
rect 443540 239362 443596 239418
rect 443732 239549 443734 239566
rect 443734 239549 443786 239566
rect 443786 239549 443788 239566
rect 443732 239510 443788 239549
rect 444308 239362 444364 239418
rect 444116 239214 444172 239270
rect 444404 239214 444460 239270
rect 443636 236106 443692 236162
rect 443636 233590 443692 233646
rect 444116 233590 444172 233646
rect 443924 233442 443980 233498
rect 443540 232110 443596 232166
rect 443636 230334 443692 230390
rect 438260 226190 438316 226246
rect 438548 226042 438604 226098
rect 439892 223970 439948 224026
rect 440660 223970 440716 224026
rect 440948 223970 441004 224026
rect 442868 224266 442924 224322
rect 445268 239362 445324 239418
rect 445364 232406 445420 232462
rect 445748 232702 445804 232758
rect 446612 239362 446668 239418
rect 446516 232258 446572 232314
rect 446708 239214 446764 239270
rect 446996 226338 447052 226394
rect 446996 225894 447052 225950
rect 447572 232850 447628 232906
rect 447956 239379 448012 239418
rect 447956 239362 447958 239379
rect 447958 239362 448010 239379
rect 448010 239362 448012 239379
rect 448148 239214 448204 239270
rect 448724 228854 448780 228910
rect 450932 230778 450988 230834
rect 451700 230630 451756 230686
rect 452084 231074 452140 231130
rect 453332 232423 453388 232462
rect 453332 232406 453334 232423
rect 453334 232406 453386 232423
rect 453386 232406 453388 232423
rect 453428 232110 453484 232166
rect 453044 228262 453100 228318
rect 453716 232406 453772 232462
rect 454004 232110 454060 232166
rect 459092 267482 459148 267538
rect 460628 273698 460684 273754
rect 460628 273402 460684 273458
rect 465524 269406 465580 269462
rect 469364 269127 469420 269166
rect 469364 269110 469366 269127
rect 469366 269110 469418 269127
rect 469418 269110 469420 269127
rect 470132 267334 470188 267390
rect 472532 270146 472588 270202
rect 480884 269127 480940 269166
rect 480884 269110 480886 269127
rect 480886 269110 480938 269127
rect 480938 269110 480940 269127
rect 480980 267186 481036 267242
rect 460820 233442 460876 233498
rect 480692 234922 480748 234978
rect 480020 234774 480076 234830
rect 481076 234626 481132 234682
rect 480980 224118 481036 224174
rect 485108 235366 485164 235422
rect 483668 235218 483724 235274
rect 483284 228114 483340 228170
rect 484436 235070 484492 235126
rect 484820 228410 484876 228466
rect 487028 236402 487084 236458
rect 486644 235958 486700 236014
rect 485876 235514 485932 235570
rect 486260 229150 486316 229206
rect 488084 235810 488140 235866
rect 487316 235662 487372 235718
rect 487028 229298 487084 229354
rect 487700 229002 487756 229058
rect 488468 230482 488524 230538
rect 489620 231222 489676 231278
rect 492692 236254 492748 236310
rect 492116 231518 492172 231574
rect 492884 229890 492940 229946
rect 493652 228706 493708 228762
rect 494324 230038 494380 230094
rect 495092 233146 495148 233202
rect 501140 255681 501142 255698
rect 501142 255681 501194 255698
rect 501194 255681 501196 255698
rect 501140 255642 501196 255681
rect 495380 234034 495436 234090
rect 495860 227670 495916 227726
rect 496532 229742 496588 229798
rect 497300 228558 497356 228614
rect 499124 233294 499180 233350
rect 498356 232998 498412 233054
rect 498164 231666 498220 231722
rect 498740 230186 498796 230242
rect 499508 229446 499564 229502
rect 499892 234478 499948 234534
rect 500660 234330 500716 234386
rect 500276 229594 500332 229650
rect 503924 232554 503980 232610
rect 501044 224118 501100 224174
rect 504308 231814 504364 231870
rect 506516 231370 506572 231426
rect 506996 231962 507052 232018
rect 508340 230926 508396 230982
rect 509876 238030 509932 238086
rect 509876 232110 509932 232166
rect 509780 224414 509836 224470
rect 514964 262154 515020 262210
rect 512852 238178 512908 238234
rect 529844 273402 529900 273458
rect 530036 273254 530092 273310
rect 538484 267186 538540 267242
rect 538484 255659 538540 255661
rect 538484 255607 538486 255659
rect 538486 255607 538538 255659
rect 538538 255607 538540 255659
rect 538484 255605 538540 255607
rect 555860 266742 555916 266798
rect 559412 267038 559468 267094
rect 561524 267186 561580 267242
rect 562964 266890 563020 266946
rect 570068 266594 570124 266650
rect 573716 266446 573772 266502
rect 590228 266781 590230 266798
rect 590230 266781 590282 266798
rect 590282 266781 590284 266798
rect 590228 266742 590284 266781
rect 590132 266594 590188 266650
rect 587924 266298 587980 266354
rect 584372 262006 584428 262062
rect 560660 260378 560716 260434
rect 557012 260230 557068 260286
rect 545204 260082 545260 260138
rect 590516 266781 590518 266798
rect 590518 266781 590570 266798
rect 590570 266781 590572 266798
rect 590516 266742 590572 266781
rect 590612 266594 590668 266650
rect 591572 261858 591628 261914
rect 595124 261710 595180 261766
rect 607028 264522 607084 264578
rect 602228 261562 602284 261618
rect 610388 266781 610390 266798
rect 610390 266781 610442 266798
rect 610442 266781 610444 266798
rect 610388 266742 610444 266781
rect 610676 266781 610678 266798
rect 610678 266781 610730 266798
rect 610730 266781 610732 266798
rect 610676 266742 610732 266781
rect 610580 264374 610636 264430
rect 609332 261414 609388 261470
rect 614132 264226 614188 264282
rect 612980 261266 613036 261322
rect 617684 264078 617740 264134
rect 623636 261118 623692 261174
rect 627188 260970 627244 261026
rect 631988 263930 632044 263986
rect 635540 263782 635596 263838
rect 634292 260822 634348 260878
rect 639092 263634 639148 263690
rect 642644 263486 642700 263542
rect 641492 260674 641548 260730
rect 645140 273106 645196 273162
rect 645044 260526 645100 260582
rect 622004 255790 622060 255846
rect 601940 255681 601942 255698
rect 601942 255681 601994 255698
rect 601994 255681 601996 255698
rect 601940 255642 601996 255681
rect 535700 234182 535756 234238
rect 521300 224562 521356 224618
rect 631316 223970 631372 224026
rect 631988 224118 632044 224174
rect 631604 223822 631660 223878
rect 633524 223970 633580 224026
rect 632372 223822 632428 223878
rect 632756 223822 632812 223878
rect 633140 223822 633196 223878
rect 204980 222638 205036 222694
rect 204884 86626 204940 86682
rect 204692 58802 204748 58858
rect 204596 58358 204652 58414
rect 204500 57174 204556 57230
rect 204692 56138 204748 56194
rect 204308 53030 204364 53086
rect 204788 55102 204844 55158
rect 204980 54658 205036 54714
rect 204884 54510 204940 54566
rect 210356 54214 210412 54270
rect 214772 54214 214828 54270
rect 214964 54214 215020 54270
rect 627092 54214 627148 54270
rect 629588 54214 629644 54270
rect 204692 51846 204748 51902
rect 187604 41782 187660 41838
rect 194324 41782 194380 41838
rect 205076 45334 205132 45390
rect 205460 45038 205516 45094
rect 205652 52142 205708 52198
rect 205844 53069 205846 53086
rect 205846 53069 205898 53086
rect 205898 53069 205900 53086
rect 205844 53030 205900 53069
rect 208532 54066 208588 54122
rect 212564 54066 212620 54122
rect 208148 53918 208204 53974
rect 206228 45482 206284 45538
rect 206132 45186 206188 45242
rect 205748 44890 205804 44946
rect 206324 44742 206380 44798
rect 206708 53474 206764 53530
rect 206708 53030 206764 53086
rect 206900 53326 206956 53382
rect 206804 51994 206860 52050
rect 207092 53585 207148 53641
rect 207572 53474 207628 53530
rect 207860 52290 207916 52346
rect 207956 46518 208012 46574
rect 207860 46387 207916 46426
rect 207860 46370 207862 46387
rect 207862 46370 207914 46387
rect 207914 46370 207916 46387
rect 208532 46557 208534 46574
rect 208534 46557 208586 46574
rect 208586 46557 208588 46574
rect 208532 46518 208588 46557
rect 209012 53474 209068 53530
rect 209300 53326 209356 53382
rect 210740 53770 210796 53826
rect 212564 53474 212620 53530
rect 213716 52882 213772 52938
rect 214484 53474 214540 53530
rect 632948 54066 633004 54122
rect 214964 51846 215020 51902
rect 628532 53918 628588 53974
rect 217076 48738 217132 48794
rect 217460 48886 217516 48942
rect 218036 52438 218092 52494
rect 218324 53030 218380 53086
rect 218228 51698 218284 51754
rect 220532 52734 220588 52790
rect 220244 52586 220300 52642
rect 209684 46370 209740 46426
rect 239828 51106 239884 51162
rect 239348 48146 239404 48202
rect 238580 47998 238636 48054
rect 236756 47850 236812 47906
rect 242036 50958 242092 51014
rect 242996 51254 243052 51310
rect 244148 50810 244204 50866
rect 264884 50366 264940 50422
rect 243764 48590 243820 48646
rect 243380 48442 243436 48498
rect 242420 48294 242476 48350
rect 241556 47702 241612 47758
rect 630644 53770 630700 53826
rect 639668 222342 639724 222398
rect 639380 221750 639436 221806
rect 635060 54214 635116 54270
rect 634868 53918 634924 53974
rect 635348 54362 635404 54418
rect 240212 47554 240268 47610
rect 208820 44594 208876 44650
rect 302516 43262 302572 43318
rect 306740 43262 306796 43318
rect 361748 43262 361804 43318
rect 364916 43262 364972 43318
rect 357140 43114 357196 43170
rect 408884 42078 408940 42134
rect 416276 42078 416332 42134
rect 406292 41782 406348 41838
rect 410804 41782 410860 41838
rect 204884 40746 204940 40802
rect 138164 40154 138220 40210
rect 465620 44742 465676 44798
rect 471092 42078 471148 42134
rect 521588 44594 521644 44650
rect 521204 42078 521260 42134
rect 636404 54066 636460 54122
rect 636308 53770 636364 53826
rect 642260 255659 642316 255698
rect 642260 255642 642262 255659
rect 642262 255642 642314 255659
rect 642314 255642 642316 255659
rect 649556 846014 649612 846070
rect 650036 892782 650092 892838
rect 649940 799098 649996 799154
rect 649844 752034 649900 752090
rect 650132 705266 650188 705322
rect 641012 222381 641014 222398
rect 641014 222381 641066 222398
rect 641066 222381 641068 222398
rect 641012 222342 641068 222381
rect 640724 221750 640780 221806
rect 639860 221306 639916 221362
rect 641300 221345 641302 221362
rect 641302 221345 641354 221362
rect 641354 221345 641356 221362
rect 641300 221306 641356 221345
rect 639764 210946 639820 211002
rect 655124 974330 655180 974386
rect 654356 950946 654412 951002
rect 673940 967522 673996 967578
rect 655220 962638 655276 962694
rect 675092 965598 675148 965654
rect 675764 965598 675820 965654
rect 675092 964858 675148 964914
rect 675092 962786 675148 962842
rect 675188 962490 675244 962546
rect 675380 962194 675436 962250
rect 675764 961454 675820 961510
rect 675476 961010 675532 961066
rect 675668 960122 675724 960178
rect 653780 939254 653836 939310
rect 654452 927453 654454 927470
rect 654454 927453 654506 927470
rect 654506 927453 654508 927470
rect 654452 927414 654508 927453
rect 654452 915722 654508 915778
rect 654452 904030 654508 904086
rect 654452 880498 654508 880554
rect 654452 868806 654508 868862
rect 654452 857114 654508 857170
rect 654452 833582 654508 833638
rect 654452 821890 654508 821946
rect 654452 810198 654508 810254
rect 654452 786666 654508 786722
rect 654452 774974 654508 775030
rect 654452 763299 654508 763338
rect 654452 763282 654454 763299
rect 654454 763282 654506 763299
rect 654506 763282 654508 763299
rect 654452 739750 654508 739806
rect 655124 728058 655180 728114
rect 654452 716218 654508 716274
rect 654836 692834 654892 692890
rect 654452 669302 654508 669358
rect 653780 658350 653836 658406
rect 654452 645918 654508 645974
rect 654452 622386 654508 622442
rect 654452 610694 654508 610750
rect 654452 599298 654508 599354
rect 654452 587162 654508 587218
rect 655316 681142 655372 681198
rect 655220 634226 655276 634282
rect 654452 575470 654508 575526
rect 654452 563778 654508 563834
rect 654452 552086 654508 552142
rect 655124 540246 655180 540302
rect 654452 528554 654508 528610
rect 654452 516862 654508 516918
rect 654452 505170 654508 505226
rect 654452 493330 654508 493386
rect 654452 481638 654508 481694
rect 654452 469985 654454 470002
rect 654454 469985 654506 470002
rect 654506 469985 654508 470002
rect 654452 469946 654508 469985
rect 654356 458254 654412 458310
rect 654452 446431 654508 446470
rect 654452 446414 654454 446431
rect 654454 446414 654506 446431
rect 654506 446414 654508 446431
rect 654356 434722 654412 434778
rect 654452 423030 654508 423086
rect 655028 411190 655084 411246
rect 654452 399498 654508 399554
rect 653876 387806 653932 387862
rect 654164 376114 654220 376170
rect 654452 364274 654508 364330
rect 655316 352582 655372 352638
rect 654164 340890 654220 340946
rect 653972 329198 654028 329254
rect 655124 317358 655180 317414
rect 653780 282282 653836 282338
rect 639956 220714 640012 220770
rect 641300 220753 641302 220770
rect 641302 220753 641354 220770
rect 641354 220753 641356 220770
rect 641300 220714 641356 220753
rect 642068 166842 642124 166898
rect 641492 165806 641548 165862
rect 642164 166398 642220 166454
rect 640148 149970 640204 150026
rect 642164 143458 642220 143514
rect 655220 305666 655276 305722
rect 655412 293974 655468 294030
rect 662324 255494 662380 255550
rect 665204 273550 665260 273606
rect 673844 941918 673900 941974
rect 670964 628306 671020 628362
rect 670868 627418 670924 627474
rect 675764 957606 675820 957662
rect 675092 953462 675148 953518
rect 675476 955978 675532 956034
rect 675188 953314 675244 953370
rect 674036 939550 674092 939606
rect 673940 937182 673996 937238
rect 674708 945322 674764 945378
rect 674708 944730 674764 944786
rect 674708 943694 674764 943750
rect 674612 943102 674668 943158
rect 674420 942601 674476 942640
rect 674420 942584 674422 942601
rect 674422 942584 674474 942601
rect 674474 942584 674476 942601
rect 674900 940586 674956 940642
rect 674132 936294 674188 936350
rect 679796 928598 679852 928654
rect 679796 928006 679852 928062
rect 675092 876354 675148 876410
rect 675764 876354 675820 876410
rect 675092 876206 675148 876262
rect 675284 875762 675340 875818
rect 674228 780450 674284 780506
rect 673652 751590 673708 751646
rect 675476 873986 675532 874042
rect 675380 873394 675436 873450
rect 675380 872802 675436 872858
rect 675572 872358 675628 872414
rect 674324 772606 674380 772662
rect 674324 765837 674326 765854
rect 674326 765837 674378 765854
rect 674378 765837 674380 765854
rect 674324 765798 674380 765837
rect 675380 869842 675436 869898
rect 675380 866882 675436 866938
rect 675476 864662 675532 864718
rect 675668 862886 675724 862942
rect 675764 787850 675820 787906
rect 675476 787406 675532 787462
rect 675764 786666 675820 786722
rect 675764 784150 675820 784206
rect 675764 781930 675820 781986
rect 674996 777490 675052 777546
rect 674804 777342 674860 777398
rect 674708 767761 674710 767778
rect 674710 767761 674762 767778
rect 674762 767761 674764 767778
rect 674708 767722 674764 767761
rect 674708 766873 674710 766890
rect 674710 766873 674762 766890
rect 674762 766873 674764 766890
rect 674708 766834 674764 766873
rect 674708 765245 674710 765262
rect 674710 765245 674762 765262
rect 674762 765245 674764 765262
rect 674708 765206 674764 765245
rect 674708 764039 674764 764078
rect 674708 764022 674710 764039
rect 674710 764022 674762 764039
rect 674762 764022 674764 764039
rect 674708 763282 674764 763338
rect 674708 762559 674764 762598
rect 674708 762542 674710 762559
rect 674710 762542 674762 762559
rect 674762 762542 674764 762559
rect 674324 722473 674326 722490
rect 674326 722473 674378 722490
rect 674378 722473 674380 722490
rect 674324 722434 674380 722473
rect 674324 720845 674326 720862
rect 674326 720845 674378 720862
rect 674378 720845 674380 720862
rect 674324 720806 674380 720845
rect 674516 717863 674572 717902
rect 674516 717846 674518 717863
rect 674518 717846 674570 717863
rect 674570 717846 674572 717863
rect 674420 714442 674476 714498
rect 674324 713702 674380 713758
rect 674228 712962 674284 713018
rect 674420 710485 674422 710502
rect 674422 710485 674474 710502
rect 674474 710485 674476 710502
rect 674420 710446 674476 710485
rect 674420 709005 674422 709022
rect 674422 709005 674474 709022
rect 674474 709005 674476 709022
rect 674420 708966 674476 709005
rect 674420 707377 674422 707394
rect 674422 707377 674474 707394
rect 674474 707377 674476 707394
rect 674420 707338 674476 707377
rect 674132 668562 674188 668618
rect 674132 630674 674188 630730
rect 673844 629786 673900 629842
rect 673844 629046 673900 629102
rect 674036 624902 674092 624958
rect 673844 617946 673900 618002
rect 673844 616318 673900 616374
rect 674420 676445 674422 676462
rect 674422 676445 674474 676462
rect 674474 676445 674476 676462
rect 674420 676406 674476 676445
rect 674420 674817 674422 674834
rect 674422 674817 674474 674834
rect 674474 674817 674476 674834
rect 674420 674778 674476 674817
rect 674420 674055 674476 674094
rect 674420 674038 674422 674055
rect 674422 674038 674474 674055
rect 674474 674038 674476 674055
rect 674324 623570 674380 623626
rect 679796 750110 679852 750166
rect 679796 749518 679852 749574
rect 675092 743302 675148 743358
rect 675764 741674 675820 741730
rect 675092 741378 675148 741434
rect 675476 740342 675532 740398
rect 675476 739306 675532 739362
rect 675380 738566 675436 738622
rect 674804 721881 674806 721898
rect 674806 721881 674858 721898
rect 674858 721881 674860 721898
rect 674804 721842 674860 721881
rect 674804 720253 674806 720270
rect 674806 720253 674858 720270
rect 674858 720253 674860 720270
rect 674804 720214 674860 720253
rect 674804 719047 674860 719086
rect 674804 719030 674806 719047
rect 674806 719030 674858 719047
rect 674858 719030 674860 719047
rect 674804 709893 674806 709910
rect 674806 709893 674858 709910
rect 674858 709893 674860 709910
rect 674804 709854 674860 709893
rect 674804 706785 674806 706802
rect 674806 706785 674858 706802
rect 674858 706785 674860 706802
rect 674804 706746 674860 706785
rect 674804 689282 674860 689338
rect 675764 736642 675820 736698
rect 675668 734422 675724 734478
rect 675188 732498 675244 732554
rect 674900 688246 674956 688302
rect 674804 679662 674860 679718
rect 674804 677481 674806 677498
rect 674806 677481 674858 677498
rect 674858 677481 674860 677498
rect 674804 677442 674860 677481
rect 674804 675853 674806 675870
rect 674806 675853 674858 675870
rect 674858 675853 674860 675870
rect 674804 675814 674860 675853
rect 674804 673167 674860 673206
rect 674804 673150 674806 673167
rect 674806 673150 674858 673167
rect 674858 673150 674860 673167
rect 674708 671078 674764 671134
rect 674612 667970 674668 668026
rect 679700 717994 679756 718050
rect 675092 716218 675148 716274
rect 679796 705118 679852 705174
rect 679796 704526 679852 704582
rect 675380 697866 675436 697922
rect 675476 697274 675532 697330
rect 675380 696830 675436 696886
rect 675764 694758 675820 694814
rect 675284 694610 675340 694666
rect 675764 693426 675820 693482
rect 675764 691650 675820 691706
rect 675764 689134 675820 689190
rect 675092 685582 675148 685638
rect 675092 672262 675148 672318
rect 674996 664714 675052 664770
rect 674708 661645 674710 661662
rect 674710 661645 674762 661662
rect 674762 661645 674764 661662
rect 674708 661606 674764 661645
rect 674996 652726 675052 652782
rect 679796 659978 679852 660034
rect 679796 659238 679852 659294
rect 675476 652578 675532 652634
rect 675476 652134 675532 652190
rect 675284 650950 675340 651006
rect 675764 649618 675820 649674
rect 675188 648286 675244 648342
rect 674516 626086 674572 626142
rect 674420 622682 674476 622738
rect 674228 619426 674284 619482
rect 674036 604774 674092 604830
rect 674708 632489 674710 632506
rect 674710 632489 674762 632506
rect 674762 632489 674764 632506
rect 674708 632450 674764 632489
rect 674708 631749 674710 631766
rect 674710 631749 674762 631766
rect 674762 631749 674764 631766
rect 674708 631710 674764 631749
rect 674900 641922 674956 641978
rect 675476 645474 675532 645530
rect 675092 640442 675148 640498
rect 674900 625642 674956 625698
rect 675764 640294 675820 640350
rect 675380 638518 675436 638574
rect 675188 637778 675244 637834
rect 676724 634966 676780 635022
rect 676052 633190 676108 633246
rect 675188 630082 675244 630138
rect 676724 630082 676780 630138
rect 676052 624754 676108 624810
rect 675092 622090 675148 622146
rect 679700 614986 679756 615042
rect 679700 614394 679756 614450
rect 675092 607734 675148 607790
rect 675092 607438 675148 607494
rect 675668 606402 675724 606458
rect 675092 604922 675148 604978
rect 675764 600186 675820 600242
rect 675764 595302 675820 595358
rect 675764 593378 675820 593434
rect 674708 586422 674764 586478
rect 674420 586313 674422 586330
rect 674422 586313 674474 586330
rect 674474 586313 674476 586330
rect 674420 586274 674476 586313
rect 674420 585425 674422 585442
rect 674422 585425 674474 585442
rect 674474 585425 674476 585442
rect 674420 585386 674476 585425
rect 674612 584833 674614 584850
rect 674614 584833 674666 584850
rect 674666 584833 674668 584850
rect 674612 584794 674668 584833
rect 674228 584498 674284 584554
rect 674708 583627 674764 583666
rect 674708 583610 674710 583627
rect 674710 583610 674762 583627
rect 674762 583610 674764 583627
rect 674708 583353 674710 583370
rect 674710 583353 674762 583370
rect 674762 583353 674764 583370
rect 674708 583314 674764 583353
rect 679700 582870 679756 582926
rect 674228 575914 674284 575970
rect 674708 575361 674710 575378
rect 674710 575361 674762 575378
rect 674762 575361 674764 575378
rect 674708 575322 674764 575361
rect 674708 574473 674710 574490
rect 674710 574473 674762 574490
rect 674762 574473 674764 574490
rect 674708 574434 674764 574473
rect 674420 573585 674422 573602
rect 674422 573585 674474 573602
rect 674474 573585 674476 573602
rect 674420 573546 674476 573585
rect 674708 572993 674710 573010
rect 674710 572993 674762 573010
rect 674762 572993 674764 573010
rect 674708 572954 674764 572993
rect 674420 571957 674422 571974
rect 674422 571957 674474 571974
rect 674474 571957 674476 571974
rect 674420 571918 674476 571957
rect 674708 571365 674710 571382
rect 674710 571365 674762 571382
rect 674762 571365 674764 571382
rect 674708 571326 674764 571365
rect 679796 569698 679852 569754
rect 679796 569106 679852 569162
rect 679988 567330 680044 567386
rect 673844 530922 673900 530978
rect 673844 530034 673900 530090
rect 673844 529294 673900 529350
rect 673748 528554 673804 528610
rect 673844 527814 673900 527870
rect 673748 526926 673804 526982
rect 673844 526186 673900 526242
rect 675092 562890 675148 562946
rect 675092 561706 675148 561762
rect 675284 561558 675340 561614
rect 675476 558894 675532 558950
rect 675764 557710 675820 557766
rect 674420 541321 674422 541338
rect 674422 541321 674474 541338
rect 674474 541321 674476 541338
rect 674420 541282 674476 541321
rect 674036 486078 674092 486134
rect 674228 490074 674284 490130
rect 674420 497291 674422 497308
rect 674422 497291 674474 497308
rect 674474 497291 674476 497308
rect 674420 497252 674476 497291
rect 674420 496477 674422 496494
rect 674422 496477 674474 496494
rect 674474 496477 674476 496494
rect 674420 496438 674476 496477
rect 674708 541578 674764 541634
rect 674708 540729 674710 540746
rect 674710 540729 674762 540746
rect 674762 540729 674764 540746
rect 674708 540690 674764 540729
rect 674708 539841 674710 539858
rect 674710 539841 674762 539858
rect 674762 539841 674764 539858
rect 674708 539802 674764 539841
rect 674804 537582 674860 537638
rect 674708 497770 674764 497826
rect 679796 547054 679852 547110
rect 676724 538618 676780 538674
rect 674612 491850 674668 491906
rect 674516 489630 674572 489686
rect 674900 488742 674956 488798
rect 674324 485264 674380 485320
rect 674132 484598 674188 484654
rect 674996 483118 675052 483174
rect 679796 537582 679852 537638
rect 679796 524706 679852 524762
rect 679796 524114 679852 524170
rect 676724 495846 676780 495902
rect 676724 494514 676780 494570
rect 676628 493034 676684 493090
rect 675092 482378 675148 482434
rect 676628 411930 676684 411986
rect 674420 409897 674422 409914
rect 674422 409897 674474 409914
rect 674474 409897 674476 409914
rect 674420 409858 674476 409897
rect 674708 409305 674710 409322
rect 674710 409305 674762 409322
rect 674762 409305 674764 409322
rect 674708 409266 674764 409305
rect 674708 408417 674710 408434
rect 674710 408417 674762 408434
rect 674762 408417 674764 408434
rect 674708 408378 674764 408417
rect 679700 494366 679756 494422
rect 679892 493478 679948 493534
rect 679796 480750 679852 480806
rect 679796 480010 679852 480066
rect 679892 475274 679948 475330
rect 676724 407638 676780 407694
rect 673844 406602 673900 406658
rect 674900 404086 674956 404142
rect 674132 401866 674188 401922
rect 674036 397130 674092 397186
rect 674612 398462 674668 398518
rect 674324 397870 674380 397926
rect 674420 396390 674476 396446
rect 674516 393726 674572 393782
rect 674804 395354 674860 395410
rect 674708 394466 674764 394522
rect 675380 402458 675436 402514
rect 675284 399350 675340 399406
rect 679796 392542 679852 392598
rect 679796 392098 679852 392154
rect 675092 374486 675148 374542
rect 675476 378778 675532 378834
rect 675476 373894 675532 373950
rect 675380 371970 675436 372026
rect 675188 371526 675244 371582
rect 674708 364422 674764 364478
rect 674420 363869 674422 363886
rect 674422 363869 674474 363886
rect 674474 363869 674476 363886
rect 674420 363830 674476 363869
rect 674612 363277 674614 363294
rect 674614 363277 674666 363294
rect 674666 363277 674668 363294
rect 674612 363238 674668 363277
rect 673844 362202 673900 362258
rect 679892 360130 679948 360186
rect 674036 359094 674092 359150
rect 674516 357170 674572 357226
rect 674324 352730 674380 352786
rect 674228 351250 674284 351306
rect 675188 356430 675244 356486
rect 675092 353322 675148 353378
rect 674900 350214 674956 350270
rect 674708 349326 674764 349382
rect 674996 348586 675052 348642
rect 675284 354062 675340 354118
rect 679796 347402 679852 347458
rect 679796 346662 679852 346718
rect 679892 345478 679948 345534
rect 675476 335118 675532 335174
rect 675476 333786 675532 333842
rect 675380 333490 675436 333546
rect 675476 330530 675532 330586
rect 675188 329494 675244 329550
rect 675380 328310 675436 328366
rect 675380 326830 675436 326886
rect 674708 319913 674710 319930
rect 674710 319913 674762 319930
rect 674762 319913 674764 319930
rect 674708 319874 674764 319913
rect 674420 318877 674422 318894
rect 674422 318877 674474 318894
rect 674474 318877 674476 318894
rect 674420 318838 674476 318877
rect 674708 318285 674710 318302
rect 674710 318285 674762 318302
rect 674762 318285 674764 318302
rect 674708 318246 674764 318285
rect 677012 313806 677068 313862
rect 674324 312474 674380 312530
rect 673940 306110 673996 306166
rect 674036 304482 674092 304538
rect 674228 303742 674284 303798
rect 676916 311438 676972 311494
rect 676820 310698 676876 310754
rect 674612 309070 674668 309126
rect 674420 308478 674476 308534
rect 675092 307442 675148 307498
rect 674996 305222 675052 305278
rect 679796 302410 679852 302466
rect 679796 301670 679852 301726
rect 675476 290126 675532 290182
rect 675380 289534 675436 289590
rect 674996 282282 675052 282338
rect 674708 274921 674710 274938
rect 674710 274921 674762 274938
rect 674762 274921 674764 274938
rect 674708 274882 674764 274921
rect 675476 285242 675532 285298
rect 675380 283614 675436 283670
rect 675380 281838 675436 281894
rect 675188 274290 675244 274346
rect 674708 274033 674710 274050
rect 674710 274033 674762 274050
rect 674762 274033 674764 274050
rect 674708 273994 674764 274033
rect 675188 273550 675244 273606
rect 674708 273293 674710 273310
rect 674710 273293 674762 273310
rect 674762 273293 674764 273310
rect 674708 273254 674764 273293
rect 674804 272662 674860 272718
rect 674420 262746 674476 262802
rect 674132 261118 674188 261174
rect 671060 255681 671062 255698
rect 671062 255681 671114 255698
rect 671114 255681 671116 255698
rect 671060 255642 671116 255681
rect 674324 258750 674380 258806
rect 680084 270886 680140 270942
rect 675380 267186 675436 267242
rect 675284 264078 675340 264134
rect 675188 263338 675244 263394
rect 674804 262154 674860 262210
rect 674900 261710 674956 261766
rect 675092 260082 675148 260138
rect 674996 259342 675052 259398
rect 676820 266446 676876 266502
rect 679700 257418 679756 257474
rect 679700 256826 679756 256882
rect 680084 256234 680140 256290
rect 675380 249574 675436 249630
rect 675284 244986 675340 245042
rect 675476 244690 675532 244746
rect 675476 243506 675532 243562
rect 675092 238918 675148 238974
rect 675668 238622 675724 238678
rect 675380 236846 675436 236902
rect 674420 229485 674422 229502
rect 674422 229485 674474 229502
rect 674474 229485 674476 229502
rect 674420 229446 674476 229485
rect 674708 228893 674710 228910
rect 674710 228893 674762 228910
rect 674762 228893 674764 228910
rect 674708 228854 674764 228893
rect 674420 227857 674422 227874
rect 674422 227857 674474 227874
rect 674474 227857 674476 227874
rect 674420 227818 674476 227857
rect 679796 225006 679852 225062
rect 676820 223674 676876 223730
rect 674516 222046 674572 222102
rect 674420 217458 674476 217514
rect 674132 215978 674188 216034
rect 674996 221158 675052 221214
rect 674612 221010 674668 221066
rect 674900 214942 674956 214998
rect 674804 214202 674860 214258
rect 674708 213314 674764 213370
rect 674612 201622 674668 201678
rect 675188 218938 675244 218994
rect 675092 218050 675148 218106
rect 679700 212130 679756 212186
rect 679700 211390 679756 211446
rect 679796 210058 679852 210114
rect 676820 206210 676876 206266
rect 675764 204434 675820 204490
rect 675476 199994 675532 200050
rect 675380 199402 675436 199458
rect 675092 193186 675148 193242
rect 675476 198366 675532 198422
rect 675476 195258 675532 195314
rect 675380 193482 675436 193538
rect 675188 193038 675244 193094
rect 675380 191558 675436 191614
rect 674420 184454 674476 184510
rect 674708 183901 674710 183918
rect 674710 183901 674762 183918
rect 674762 183901 674764 183918
rect 674708 183862 674764 183901
rect 674420 182865 674422 182882
rect 674422 182865 674474 182882
rect 674474 182865 674476 182882
rect 674420 182826 674476 182865
rect 676916 178682 676972 178738
rect 674516 177054 674572 177110
rect 674036 170986 674092 171042
rect 674228 169358 674284 169414
rect 676820 176166 676876 176222
rect 675668 173946 675724 174002
rect 674900 173058 674956 173114
rect 674516 168322 674572 168378
rect 674708 167286 674764 167342
rect 674612 166694 674668 166750
rect 674708 165658 674764 165714
rect 674996 172318 675052 172374
rect 675092 169950 675148 170006
rect 677012 175574 677068 175630
rect 677012 161366 677068 161422
rect 675284 155150 675340 155206
rect 675476 155002 675532 155058
rect 675764 153374 675820 153430
rect 675476 150266 675532 150322
rect 675476 148490 675532 148546
rect 675380 146418 675436 146474
rect 674324 142718 674380 142774
rect 674708 138722 674764 138778
rect 674420 138443 674476 138482
rect 674420 138426 674422 138443
rect 674422 138426 674474 138443
rect 674474 138426 674476 138443
rect 674708 137094 674764 137150
rect 674708 135466 674764 135522
rect 679700 135466 679756 135522
rect 674420 134504 674476 134560
rect 675284 133394 675340 133450
rect 675188 131766 675244 131822
rect 674132 131174 674188 131230
rect 673364 126734 673420 126790
rect 674036 125846 674092 125902
rect 642068 121702 642124 121758
rect 642164 121149 642166 121166
rect 642166 121149 642218 121166
rect 642218 121149 642220 121166
rect 642164 121110 642220 121149
rect 641396 120666 641452 120722
rect 640724 120074 640780 120130
rect 665204 112230 665260 112286
rect 640148 60282 640204 60338
rect 640820 58654 640876 58710
rect 668180 111194 668236 111250
rect 675092 128658 675148 128714
rect 674420 128066 674476 128122
rect 674324 127326 674380 127382
rect 674228 126438 674284 126494
rect 674996 124810 675052 124866
rect 674900 123922 674956 123978
rect 674516 123182 674572 123238
rect 674804 122146 674860 122202
rect 674612 121554 674668 121610
rect 674708 121275 674764 121314
rect 674708 121258 674710 121275
rect 674710 121258 674762 121275
rect 674762 121258 674764 121275
rect 674900 110750 674956 110806
rect 675572 110010 675628 110066
rect 675380 108086 675436 108142
rect 675380 103202 675436 103258
rect 675380 101426 675436 101482
rect 652628 86922 652684 86978
rect 653588 86182 653644 86238
rect 653492 85294 653548 85350
rect 641012 61318 641068 61374
rect 640916 57470 640972 57526
rect 663380 85590 663436 85646
rect 653684 84258 653740 84314
rect 653588 83370 653644 83426
rect 641204 58062 641260 58118
rect 653684 82630 653740 82686
rect 662420 81150 662476 81206
rect 641396 59542 641452 59598
rect 641300 57026 641356 57082
rect 641108 56434 641164 56490
rect 640724 55398 640780 55454
rect 641588 59690 641644 59746
rect 642164 75526 642220 75582
rect 641684 56286 641740 56342
rect 641492 54806 641548 54862
rect 663284 83962 663340 84018
rect 663284 82038 663340 82094
rect 663572 84702 663628 84758
rect 663476 82778 663532 82834
rect 523892 43114 523948 43170
rect 529268 43114 529324 43170
rect 525908 42078 525964 42134
rect 518516 41782 518572 41838
rect 512564 40746 512620 40802
rect 613460 40598 613516 40654
<< metal3 >>
rect 549570 1019912 550782 1019972
rect 549570 1019824 549630 1019912
rect 549216 1019794 549630 1019824
rect 550722 1019794 550782 1019912
rect 549186 1019764 549630 1019794
rect 108687 1005468 108753 1005471
rect 115215 1005468 115281 1005471
rect 321039 1005468 321105 1005471
rect 108687 1005466 109152 1005468
rect 108687 1005410 108692 1005466
rect 108748 1005410 109152 1005466
rect 108687 1005408 109152 1005410
rect 115215 1005466 115488 1005468
rect 115215 1005410 115220 1005466
rect 115276 1005410 115488 1005466
rect 115215 1005408 115488 1005410
rect 320448 1005466 321105 1005468
rect 320448 1005410 321044 1005466
rect 321100 1005410 321105 1005466
rect 320448 1005408 321105 1005410
rect 108687 1005405 108753 1005408
rect 115215 1005405 115281 1005408
rect 321039 1005405 321105 1005408
rect 321423 1005468 321489 1005471
rect 325455 1005468 325521 1005471
rect 358671 1005468 358737 1005471
rect 431631 1005468 431697 1005471
rect 433263 1005468 433329 1005471
rect 504591 1005468 504657 1005471
rect 321423 1005466 325521 1005468
rect 321423 1005410 321428 1005466
rect 321484 1005410 325460 1005466
rect 325516 1005410 325521 1005466
rect 321423 1005408 325521 1005410
rect 358176 1005466 358737 1005468
rect 358176 1005410 358676 1005466
rect 358732 1005410 358737 1005466
rect 358176 1005408 358737 1005410
rect 431040 1005466 431697 1005468
rect 431040 1005410 431636 1005466
rect 431692 1005410 431697 1005466
rect 431040 1005408 431697 1005410
rect 432672 1005466 433329 1005468
rect 432672 1005410 433268 1005466
rect 433324 1005410 433329 1005466
rect 432672 1005408 433329 1005410
rect 504096 1005466 504657 1005468
rect 504096 1005410 504596 1005466
rect 504652 1005410 504657 1005466
rect 504096 1005408 504657 1005410
rect 321423 1005405 321489 1005408
rect 325455 1005405 325521 1005408
rect 358671 1005405 358737 1005408
rect 431631 1005405 431697 1005408
rect 433263 1005405 433329 1005408
rect 504591 1005405 504657 1005408
rect 106575 1005320 106641 1005323
rect 109455 1005320 109521 1005323
rect 217263 1005320 217329 1005323
rect 106575 1005318 106752 1005320
rect 106575 1005262 106580 1005318
rect 106636 1005262 106752 1005318
rect 106575 1005260 106752 1005262
rect 109455 1005318 109920 1005320
rect 109455 1005262 109460 1005318
rect 109516 1005262 109920 1005318
rect 109455 1005260 109920 1005262
rect 216672 1005318 217329 1005320
rect 216672 1005262 217268 1005318
rect 217324 1005262 217329 1005318
rect 216672 1005260 217329 1005262
rect 106575 1005257 106641 1005260
rect 109455 1005257 109521 1005260
rect 217263 1005257 217329 1005260
rect 218895 1005320 218961 1005323
rect 223119 1005320 223185 1005323
rect 218895 1005318 223185 1005320
rect 218895 1005262 218900 1005318
rect 218956 1005262 223124 1005318
rect 223180 1005262 223185 1005318
rect 218895 1005260 223185 1005262
rect 218895 1005257 218961 1005260
rect 223119 1005257 223185 1005260
rect 308751 1005320 308817 1005323
rect 309615 1005320 309681 1005323
rect 365007 1005320 365073 1005323
rect 424527 1005320 424593 1005323
rect 425295 1005320 425361 1005323
rect 434799 1005320 434865 1005323
rect 438735 1005320 438801 1005323
rect 308751 1005318 309312 1005320
rect 308751 1005262 308756 1005318
rect 308812 1005262 309312 1005318
rect 308751 1005260 309312 1005262
rect 309615 1005318 310176 1005320
rect 309615 1005262 309620 1005318
rect 309676 1005262 310176 1005318
rect 309615 1005260 310176 1005262
rect 364512 1005318 365073 1005320
rect 364512 1005262 365012 1005318
rect 365068 1005262 365073 1005318
rect 364512 1005260 365073 1005262
rect 424032 1005318 424593 1005320
rect 424032 1005262 424532 1005318
rect 424588 1005262 424593 1005318
rect 424032 1005260 424593 1005262
rect 424800 1005318 425361 1005320
rect 424800 1005262 425300 1005318
rect 425356 1005262 425361 1005318
rect 424800 1005260 425361 1005262
rect 434304 1005318 434865 1005320
rect 434304 1005262 434804 1005318
rect 434860 1005262 434865 1005318
rect 434304 1005260 434865 1005262
rect 438240 1005318 438801 1005320
rect 438240 1005262 438740 1005318
rect 438796 1005262 438801 1005318
rect 438240 1005260 438801 1005262
rect 308751 1005257 308817 1005260
rect 309615 1005257 309681 1005260
rect 365007 1005257 365073 1005260
rect 424527 1005257 424593 1005260
rect 425295 1005257 425361 1005260
rect 434799 1005257 434865 1005260
rect 438735 1005257 438801 1005260
rect 439695 1005320 439761 1005323
rect 444879 1005320 444945 1005323
rect 502287 1005320 502353 1005323
rect 439695 1005318 444945 1005320
rect 439695 1005262 439700 1005318
rect 439756 1005262 444884 1005318
rect 444940 1005262 444945 1005318
rect 439695 1005260 444945 1005262
rect 501792 1005318 502353 1005320
rect 501792 1005262 502292 1005318
rect 502348 1005262 502353 1005318
rect 501792 1005260 502353 1005262
rect 439695 1005257 439761 1005260
rect 444879 1005257 444945 1005260
rect 502287 1005257 502353 1005260
rect 114159 1005172 114225 1005175
rect 207279 1005172 207345 1005175
rect 221871 1005172 221937 1005175
rect 114159 1005170 114720 1005172
rect 114159 1005114 114164 1005170
rect 114220 1005114 114720 1005170
rect 114159 1005112 114720 1005114
rect 207279 1005170 207936 1005172
rect 207279 1005114 207284 1005170
rect 207340 1005114 207936 1005170
rect 207279 1005112 207936 1005114
rect 218304 1005170 221937 1005172
rect 218304 1005114 221876 1005170
rect 221932 1005114 221937 1005170
rect 218304 1005112 221937 1005114
rect 114159 1005109 114225 1005112
rect 207279 1005109 207345 1005112
rect 221871 1005109 221937 1005112
rect 314223 1005172 314289 1005175
rect 357999 1005172 358065 1005175
rect 426063 1005172 426129 1005175
rect 435567 1005172 435633 1005175
rect 445071 1005172 445137 1005175
rect 498351 1005172 498417 1005175
rect 314223 1005170 314880 1005172
rect 314223 1005114 314228 1005170
rect 314284 1005114 314880 1005170
rect 314223 1005112 314880 1005114
rect 357408 1005170 358065 1005172
rect 357408 1005114 358004 1005170
rect 358060 1005114 358065 1005170
rect 357408 1005112 358065 1005114
rect 425568 1005170 426129 1005172
rect 425568 1005114 426068 1005170
rect 426124 1005114 426129 1005170
rect 425568 1005112 426129 1005114
rect 435168 1005170 435633 1005172
rect 435168 1005114 435572 1005170
rect 435628 1005114 435633 1005170
rect 435168 1005112 435633 1005114
rect 439104 1005170 445137 1005172
rect 439104 1005114 445076 1005170
rect 445132 1005114 445137 1005170
rect 439104 1005112 445137 1005114
rect 497856 1005170 498417 1005172
rect 497856 1005114 498356 1005170
rect 498412 1005114 498417 1005170
rect 497856 1005112 498417 1005114
rect 314223 1005109 314289 1005112
rect 357999 1005109 358065 1005112
rect 426063 1005109 426129 1005112
rect 435567 1005109 435633 1005112
rect 445071 1005109 445137 1005112
rect 498351 1005109 498417 1005112
rect 498735 1005172 498801 1005175
rect 508623 1005172 508689 1005175
rect 498735 1005170 499296 1005172
rect 498735 1005114 498740 1005170
rect 498796 1005114 499296 1005170
rect 498735 1005112 499296 1005114
rect 508032 1005170 508689 1005172
rect 508032 1005114 508628 1005170
rect 508684 1005114 508689 1005170
rect 508032 1005112 508689 1005114
rect 498735 1005109 498801 1005112
rect 508623 1005109 508689 1005112
rect 547119 1005172 547185 1005175
rect 549186 1005172 549246 1019764
rect 554511 1005320 554577 1005323
rect 554016 1005318 554577 1005320
rect 554016 1005262 554516 1005318
rect 554572 1005262 554577 1005318
rect 554016 1005260 554577 1005262
rect 554511 1005257 554577 1005260
rect 553743 1005172 553809 1005175
rect 562479 1005172 562545 1005175
rect 547119 1005170 549246 1005172
rect 547119 1005114 547124 1005170
rect 547180 1005142 549246 1005170
rect 553248 1005170 553809 1005172
rect 547180 1005114 549216 1005142
rect 547119 1005112 549216 1005114
rect 553248 1005114 553748 1005170
rect 553804 1005114 553809 1005170
rect 553248 1005112 553809 1005114
rect 561888 1005170 562545 1005172
rect 561888 1005114 562484 1005170
rect 562540 1005114 562545 1005170
rect 561888 1005112 562545 1005114
rect 547119 1005109 547185 1005112
rect 553743 1005109 553809 1005112
rect 562479 1005109 562545 1005112
rect 356751 1003988 356817 1003991
rect 356640 1003986 356817 1003988
rect 356640 1003930 356756 1003986
rect 356812 1003930 356817 1003986
rect 356640 1003928 356817 1003930
rect 356751 1003925 356817 1003928
rect 355983 1003840 356049 1003843
rect 359055 1003840 359121 1003843
rect 423375 1003840 423441 1003843
rect 428079 1003840 428145 1003843
rect 501135 1003840 501201 1003843
rect 551727 1003840 551793 1003843
rect 556527 1003840 556593 1003843
rect 355776 1003838 356049 1003840
rect 355776 1003782 355988 1003838
rect 356044 1003782 356049 1003838
rect 355776 1003780 356049 1003782
rect 358944 1003838 359121 1003840
rect 358944 1003782 359060 1003838
rect 359116 1003782 359121 1003838
rect 358944 1003780 359121 1003782
rect 423168 1003838 423441 1003840
rect 423168 1003782 423380 1003838
rect 423436 1003782 423441 1003838
rect 423168 1003780 423441 1003782
rect 427872 1003838 428145 1003840
rect 427872 1003782 428084 1003838
rect 428140 1003782 428145 1003838
rect 427872 1003780 428145 1003782
rect 501024 1003838 501201 1003840
rect 501024 1003782 501140 1003838
rect 501196 1003782 501201 1003838
rect 501024 1003780 501201 1003782
rect 551520 1003838 551793 1003840
rect 551520 1003782 551732 1003838
rect 551788 1003782 551793 1003838
rect 551520 1003780 551793 1003782
rect 556320 1003838 556593 1003840
rect 556320 1003782 556532 1003838
rect 556588 1003782 556593 1003838
rect 556320 1003780 556593 1003782
rect 355983 1003777 356049 1003780
rect 359055 1003777 359121 1003780
rect 423375 1003777 423441 1003780
rect 428079 1003777 428145 1003780
rect 501135 1003777 501201 1003780
rect 551727 1003777 551793 1003780
rect 556527 1003777 556593 1003780
rect 211695 1003692 211761 1003695
rect 359919 1003692 359985 1003695
rect 426447 1003692 426513 1003695
rect 500367 1003692 500433 1003695
rect 552591 1003692 552657 1003695
rect 211695 1003690 211872 1003692
rect 211695 1003634 211700 1003690
rect 211756 1003634 211872 1003690
rect 211695 1003632 211872 1003634
rect 359712 1003690 359985 1003692
rect 359712 1003634 359924 1003690
rect 359980 1003634 359985 1003690
rect 359712 1003632 359985 1003634
rect 426336 1003690 426513 1003692
rect 426336 1003634 426452 1003690
rect 426508 1003634 426513 1003690
rect 426336 1003632 426513 1003634
rect 500160 1003690 500433 1003692
rect 500160 1003634 500372 1003690
rect 500428 1003634 500433 1003690
rect 500160 1003632 500433 1003634
rect 552384 1003690 552657 1003692
rect 552384 1003634 552596 1003690
rect 552652 1003634 552657 1003690
rect 552384 1003632 552657 1003634
rect 211695 1003629 211761 1003632
rect 359919 1003629 359985 1003632
rect 426447 1003629 426513 1003632
rect 500367 1003629 500433 1003632
rect 552591 1003629 552657 1003632
rect 151503 1002656 151569 1002659
rect 151503 1002654 151776 1002656
rect 151503 1002598 151508 1002654
rect 151564 1002598 151776 1002654
rect 151503 1002596 151776 1002598
rect 151503 1002593 151569 1002596
rect 152847 1002508 152913 1002511
rect 153615 1002508 153681 1002511
rect 502767 1002508 502833 1002511
rect 503439 1002508 503505 1002511
rect 559119 1002508 559185 1002511
rect 559887 1002508 559953 1002511
rect 152847 1002506 153408 1002508
rect 152847 1002450 152852 1002506
rect 152908 1002450 153408 1002506
rect 152847 1002448 153408 1002450
rect 153615 1002506 154080 1002508
rect 153615 1002450 153620 1002506
rect 153676 1002450 154080 1002506
rect 153615 1002448 154080 1002450
rect 502560 1002506 502833 1002508
rect 502560 1002450 502772 1002506
rect 502828 1002450 502833 1002506
rect 502560 1002448 502833 1002450
rect 503328 1002506 503505 1002508
rect 503328 1002450 503444 1002506
rect 503500 1002450 503505 1002506
rect 503328 1002448 503505 1002450
rect 558816 1002506 559185 1002508
rect 558816 1002450 559124 1002506
rect 559180 1002450 559185 1002506
rect 558816 1002448 559185 1002450
rect 559488 1002506 559953 1002508
rect 559488 1002450 559892 1002506
rect 559948 1002450 559953 1002506
rect 559488 1002448 559953 1002450
rect 152847 1002445 152913 1002448
rect 153615 1002445 153681 1002448
rect 502767 1002445 502833 1002448
rect 503439 1002445 503505 1002448
rect 559119 1002445 559185 1002448
rect 559887 1002445 559953 1002448
rect 150351 1002360 150417 1002363
rect 505071 1002360 505137 1002363
rect 560559 1002360 560625 1002363
rect 561519 1002360 561585 1002363
rect 564783 1002360 564849 1002363
rect 150351 1002358 151008 1002360
rect 150351 1002302 150356 1002358
rect 150412 1002302 151008 1002358
rect 150351 1002300 151008 1002302
rect 504960 1002358 505137 1002360
rect 504960 1002302 505076 1002358
rect 505132 1002302 505137 1002358
rect 504960 1002300 505137 1002302
rect 560256 1002358 560625 1002360
rect 560256 1002302 560564 1002358
rect 560620 1002302 560625 1002358
rect 560256 1002300 560625 1002302
rect 561120 1002358 561585 1002360
rect 561120 1002302 561524 1002358
rect 561580 1002302 561585 1002358
rect 561120 1002300 561585 1002302
rect 564192 1002358 564849 1002360
rect 564192 1002302 564788 1002358
rect 564844 1002302 564849 1002358
rect 564192 1002300 564849 1002302
rect 150351 1002297 150417 1002300
rect 505071 1002297 505137 1002300
rect 560559 1002297 560625 1002300
rect 561519 1002297 561585 1002300
rect 564783 1002297 564849 1002300
rect 434031 1001176 434097 1001179
rect 433536 1001174 434097 1001176
rect 433536 1001118 434036 1001174
rect 434092 1001118 434097 1001174
rect 433536 1001116 434097 1001118
rect 434031 1001113 434097 1001116
rect 430863 1001028 430929 1001031
rect 432495 1001028 432561 1001031
rect 510927 1001028 510993 1001031
rect 430368 1001026 430929 1001028
rect 430368 1000970 430868 1001026
rect 430924 1000970 430929 1001026
rect 430368 1000968 430929 1000970
rect 431904 1001026 432561 1001028
rect 431904 1000970 432500 1001026
rect 432556 1000970 432561 1001026
rect 431904 1000968 432561 1000970
rect 510528 1001026 510993 1001028
rect 510528 1000970 510932 1001026
rect 510988 1000970 510993 1001026
rect 510528 1000968 510993 1000970
rect 430863 1000965 430929 1000968
rect 432495 1000965 432561 1000968
rect 510927 1000965 510993 1000968
rect 516687 1001028 516753 1001031
rect 523599 1001028 523665 1001031
rect 516687 1001026 523665 1001028
rect 516687 1000970 516692 1001026
rect 516748 1000970 523604 1001026
rect 523660 1000970 523665 1001026
rect 516687 1000968 523665 1000970
rect 516687 1000965 516753 1000968
rect 523599 1000965 523665 1000968
rect 160239 1000880 160305 1000883
rect 208143 1000880 208209 1000883
rect 361551 1000880 361617 1000883
rect 427311 1000880 427377 1000883
rect 428943 1000880 429009 1000883
rect 509295 1000880 509361 1000883
rect 160239 1000878 160512 1000880
rect 160239 1000822 160244 1000878
rect 160300 1000822 160512 1000878
rect 160239 1000820 160512 1000822
rect 208143 1000878 208800 1000880
rect 208143 1000822 208148 1000878
rect 208204 1000822 208800 1000878
rect 208143 1000820 208800 1000822
rect 361344 1000878 361617 1000880
rect 361344 1000822 361556 1000878
rect 361612 1000822 361617 1000878
rect 361344 1000820 361617 1000822
rect 427104 1000878 427377 1000880
rect 427104 1000822 427316 1000878
rect 427372 1000822 427377 1000878
rect 427104 1000820 427377 1000822
rect 428736 1000878 429009 1000880
rect 428736 1000822 428948 1000878
rect 429004 1000822 429009 1000878
rect 428736 1000820 429009 1000822
rect 508896 1000878 509361 1000880
rect 508896 1000822 509300 1000878
rect 509356 1000822 509361 1000878
rect 508896 1000820 509361 1000822
rect 160239 1000817 160305 1000820
rect 208143 1000817 208209 1000820
rect 361551 1000817 361617 1000820
rect 427311 1000817 427377 1000820
rect 428943 1000817 429009 1000820
rect 509295 1000817 509361 1000820
rect 516687 1000880 516753 1000883
rect 523695 1000880 523761 1000883
rect 516687 1000878 523761 1000880
rect 516687 1000822 516692 1000878
rect 516748 1000822 523700 1000878
rect 523756 1000822 523761 1000878
rect 516687 1000820 523761 1000822
rect 516687 1000817 516753 1000820
rect 523695 1000817 523761 1000820
rect 516783 1000732 516849 1000735
rect 523503 1000732 523569 1000735
rect 516783 1000730 523569 1000732
rect 516783 1000674 516788 1000730
rect 516844 1000674 523508 1000730
rect 523564 1000674 523569 1000730
rect 516783 1000672 523569 1000674
rect 516783 1000669 516849 1000672
rect 523503 1000669 523569 1000672
rect 523407 999992 523473 999995
rect 521154 999990 523473 999992
rect 521154 999934 523412 999990
rect 523468 999934 523473 999990
rect 521154 999932 523473 999934
rect 155151 999548 155217 999551
rect 258831 999548 258897 999551
rect 260751 999548 260817 999551
rect 516687 999548 516753 999551
rect 521154 999548 521214 999932
rect 523407 999929 523473 999932
rect 521391 999696 521457 999699
rect 523887 999696 523953 999699
rect 521391 999694 523953 999696
rect 521391 999638 521396 999694
rect 521452 999638 523892 999694
rect 523948 999638 523953 999694
rect 521391 999636 523953 999638
rect 521391 999633 521457 999636
rect 523887 999633 523953 999636
rect 155151 999546 155712 999548
rect 155151 999490 155156 999546
rect 155212 999490 155712 999546
rect 155151 999488 155712 999490
rect 258831 999546 259296 999548
rect 258831 999490 258836 999546
rect 258892 999490 259296 999546
rect 258831 999488 259296 999490
rect 260751 999546 261024 999548
rect 260751 999490 260756 999546
rect 260812 999490 261024 999546
rect 260751 999488 261024 999490
rect 516687 999546 521214 999548
rect 516687 999490 516692 999546
rect 516748 999490 521214 999546
rect 516687 999488 521214 999490
rect 521487 999548 521553 999551
rect 524079 999548 524145 999551
rect 521487 999546 524145 999548
rect 521487 999490 521492 999546
rect 521548 999490 524084 999546
rect 524140 999490 524145 999546
rect 521487 999488 524145 999490
rect 155151 999485 155217 999488
rect 258831 999485 258897 999488
rect 260751 999485 260817 999488
rect 516687 999485 516753 999488
rect 521487 999485 521553 999488
rect 524079 999485 524145 999488
rect 156879 999400 156945 999403
rect 259599 999400 259665 999403
rect 311247 999400 311313 999403
rect 488847 999400 488913 999403
rect 497583 999400 497649 999403
rect 506319 999400 506385 999403
rect 156879 999398 157344 999400
rect 156879 999342 156884 999398
rect 156940 999342 157344 999398
rect 156879 999340 157344 999342
rect 259599 999398 260160 999400
rect 259599 999342 259604 999398
rect 259660 999342 260160 999398
rect 259599 999340 260160 999342
rect 311247 999398 311712 999400
rect 311247 999342 311252 999398
rect 311308 999342 311712 999398
rect 311247 999340 311712 999342
rect 488847 999398 497649 999400
rect 488847 999342 488852 999398
rect 488908 999342 497588 999398
rect 497644 999342 497649 999398
rect 488847 999340 497649 999342
rect 505728 999398 506385 999400
rect 505728 999342 506324 999398
rect 506380 999342 506385 999398
rect 505728 999340 506385 999342
rect 156879 999337 156945 999340
rect 259599 999337 259665 999340
rect 311247 999337 311313 999340
rect 488847 999337 488913 999340
rect 497583 999337 497649 999340
rect 506319 999337 506385 999340
rect 516687 999400 516753 999403
rect 523791 999400 523857 999403
rect 516687 999398 523857 999400
rect 516687 999342 516692 999398
rect 516748 999342 523796 999398
rect 523852 999342 523857 999398
rect 516687 999340 523857 999342
rect 516687 999337 516753 999340
rect 523791 999337 523857 999340
rect 209391 997920 209457 997923
rect 367887 997920 367953 997923
rect 555183 997920 555249 997923
rect 557295 997920 557361 997923
rect 209391 997918 209568 997920
rect 209391 997862 209396 997918
rect 209452 997862 209568 997918
rect 209391 997860 209568 997862
rect 367776 997918 367953 997920
rect 367776 997862 367892 997918
rect 367948 997862 367953 997918
rect 367776 997860 367953 997862
rect 554688 997918 555249 997920
rect 554688 997862 555188 997918
rect 555244 997862 555249 997918
rect 554688 997860 555249 997862
rect 557088 997918 557361 997920
rect 557088 997862 557300 997918
rect 557356 997862 557361 997918
rect 557088 997860 557361 997862
rect 209391 997857 209457 997860
rect 367887 997857 367953 997860
rect 555183 997857 555249 997860
rect 557295 997857 557361 997860
rect 318447 997772 318513 997775
rect 318048 997770 318513 997772
rect 318048 997714 318452 997770
rect 318508 997714 318513 997770
rect 318048 997712 318513 997714
rect 318447 997709 318513 997712
rect 369039 997772 369105 997775
rect 556143 997772 556209 997775
rect 369039 997770 369216 997772
rect 369039 997714 369044 997770
rect 369100 997714 369216 997770
rect 369039 997712 369216 997714
rect 555552 997770 556209 997772
rect 555552 997714 556148 997770
rect 556204 997714 556209 997770
rect 555552 997712 556209 997714
rect 369039 997709 369105 997712
rect 556143 997709 556209 997712
rect 74703 997328 74769 997331
rect 74895 997328 74961 997331
rect 74703 997326 74992 997328
rect 74703 997270 74708 997326
rect 74764 997270 74900 997326
rect 74956 997270 74992 997326
rect 74703 997268 74992 997270
rect 74703 997265 74769 997268
rect 74895 997265 74961 997268
rect 263919 996588 263985 996591
rect 507855 996588 507921 996591
rect 510255 996588 510321 996591
rect 263919 996586 264096 996588
rect 263919 996530 263924 996586
rect 263980 996530 264096 996586
rect 263919 996528 264096 996530
rect 507360 996586 507921 996588
rect 507360 996530 507860 996586
rect 507916 996530 507921 996586
rect 507360 996528 507921 996530
rect 509664 996586 510321 996588
rect 509664 996530 510260 996586
rect 510316 996530 510321 996586
rect 509664 996528 510321 996530
rect 263919 996525 263985 996528
rect 507855 996525 507921 996528
rect 510255 996525 510321 996528
rect 92559 996144 92625 996147
rect 164079 996144 164145 996147
rect 84546 996142 92625 996144
rect 84546 996086 92564 996142
rect 92620 996086 92625 996142
rect 84546 996084 92625 996086
rect 163680 996142 164145 996144
rect 163680 996086 164084 996142
rect 164140 996086 164145 996142
rect 163680 996084 164145 996086
rect 78639 995848 78705 995851
rect 84546 995848 84606 996084
rect 92559 996081 92625 996084
rect 164079 996081 164145 996084
rect 213327 996144 213393 996147
rect 215631 996144 215697 996147
rect 265071 996144 265137 996147
rect 266991 996144 267057 996147
rect 213327 996142 213504 996144
rect 213327 996086 213332 996142
rect 213388 996086 213504 996142
rect 213327 996084 213504 996086
rect 215631 996142 215808 996144
rect 215631 996086 215636 996142
rect 215692 996086 215808 996142
rect 215631 996084 215808 996086
rect 264864 996142 265137 996144
rect 264864 996086 265076 996142
rect 265132 996086 265137 996142
rect 264864 996084 265137 996086
rect 266400 996142 267057 996144
rect 266400 996086 266996 996142
rect 267052 996086 267057 996142
rect 266400 996084 267057 996086
rect 213327 996081 213393 996084
rect 215631 996081 215697 996084
rect 265071 996081 265137 996084
rect 266991 996081 267057 996084
rect 316335 996144 316401 996147
rect 318639 996144 318705 996147
rect 367119 996144 367185 996147
rect 316335 996142 316512 996144
rect 316335 996086 316340 996142
rect 316396 996086 316512 996142
rect 316335 996084 316512 996086
rect 318639 996142 318816 996144
rect 318639 996086 318644 996142
rect 318700 996086 318816 996142
rect 318639 996084 318816 996086
rect 366912 996142 367185 996144
rect 366912 996086 367124 996142
rect 367180 996086 367185 996142
rect 366912 996084 367185 996086
rect 316335 996081 316401 996084
rect 318639 996081 318705 996084
rect 367119 996081 367185 996084
rect 380271 996144 380337 996147
rect 385978 996144 385984 996146
rect 380271 996142 385984 996144
rect 380271 996086 380276 996142
rect 380332 996086 385984 996142
rect 380271 996084 385984 996086
rect 380271 996081 380337 996084
rect 385978 996082 385984 996084
rect 386048 996082 386054 996146
rect 436431 996144 436497 996147
rect 435840 996142 436497 996144
rect 435840 996086 436436 996142
rect 436492 996086 436497 996142
rect 435840 996084 436497 996086
rect 436431 996081 436497 996084
rect 511119 996144 511185 996147
rect 513423 996144 513489 996147
rect 511119 996142 511296 996144
rect 511119 996086 511124 996142
rect 511180 996086 511296 996142
rect 511119 996084 511296 996086
rect 513423 996142 513696 996144
rect 513423 996086 513428 996142
rect 513484 996086 513696 996142
rect 513423 996084 513696 996086
rect 511119 996081 511185 996084
rect 513423 996081 513489 996084
rect 101487 995996 101553 995999
rect 103887 995996 103953 995999
rect 106959 995996 107025 995999
rect 113391 995996 113457 995999
rect 144207 995996 144273 995999
rect 101487 995994 102048 995996
rect 101487 995938 101492 995994
rect 101548 995938 102048 995994
rect 101487 995936 102048 995938
rect 103887 995994 104352 995996
rect 103887 995938 103892 995994
rect 103948 995938 104352 995994
rect 103887 995936 104352 995938
rect 106959 995994 107424 995996
rect 106959 995938 106964 995994
rect 107020 995938 107424 995994
rect 106959 995936 107424 995938
rect 113391 995994 113856 995996
rect 113391 995938 113396 995994
rect 113452 995938 113856 995994
rect 113391 995936 113856 995938
rect 136770 995994 144273 995996
rect 136770 995938 144212 995994
rect 144268 995938 144273 995994
rect 136770 995936 144273 995938
rect 101487 995933 101553 995936
rect 103887 995933 103953 995936
rect 106959 995933 107025 995936
rect 113391 995933 113457 995936
rect 136770 995851 136830 995936
rect 144207 995933 144273 995936
rect 145263 995996 145329 995999
rect 149103 995996 149169 995999
rect 145263 995994 149169 995996
rect 145263 995938 145268 995994
rect 145324 995938 149108 995994
rect 149164 995938 149169 995994
rect 145263 995936 149169 995938
rect 145263 995933 145329 995936
rect 149103 995933 149169 995936
rect 149487 995996 149553 995999
rect 151983 995996 152049 995999
rect 159471 995996 159537 995999
rect 164175 995996 164241 995999
rect 195375 995996 195441 995999
rect 200271 995996 200337 995999
rect 149487 995994 150144 995996
rect 149487 995938 149492 995994
rect 149548 995938 150144 995994
rect 149487 995936 150144 995938
rect 151983 995994 152544 995996
rect 151983 995938 151988 995994
rect 152044 995938 152544 995994
rect 151983 995936 152544 995938
rect 159471 995994 159648 995996
rect 159471 995938 159476 995994
rect 159532 995938 159648 995994
rect 159471 995936 159648 995938
rect 164175 995994 164448 995996
rect 164175 995938 164180 995994
rect 164236 995938 164448 995994
rect 164175 995936 164448 995938
rect 192258 995994 195441 995996
rect 192258 995938 195380 995994
rect 195436 995938 195441 995994
rect 192258 995936 195441 995938
rect 200064 995994 200337 995996
rect 200064 995938 200276 995994
rect 200332 995938 200337 995994
rect 200064 995936 200337 995938
rect 149487 995933 149553 995936
rect 151983 995933 152049 995936
rect 159471 995933 159537 995936
rect 164175 995933 164241 995936
rect 95055 995848 95121 995851
rect 78639 995846 84606 995848
rect 78639 995790 78644 995846
rect 78700 995790 84606 995846
rect 78639 995788 84606 995790
rect 94722 995846 95121 995848
rect 94722 995790 95060 995846
rect 95116 995790 95121 995846
rect 99759 995848 99825 995851
rect 105423 995848 105489 995851
rect 113391 995848 113457 995851
rect 99759 995846 100416 995848
rect 94722 995788 95121 995790
rect 78639 995785 78705 995788
rect 89679 995700 89745 995703
rect 94722 995700 94782 995788
rect 95055 995785 95121 995788
rect 89679 995698 94782 995700
rect 89679 995642 89684 995698
rect 89740 995642 94782 995698
rect 89679 995640 94782 995642
rect 94959 995700 95025 995703
rect 97218 995700 97278 995818
rect 98754 995700 98814 995818
rect 94959 995698 98814 995700
rect 94959 995642 94964 995698
rect 95020 995642 98814 995698
rect 94959 995640 98814 995642
rect 98895 995700 98961 995703
rect 99522 995700 99582 995818
rect 99759 995790 99764 995846
rect 99820 995790 100416 995846
rect 105423 995846 105984 995848
rect 99759 995788 100416 995790
rect 99759 995785 99825 995788
rect 98895 995698 99582 995700
rect 98895 995642 98900 995698
rect 98956 995642 99582 995698
rect 98895 995640 99582 995642
rect 99663 995700 99729 995703
rect 101154 995700 101214 995818
rect 99663 995698 101214 995700
rect 99663 995642 99668 995698
rect 99724 995642 101214 995698
rect 99663 995640 101214 995642
rect 89679 995637 89745 995640
rect 94959 995637 95025 995640
rect 98895 995637 98961 995640
rect 99663 995637 99729 995640
rect 86511 995404 86577 995407
rect 98895 995404 98961 995407
rect 86511 995402 98961 995404
rect 86511 995346 86516 995402
rect 86572 995346 98900 995402
rect 98956 995346 98961 995402
rect 86511 995344 98961 995346
rect 86511 995341 86577 995344
rect 98895 995341 98961 995344
rect 87855 995256 87921 995259
rect 102690 995256 102750 995818
rect 103119 995700 103185 995703
rect 103458 995700 103518 995818
rect 103119 995698 103518 995700
rect 103119 995642 103124 995698
rect 103180 995642 103518 995698
rect 103119 995640 103518 995642
rect 103119 995637 103185 995640
rect 87855 995254 102750 995256
rect 87855 995198 87860 995254
rect 87916 995198 102750 995254
rect 87855 995196 102750 995198
rect 87855 995193 87921 995196
rect 100719 995108 100785 995111
rect 105090 995108 105150 995818
rect 105423 995790 105428 995846
rect 105484 995790 105984 995846
rect 105423 995788 105984 995790
rect 105423 995785 105489 995788
rect 108258 995555 108318 995818
rect 110688 995788 111294 995848
rect 112992 995846 113457 995848
rect 108207 995550 108318 995555
rect 108207 995494 108212 995550
rect 108268 995494 108318 995550
rect 108207 995492 108318 995494
rect 108207 995489 108273 995492
rect 111234 995404 111294 995788
rect 111522 995552 111582 995818
rect 112194 995700 112254 995818
rect 112992 995790 113396 995846
rect 113452 995790 113457 995846
rect 112992 995788 113457 995790
rect 113391 995785 113457 995788
rect 123855 995848 123921 995851
rect 134511 995848 134577 995851
rect 123855 995846 134577 995848
rect 123855 995790 123860 995846
rect 123916 995790 134516 995846
rect 134572 995790 134577 995846
rect 123855 995788 134577 995790
rect 123855 995785 123921 995788
rect 134511 995785 134577 995788
rect 136719 995846 136830 995851
rect 136719 995790 136724 995846
rect 136780 995790 136830 995846
rect 136719 995788 136830 995790
rect 137967 995848 138033 995851
rect 144015 995848 144081 995851
rect 137967 995846 144081 995848
rect 137967 995790 137972 995846
rect 138028 995790 144020 995846
rect 144076 995790 144081 995846
rect 158607 995848 158673 995851
rect 165615 995848 165681 995851
rect 166191 995848 166257 995851
rect 178479 995848 178545 995851
rect 185199 995848 185265 995851
rect 158607 995846 158880 995848
rect 137967 995788 144081 995790
rect 136719 995785 136785 995788
rect 137967 995785 138033 995788
rect 144015 995785 144081 995788
rect 115215 995700 115281 995703
rect 112194 995698 115281 995700
rect 112194 995642 115220 995698
rect 115276 995642 115281 995698
rect 112194 995640 115281 995642
rect 115215 995637 115281 995640
rect 137391 995700 137457 995703
rect 143631 995700 143697 995703
rect 137391 995698 143697 995700
rect 137391 995642 137396 995698
rect 137452 995642 143636 995698
rect 143692 995642 143697 995698
rect 137391 995640 143697 995642
rect 137391 995637 137457 995640
rect 143631 995637 143697 995640
rect 146799 995700 146865 995703
rect 154914 995700 154974 995818
rect 146799 995698 154974 995700
rect 146799 995642 146804 995698
rect 146860 995642 154974 995698
rect 146799 995640 154974 995642
rect 146799 995637 146865 995640
rect 115311 995552 115377 995555
rect 111522 995550 115377 995552
rect 111522 995494 115316 995550
rect 115372 995494 115377 995550
rect 111522 995492 115377 995494
rect 115311 995489 115377 995492
rect 146799 995552 146865 995555
rect 156546 995552 156606 995818
rect 146799 995550 156606 995552
rect 146799 995494 146804 995550
rect 146860 995494 156606 995550
rect 146799 995492 156606 995494
rect 146799 995489 146865 995492
rect 115215 995404 115281 995407
rect 111234 995402 115281 995404
rect 111234 995346 115220 995402
rect 115276 995346 115281 995402
rect 111234 995344 115281 995346
rect 115215 995341 115281 995344
rect 100719 995106 105150 995108
rect 100719 995050 100724 995106
rect 100780 995050 105150 995106
rect 100719 995048 105150 995050
rect 100719 995045 100785 995048
rect 136143 994368 136209 994371
rect 158178 994368 158238 995818
rect 158607 995790 158612 995846
rect 158668 995790 158880 995846
rect 158607 995788 158880 995790
rect 158607 995785 158673 995788
rect 158319 995700 158385 995703
rect 161250 995700 161310 995818
rect 158319 995698 161310 995700
rect 158319 995642 158324 995698
rect 158380 995642 161310 995698
rect 158319 995640 161310 995642
rect 158319 995637 158385 995640
rect 162114 995552 162174 995818
rect 162882 995703 162942 995818
rect 165216 995788 165438 995848
rect 162882 995698 162993 995703
rect 162882 995642 162932 995698
rect 162988 995642 162993 995698
rect 162882 995640 162993 995642
rect 165378 995700 165438 995788
rect 165615 995846 166080 995848
rect 165615 995790 165620 995846
rect 165676 995790 166080 995846
rect 165615 995788 166080 995790
rect 166191 995846 166944 995848
rect 166191 995790 166196 995846
rect 166252 995790 166944 995846
rect 166191 995788 166944 995790
rect 178479 995846 185265 995848
rect 178479 995790 178484 995846
rect 178540 995790 185204 995846
rect 185260 995790 185265 995846
rect 178479 995788 185265 995790
rect 165615 995785 165681 995788
rect 166191 995785 166257 995788
rect 178479 995785 178545 995788
rect 185199 995785 185265 995788
rect 187599 995848 187665 995851
rect 192258 995848 192318 995936
rect 195375 995933 195441 995936
rect 200271 995933 200337 995936
rect 200943 995996 201009 995999
rect 204207 995996 204273 995999
rect 206607 995996 206673 995999
rect 216783 995996 216849 995999
rect 246639 995996 246705 995999
rect 200943 995994 201504 995996
rect 200943 995938 200948 995994
rect 201004 995938 201504 995994
rect 200943 995936 201504 995938
rect 204207 995994 204768 995996
rect 204207 995938 204212 995994
rect 204268 995938 204768 995994
rect 204207 995936 204768 995938
rect 206607 995994 207072 995996
rect 206607 995938 206612 995994
rect 206668 995938 207072 995994
rect 206607 995936 207072 995938
rect 216783 995994 217440 995996
rect 216783 995938 216788 995994
rect 216844 995938 217440 995994
rect 216783 995936 217440 995938
rect 239298 995994 246705 995996
rect 239298 995938 246644 995994
rect 246700 995938 246705 995994
rect 239298 995936 246705 995938
rect 200943 995933 201009 995936
rect 204207 995933 204273 995936
rect 206607 995933 206673 995936
rect 216783 995933 216849 995936
rect 187599 995846 192318 995848
rect 187599 995790 187604 995846
rect 187660 995790 192318 995846
rect 187599 995788 192318 995790
rect 192495 995848 192561 995851
rect 195279 995848 195345 995851
rect 192495 995846 195345 995848
rect 192495 995790 192500 995846
rect 192556 995790 195284 995846
rect 195340 995790 195345 995846
rect 202863 995848 202929 995851
rect 203343 995848 203409 995851
rect 238863 995848 238929 995851
rect 239298 995848 239358 995936
rect 246639 995933 246705 995936
rect 247599 995996 247665 995999
rect 266895 995996 266961 995999
rect 305679 995996 305745 995999
rect 313839 995996 313905 995999
rect 326799 995996 326865 995999
rect 362319 995996 362385 995999
rect 370191 995996 370257 995999
rect 377487 995996 377553 995999
rect 429711 995996 429777 995999
rect 247599 995994 251424 995996
rect 247599 995938 247604 995994
rect 247660 995966 251424 995994
rect 266895 995994 267264 995996
rect 247660 995938 251454 995966
rect 247599 995936 251454 995938
rect 247599 995933 247665 995936
rect 202863 995846 203232 995848
rect 192495 995788 195345 995790
rect 187599 995785 187665 995788
rect 192495 995785 192561 995788
rect 195279 995785 195345 995788
rect 170223 995700 170289 995703
rect 165378 995698 170289 995700
rect 165378 995642 170228 995698
rect 170284 995642 170289 995698
rect 165378 995640 170289 995642
rect 162927 995637 162993 995640
rect 170223 995637 170289 995640
rect 189423 995700 189489 995703
rect 202338 995700 202398 995818
rect 202863 995790 202868 995846
rect 202924 995790 203232 995846
rect 202863 995788 203232 995790
rect 203343 995846 204000 995848
rect 203343 995790 203348 995846
rect 203404 995790 204000 995846
rect 203343 995788 204000 995790
rect 205314 995788 205536 995848
rect 238863 995846 239358 995848
rect 202863 995785 202929 995788
rect 203343 995785 203409 995788
rect 205314 995700 205374 995788
rect 189423 995698 202398 995700
rect 189423 995642 189428 995698
rect 189484 995642 202398 995698
rect 189423 995640 202398 995642
rect 202626 995640 205374 995700
rect 189423 995637 189489 995640
rect 162639 995552 162705 995555
rect 162114 995550 162705 995552
rect 162114 995494 162644 995550
rect 162700 995494 162705 995550
rect 162114 995492 162705 995494
rect 162639 995489 162705 995492
rect 185103 995552 185169 995555
rect 190575 995552 190641 995555
rect 202626 995552 202686 995640
rect 185103 995550 190398 995552
rect 185103 995494 185108 995550
rect 185164 995494 190398 995550
rect 185103 995492 190398 995494
rect 185103 995489 185169 995492
rect 190338 995404 190398 995492
rect 190575 995550 202686 995552
rect 190575 995494 190580 995550
rect 190636 995494 202686 995550
rect 190575 995492 202686 995494
rect 190575 995489 190641 995492
rect 203343 995404 203409 995407
rect 190338 995402 203409 995404
rect 190338 995346 203348 995402
rect 203404 995346 203409 995402
rect 190338 995344 203409 995346
rect 203343 995341 203409 995344
rect 201519 995256 201585 995259
rect 206274 995256 206334 995818
rect 210210 995259 210270 995818
rect 211074 995259 211134 995818
rect 212706 995407 212766 995818
rect 212655 995402 212766 995407
rect 212655 995346 212660 995402
rect 212716 995346 212766 995402
rect 212655 995344 212766 995346
rect 214338 995407 214398 995818
rect 215010 995700 215070 995818
rect 238863 995790 238868 995846
rect 238924 995790 239358 995846
rect 238863 995788 239358 995790
rect 239535 995848 239601 995851
rect 250479 995848 250545 995851
rect 239535 995846 250545 995848
rect 239535 995790 239540 995846
rect 239596 995790 250484 995846
rect 250540 995790 250545 995846
rect 251394 995848 251454 995936
rect 266895 995938 266900 995994
rect 266956 995938 267264 995994
rect 266895 995936 267264 995938
rect 305679 995994 306144 995996
rect 305679 995938 305684 995994
rect 305740 995938 306144 995994
rect 305679 995936 306144 995938
rect 313839 995994 314016 995996
rect 313839 995938 313844 995994
rect 313900 995938 314016 995994
rect 313839 995936 314016 995938
rect 321312 995994 326865 995996
rect 321312 995938 326804 995994
rect 326860 995938 326865 995994
rect 321312 995936 326865 995938
rect 362208 995994 362385 995996
rect 362208 995938 362324 995994
rect 362380 995938 362385 995994
rect 362208 995936 362385 995938
rect 370080 995994 370257 995996
rect 370080 995938 370196 995994
rect 370252 995938 370257 995994
rect 370080 995936 370257 995938
rect 371712 995994 377553 995996
rect 371712 995938 377492 995994
rect 377548 995938 377553 995994
rect 371712 995936 377553 995938
rect 266895 995933 266961 995936
rect 305679 995933 305745 995936
rect 313839 995933 313905 995936
rect 326799 995933 326865 995936
rect 362319 995933 362385 995936
rect 370191 995933 370257 995936
rect 377487 995933 377553 995936
rect 378498 995936 392958 995996
rect 429600 995994 429777 995996
rect 429600 995938 429716 995994
rect 429772 995938 429777 995994
rect 429600 995936 429777 995938
rect 254031 995848 254097 995851
rect 254895 995848 254961 995851
rect 255663 995848 255729 995851
rect 257295 995848 257361 995851
rect 262671 995848 262737 995851
rect 268527 995848 268593 995851
rect 273615 995848 273681 995851
rect 251394 995818 251838 995848
rect 239535 995788 250545 995790
rect 251424 995788 251838 995818
rect 238863 995785 238929 995788
rect 239535 995785 239601 995788
rect 250479 995785 250545 995788
rect 218895 995700 218961 995703
rect 215010 995698 218961 995700
rect 215010 995642 218900 995698
rect 218956 995642 218961 995698
rect 215010 995640 218961 995642
rect 218895 995637 218961 995640
rect 240207 995700 240273 995703
rect 250383 995700 250449 995703
rect 240207 995698 250449 995700
rect 240207 995642 240212 995698
rect 240268 995642 250388 995698
rect 250444 995642 250449 995698
rect 240207 995640 250449 995642
rect 251778 995700 251838 995788
rect 252930 995700 252990 995818
rect 253728 995788 253950 995848
rect 253890 995700 253950 995788
rect 254031 995846 254592 995848
rect 254031 995790 254036 995846
rect 254092 995790 254592 995846
rect 254031 995788 254592 995790
rect 254895 995846 255456 995848
rect 254895 995790 254900 995846
rect 254956 995790 255456 995846
rect 254895 995788 255456 995790
rect 255663 995846 256224 995848
rect 255663 995790 255668 995846
rect 255724 995790 256224 995846
rect 257295 995846 257760 995848
rect 255663 995788 256224 995790
rect 254031 995785 254097 995788
rect 254895 995785 254961 995788
rect 255663 995785 255729 995788
rect 251778 995640 252990 995700
rect 253698 995640 253950 995700
rect 240207 995637 240273 995640
rect 250383 995637 250449 995640
rect 240783 995552 240849 995555
rect 253698 995552 253758 995640
rect 240783 995550 253758 995552
rect 240783 995494 240788 995550
rect 240844 995494 253758 995550
rect 240783 995492 253758 995494
rect 240783 995489 240849 995492
rect 214338 995402 214449 995407
rect 214338 995346 214388 995402
rect 214444 995346 214449 995402
rect 214338 995344 214449 995346
rect 212655 995341 212721 995344
rect 214383 995341 214449 995344
rect 241839 995404 241905 995407
rect 256866 995404 256926 995818
rect 257295 995790 257300 995846
rect 257356 995790 257760 995846
rect 257295 995788 257760 995790
rect 257295 995785 257361 995788
rect 241839 995402 256926 995404
rect 241839 995346 241844 995402
rect 241900 995346 256926 995402
rect 241839 995344 256926 995346
rect 241839 995341 241905 995344
rect 201519 995254 206334 995256
rect 201519 995198 201524 995254
rect 201580 995198 206334 995254
rect 201519 995196 206334 995198
rect 210159 995254 210270 995259
rect 210159 995198 210164 995254
rect 210220 995198 210270 995254
rect 210159 995196 210270 995198
rect 211023 995254 211134 995259
rect 211023 995198 211028 995254
rect 211084 995198 211134 995254
rect 211023 995196 211134 995198
rect 201519 995193 201585 995196
rect 210159 995193 210225 995196
rect 211023 995193 211089 995196
rect 250479 995108 250545 995111
rect 258498 995108 258558 995818
rect 261600 995788 261822 995848
rect 262671 995846 263328 995848
rect 261762 995700 261822 995788
rect 250479 995106 258558 995108
rect 250479 995050 250484 995106
rect 250540 995050 258558 995106
rect 250479 995048 258558 995050
rect 261570 995640 261822 995700
rect 250479 995045 250545 995048
rect 261570 994960 261630 995640
rect 238722 994900 261630 994960
rect 234351 994516 234417 994519
rect 238722 994516 238782 994900
rect 262434 994812 262494 995818
rect 262671 995790 262676 995846
rect 262732 995790 263328 995846
rect 268032 995846 268593 995848
rect 262671 995788 263328 995790
rect 262671 995785 262737 995788
rect 265698 995703 265758 995818
rect 268032 995790 268532 995846
rect 268588 995790 268593 995846
rect 269664 995846 273681 995848
rect 268032 995788 268593 995790
rect 268527 995785 268593 995788
rect 265698 995698 265809 995703
rect 265698 995642 265748 995698
rect 265804 995642 265809 995698
rect 265698 995640 265809 995642
rect 265743 995637 265809 995640
rect 268047 995700 268113 995703
rect 268866 995700 268926 995818
rect 269664 995790 273620 995846
rect 273676 995790 273681 995846
rect 269664 995788 273681 995790
rect 273615 995785 273681 995788
rect 292527 995848 292593 995851
rect 299439 995848 299505 995851
rect 304719 995848 304785 995851
rect 307311 995848 307377 995851
rect 310287 995848 310353 995851
rect 317487 995848 317553 995851
rect 292527 995846 299505 995848
rect 292527 995790 292532 995846
rect 292588 995790 299444 995846
rect 299500 995790 299505 995846
rect 292527 995788 299505 995790
rect 292527 995785 292593 995788
rect 299439 995785 299505 995788
rect 268047 995698 268926 995700
rect 268047 995642 268052 995698
rect 268108 995642 268926 995698
rect 268047 995640 268926 995642
rect 295407 995700 295473 995703
rect 298191 995700 298257 995703
rect 295407 995698 298257 995700
rect 295407 995642 295412 995698
rect 295468 995642 298196 995698
rect 298252 995642 298257 995698
rect 295407 995640 298257 995642
rect 268047 995637 268113 995640
rect 295407 995637 295473 995640
rect 298191 995637 298257 995640
rect 298479 995700 298545 995703
rect 303042 995700 303102 995818
rect 304002 995788 304608 995848
rect 304719 995846 305376 995848
rect 304719 995790 304724 995846
rect 304780 995790 305376 995846
rect 307311 995846 307872 995848
rect 304719 995788 305376 995790
rect 304002 995700 304062 995788
rect 304719 995785 304785 995788
rect 298479 995698 304062 995700
rect 298479 995642 298484 995698
rect 298540 995642 304062 995698
rect 298479 995640 304062 995642
rect 298479 995637 298545 995640
rect 286767 995552 286833 995555
rect 299535 995552 299601 995555
rect 286767 995550 299601 995552
rect 286767 995494 286772 995550
rect 286828 995494 299540 995550
rect 299596 995494 299601 995550
rect 286767 995492 299601 995494
rect 286767 995489 286833 995492
rect 299535 995489 299601 995492
rect 302319 995552 302385 995555
rect 306978 995552 307038 995818
rect 307311 995790 307316 995846
rect 307372 995790 307872 995846
rect 307311 995788 307872 995790
rect 308448 995788 308670 995848
rect 307311 995785 307377 995788
rect 308610 995700 308670 995788
rect 310287 995846 310944 995848
rect 310287 995790 310292 995846
rect 310348 995790 310944 995846
rect 310287 995788 310944 995790
rect 310287 995785 310353 995788
rect 302319 995550 307038 995552
rect 302319 995494 302324 995550
rect 302380 995494 307038 995550
rect 302319 995492 307038 995494
rect 308418 995640 308670 995700
rect 309231 995700 309297 995703
rect 312546 995700 312606 995818
rect 309231 995698 312606 995700
rect 309231 995642 309236 995698
rect 309292 995642 312606 995698
rect 309231 995640 312606 995642
rect 302319 995489 302385 995492
rect 293583 995404 293649 995407
rect 308418 995404 308478 995640
rect 309231 995637 309297 995640
rect 293583 995402 308478 995404
rect 293583 995346 293588 995402
rect 293644 995346 308478 995402
rect 293583 995344 308478 995346
rect 293583 995341 293649 995344
rect 290319 994812 290385 994815
rect 309231 994812 309297 994815
rect 262434 994752 262974 994812
rect 243567 994664 243633 994667
rect 262671 994664 262737 994667
rect 243567 994662 262737 994664
rect 243567 994606 243572 994662
rect 243628 994606 262676 994662
rect 262732 994606 262737 994662
rect 243567 994604 262737 994606
rect 243567 994601 243633 994604
rect 262671 994601 262737 994604
rect 234351 994514 238782 994516
rect 234351 994458 234356 994514
rect 234412 994458 238782 994514
rect 234351 994456 238782 994458
rect 234351 994453 234417 994456
rect 136143 994366 158238 994368
rect 136143 994310 136148 994366
rect 136204 994310 158238 994366
rect 136143 994308 158238 994310
rect 231471 994368 231537 994371
rect 262914 994368 262974 994752
rect 290319 994810 309297 994812
rect 290319 994754 290324 994810
rect 290380 994754 309236 994810
rect 309292 994754 309297 994810
rect 290319 994752 309297 994754
rect 290319 994749 290385 994752
rect 309231 994749 309297 994752
rect 286287 994664 286353 994667
rect 313218 994664 313278 995818
rect 315138 995788 315744 995848
rect 317280 995846 317553 995848
rect 317280 995790 317492 995846
rect 317548 995790 317553 995846
rect 350127 995848 350193 995851
rect 360975 995848 361041 995851
rect 365871 995848 365937 995851
rect 377295 995848 377361 995851
rect 378498 995848 378558 995936
rect 350127 995846 353472 995848
rect 317280 995788 317553 995790
rect 313359 995700 313425 995703
rect 315138 995700 315198 995788
rect 317487 995785 317553 995788
rect 313359 995698 315198 995700
rect 313359 995642 313364 995698
rect 313420 995642 315198 995698
rect 313359 995640 315198 995642
rect 319650 995700 319710 995818
rect 350127 995790 350132 995846
rect 350188 995818 353472 995846
rect 350188 995790 353502 995818
rect 350127 995788 353502 995790
rect 354912 995788 355134 995848
rect 360480 995846 361041 995848
rect 360480 995790 360980 995846
rect 361036 995790 361041 995846
rect 365280 995846 365937 995848
rect 360480 995788 361041 995790
rect 350127 995785 350193 995788
rect 323919 995700 323985 995703
rect 319650 995698 323985 995700
rect 319650 995642 323924 995698
rect 323980 995642 323985 995698
rect 319650 995640 323985 995642
rect 353442 995700 353502 995788
rect 355074 995700 355134 995788
rect 360975 995785 361041 995788
rect 353442 995640 355134 995700
rect 313359 995637 313425 995640
rect 323919 995637 323985 995640
rect 362946 995256 363006 995818
rect 363618 995404 363678 995818
rect 365280 995790 365876 995846
rect 365932 995790 365937 995846
rect 365280 995788 365937 995790
rect 366048 995788 366654 995848
rect 377295 995846 378558 995848
rect 365871 995785 365937 995788
rect 366594 995552 366654 995788
rect 368418 995700 368478 995818
rect 368847 995700 368913 995703
rect 368418 995698 368913 995700
rect 368418 995642 368852 995698
rect 368908 995642 368913 995698
rect 368418 995640 368913 995642
rect 370818 995700 370878 995818
rect 377295 995790 377300 995846
rect 377356 995790 378558 995846
rect 377295 995788 378558 995790
rect 380175 995848 380241 995851
rect 388815 995848 388881 995851
rect 380175 995846 388881 995848
rect 380175 995790 380180 995846
rect 380236 995790 388820 995846
rect 388876 995790 388881 995846
rect 380175 995788 388881 995790
rect 392898 995848 392958 995936
rect 429711 995933 429777 995936
rect 436431 995996 436497 995999
rect 472047 995996 472113 995999
rect 511887 995996 511953 995999
rect 513423 995996 513489 995999
rect 521391 995996 521457 995999
rect 436431 995994 436608 995996
rect 436431 995938 436436 995994
rect 436492 995938 436608 995994
rect 436431 995936 436608 995938
rect 472047 995994 478206 995996
rect 472047 995938 472052 995994
rect 472108 995938 478206 995994
rect 472047 995936 478206 995938
rect 436431 995933 436497 995936
rect 472047 995933 472113 995936
rect 396687 995848 396753 995851
rect 466479 995848 466545 995851
rect 477039 995848 477105 995851
rect 392898 995846 396753 995848
rect 392898 995790 396692 995846
rect 396748 995790 396753 995846
rect 392898 995788 396753 995790
rect 377295 995785 377361 995788
rect 380175 995785 380241 995788
rect 388815 995785 388881 995788
rect 396687 995785 396753 995788
rect 374415 995700 374481 995703
rect 370818 995698 374481 995700
rect 370818 995642 374420 995698
rect 374476 995642 374481 995698
rect 370818 995640 374481 995642
rect 368847 995637 368913 995640
rect 374415 995637 374481 995640
rect 381423 995700 381489 995703
rect 393039 995700 393105 995703
rect 381423 995698 393105 995700
rect 381423 995642 381428 995698
rect 381484 995642 393044 995698
rect 393100 995642 393105 995698
rect 381423 995640 393105 995642
rect 381423 995637 381489 995640
rect 393039 995637 393105 995640
rect 410319 995700 410385 995703
rect 420834 995700 420894 995818
rect 422304 995788 422526 995848
rect 466479 995846 477105 995848
rect 422466 995700 422526 995788
rect 410319 995698 422526 995700
rect 410319 995642 410324 995698
rect 410380 995642 422526 995698
rect 410319 995640 422526 995642
rect 437442 995700 437502 995818
rect 466479 995790 466484 995846
rect 466540 995790 477044 995846
rect 477100 995790 477105 995846
rect 466479 995788 477105 995790
rect 478146 995848 478206 995936
rect 511887 995994 512160 995996
rect 511887 995938 511892 995994
rect 511948 995938 512160 995994
rect 511887 995936 512160 995938
rect 512832 995994 513489 995996
rect 512832 995938 513428 995994
rect 513484 995938 513489 995994
rect 512832 995936 513489 995938
rect 516096 995994 521457 995996
rect 516096 995938 521396 995994
rect 521452 995938 521457 995994
rect 516096 995936 521457 995938
rect 511887 995933 511953 995936
rect 513423 995933 513489 995936
rect 521391 995933 521457 995936
rect 564783 995996 564849 995999
rect 564783 995994 565056 995996
rect 564783 995938 564788 995994
rect 564844 995938 565056 995994
rect 564783 995936 565056 995938
rect 564783 995933 564849 995936
rect 481455 995848 481521 995851
rect 519471 995848 519537 995851
rect 532815 995848 532881 995851
rect 563727 995848 563793 995851
rect 573135 995848 573201 995851
rect 478146 995846 481521 995848
rect 478146 995790 481460 995846
rect 481516 995790 481521 995846
rect 478146 995788 481521 995790
rect 466479 995785 466545 995788
rect 477039 995785 477105 995788
rect 481455 995785 481521 995788
rect 440655 995700 440721 995703
rect 437442 995698 440721 995700
rect 437442 995642 440660 995698
rect 440716 995642 440721 995698
rect 437442 995640 440721 995642
rect 410319 995637 410385 995640
rect 440655 995637 440721 995640
rect 480111 995700 480177 995703
rect 488847 995700 488913 995703
rect 480111 995698 488913 995700
rect 480111 995642 480116 995698
rect 480172 995642 488852 995698
rect 488908 995642 488913 995698
rect 480111 995640 488913 995642
rect 480111 995637 480177 995640
rect 488847 995637 488913 995640
rect 385839 995552 385905 995555
rect 366594 995550 385905 995552
rect 366594 995494 385844 995550
rect 385900 995494 385905 995550
rect 366594 995492 385905 995494
rect 385839 995489 385905 995492
rect 385978 995490 385984 995554
rect 386048 995552 386054 995554
rect 394863 995552 394929 995555
rect 386048 995550 394929 995552
rect 386048 995494 394868 995550
rect 394924 995494 394929 995550
rect 386048 995492 394929 995494
rect 386048 995490 386054 995492
rect 394863 995489 394929 995492
rect 506562 995407 506622 995818
rect 514434 995552 514494 995818
rect 515232 995788 515454 995848
rect 515394 995700 515454 995788
rect 519471 995846 532881 995848
rect 519471 995790 519476 995846
rect 519532 995790 532820 995846
rect 532876 995790 532881 995846
rect 563520 995846 563793 995848
rect 519471 995788 532881 995790
rect 519471 995785 519537 995788
rect 532815 995785 532881 995788
rect 518415 995700 518481 995703
rect 515394 995698 518481 995700
rect 515394 995642 518420 995698
rect 518476 995642 518481 995698
rect 515394 995640 518481 995642
rect 518415 995637 518481 995640
rect 521199 995700 521265 995703
rect 532239 995700 532305 995703
rect 521199 995698 532305 995700
rect 521199 995642 521204 995698
rect 521260 995642 532244 995698
rect 532300 995642 532305 995698
rect 521199 995640 532305 995642
rect 521199 995637 521265 995640
rect 532239 995637 532305 995640
rect 518511 995552 518577 995555
rect 514434 995550 518577 995552
rect 514434 995494 518516 995550
rect 518572 995494 518577 995550
rect 514434 995492 518577 995494
rect 518511 995489 518577 995492
rect 521007 995552 521073 995555
rect 534063 995552 534129 995555
rect 521007 995550 534129 995552
rect 521007 995494 521012 995550
rect 521068 995494 534068 995550
rect 534124 995494 534129 995550
rect 521007 995492 534129 995494
rect 521007 995489 521073 995492
rect 534063 995489 534129 995492
rect 557922 995407 557982 995818
rect 562722 995703 562782 995818
rect 563520 995790 563732 995846
rect 563788 995790 563793 995846
rect 567456 995846 573201 995848
rect 563520 995788 563793 995790
rect 563727 995785 563793 995788
rect 562722 995698 562833 995703
rect 562722 995642 562772 995698
rect 562828 995642 562833 995698
rect 562722 995640 562833 995642
rect 562767 995637 562833 995640
rect 565794 995552 565854 995818
rect 566658 995700 566718 995818
rect 567456 995790 573140 995846
rect 573196 995790 573201 995846
rect 567456 995788 573201 995790
rect 573135 995785 573201 995788
rect 570255 995700 570321 995703
rect 566658 995698 570321 995700
rect 566658 995642 570260 995698
rect 570316 995642 570321 995698
rect 566658 995640 570321 995642
rect 570255 995637 570321 995640
rect 570447 995552 570513 995555
rect 565794 995550 570513 995552
rect 565794 995494 570452 995550
rect 570508 995494 570513 995550
rect 565794 995492 570513 995494
rect 570447 995489 570513 995492
rect 387471 995404 387537 995407
rect 363618 995402 387537 995404
rect 363618 995346 387476 995402
rect 387532 995346 387537 995402
rect 363618 995344 387537 995346
rect 506562 995402 506673 995407
rect 506562 995346 506612 995402
rect 506668 995346 506673 995402
rect 506562 995344 506673 995346
rect 387471 995341 387537 995344
rect 506607 995341 506673 995344
rect 523407 995404 523473 995407
rect 530895 995404 530961 995407
rect 523407 995402 530961 995404
rect 523407 995346 523412 995402
rect 523468 995346 530900 995402
rect 530956 995346 530961 995402
rect 523407 995344 530961 995346
rect 557922 995402 558033 995407
rect 557922 995346 557972 995402
rect 558028 995346 558033 995402
rect 557922 995344 558033 995346
rect 523407 995341 523473 995344
rect 530895 995341 530961 995344
rect 557967 995341 558033 995344
rect 392079 995256 392145 995259
rect 362946 995254 392145 995256
rect 362946 995198 392084 995254
rect 392140 995198 392145 995254
rect 362946 995196 392145 995198
rect 392079 995193 392145 995196
rect 381999 995108 382065 995111
rect 392655 995108 392721 995111
rect 381999 995106 392721 995108
rect 381999 995050 382004 995106
rect 382060 995050 392660 995106
rect 392716 995050 392721 995106
rect 381999 995048 392721 995050
rect 381999 995045 382065 995048
rect 392655 995045 392721 995048
rect 379023 994960 379089 994963
rect 393711 994960 393777 994963
rect 379023 994958 393777 994960
rect 379023 994902 379028 994958
rect 379084 994902 393716 994958
rect 393772 994902 393777 994958
rect 379023 994900 393777 994902
rect 379023 994897 379089 994900
rect 393711 994897 393777 994900
rect 570831 994960 570897 994963
rect 629967 994960 630033 994963
rect 570831 994958 630033 994960
rect 570831 994902 570836 994958
rect 570892 994902 629972 994958
rect 630028 994902 630033 994958
rect 570831 994900 630033 994902
rect 570831 994897 570897 994900
rect 629967 994897 630033 994900
rect 570351 994812 570417 994815
rect 634287 994812 634353 994815
rect 570351 994810 634353 994812
rect 570351 994754 570356 994810
rect 570412 994754 634292 994810
rect 634348 994754 634353 994810
rect 570351 994752 634353 994754
rect 570351 994749 570417 994752
rect 634287 994749 634353 994752
rect 286287 994662 313278 994664
rect 286287 994606 286292 994662
rect 286348 994606 313278 994662
rect 286287 994604 313278 994606
rect 469551 994664 469617 994667
rect 485967 994664 486033 994667
rect 469551 994662 486033 994664
rect 469551 994606 469556 994662
rect 469612 994606 485972 994662
rect 486028 994606 486033 994662
rect 469551 994604 486033 994606
rect 286287 994601 286353 994604
rect 469551 994601 469617 994604
rect 485967 994601 486033 994604
rect 515535 994664 515601 994667
rect 533679 994664 533745 994667
rect 515535 994662 533745 994664
rect 515535 994606 515540 994662
rect 515596 994606 533684 994662
rect 533740 994606 533745 994662
rect 515535 994604 533745 994606
rect 515535 994601 515601 994604
rect 533679 994601 533745 994604
rect 571023 994664 571089 994667
rect 639183 994664 639249 994667
rect 571023 994662 639249 994664
rect 571023 994606 571028 994662
rect 571084 994606 639188 994662
rect 639244 994606 639249 994662
rect 571023 994604 639249 994606
rect 571023 994601 571089 994604
rect 639183 994601 639249 994604
rect 284367 994516 284433 994519
rect 313359 994516 313425 994519
rect 284367 994514 313425 994516
rect 284367 994458 284372 994514
rect 284428 994458 313364 994514
rect 313420 994458 313425 994514
rect 284367 994456 313425 994458
rect 284367 994453 284433 994456
rect 313359 994453 313425 994456
rect 365775 994516 365841 994519
rect 388335 994516 388401 994519
rect 391119 994516 391185 994519
rect 479823 994516 479889 994519
rect 365775 994514 388401 994516
rect 365775 994458 365780 994514
rect 365836 994458 388340 994514
rect 388396 994458 388401 994514
rect 365775 994456 388401 994458
rect 365775 994453 365841 994456
rect 388335 994453 388401 994456
rect 390978 994514 479889 994516
rect 390978 994458 391124 994514
rect 391180 994458 479828 994514
rect 479884 994458 479889 994514
rect 390978 994456 479889 994458
rect 390978 994368 391038 994456
rect 391119 994453 391185 994456
rect 479823 994453 479889 994456
rect 531183 994516 531249 994519
rect 630735 994516 630801 994519
rect 632751 994516 632817 994519
rect 531183 994514 632817 994516
rect 531183 994458 531188 994514
rect 531244 994458 630740 994514
rect 630796 994458 632756 994514
rect 632812 994458 632817 994514
rect 531183 994456 632817 994458
rect 531183 994453 531249 994456
rect 630735 994453 630801 994456
rect 632751 994453 632817 994456
rect 231471 994366 262974 994368
rect 231471 994310 231476 994366
rect 231532 994310 262974 994366
rect 231471 994308 262974 994310
rect 294402 994308 391038 994368
rect 396303 994368 396369 994371
rect 638511 994368 638577 994371
rect 396303 994366 638577 994368
rect 396303 994310 396308 994366
rect 396364 994310 638516 994366
rect 638572 994310 638577 994366
rect 396303 994308 638577 994310
rect 136143 994305 136209 994308
rect 231471 994305 231537 994308
rect 129711 994220 129777 994223
rect 158319 994220 158385 994223
rect 129711 994218 158385 994220
rect 129711 994162 129716 994218
rect 129772 994162 158324 994218
rect 158380 994162 158385 994218
rect 129711 994160 158385 994162
rect 129711 994157 129777 994160
rect 158319 994157 158385 994160
rect 185391 994220 185457 994223
rect 227535 994220 227601 994223
rect 288975 994220 289041 994223
rect 294402 994220 294462 994308
rect 396303 994305 396369 994308
rect 638511 994305 638577 994308
rect 185391 994218 227601 994220
rect 185391 994162 185396 994218
rect 185452 994162 227540 994218
rect 227596 994162 227601 994218
rect 185391 994160 227601 994162
rect 185391 994157 185457 994160
rect 227535 994157 227601 994160
rect 242946 994218 294462 994220
rect 242946 994162 288980 994218
rect 289036 994162 294462 994218
rect 242946 994160 294462 994162
rect 294543 994220 294609 994223
rect 640719 994220 640785 994223
rect 294543 994218 640785 994220
rect 294543 994162 294548 994218
rect 294604 994162 640724 994218
rect 640780 994162 640785 994218
rect 294543 994160 640785 994162
rect 134607 994072 134673 994075
rect 185967 994072 186033 994075
rect 237423 994072 237489 994075
rect 242946 994072 243006 994160
rect 288975 994157 289041 994160
rect 294543 994157 294609 994160
rect 640719 994157 640785 994160
rect 134607 994070 243006 994072
rect 134607 994014 134612 994070
rect 134668 994014 185972 994070
rect 186028 994014 237428 994070
rect 237484 994014 243006 994070
rect 134607 994012 243006 994014
rect 243183 994072 243249 994075
rect 650031 994072 650097 994075
rect 243183 994070 650097 994072
rect 243183 994014 243188 994070
rect 243244 994014 650036 994070
rect 650092 994014 650097 994070
rect 243183 994012 650097 994014
rect 134607 994009 134673 994012
rect 185967 994009 186033 994012
rect 237423 994009 237489 994012
rect 243183 994009 243249 994012
rect 650031 994009 650097 994012
rect 88719 993924 88785 993927
rect 576015 993924 576081 993927
rect 88719 993922 576081 993924
rect 88719 993866 88724 993922
rect 88780 993866 576020 993922
rect 576076 993866 576081 993922
rect 88719 993864 576081 993866
rect 88719 993861 88785 993864
rect 576015 993861 576081 993864
rect 80175 993776 80241 993779
rect 106959 993776 107025 993779
rect 80175 993774 107025 993776
rect 80175 993718 80180 993774
rect 80236 993718 106964 993774
rect 107020 993718 107025 993774
rect 80175 993716 107025 993718
rect 80175 993713 80241 993716
rect 106959 993713 107025 993716
rect 140367 993776 140433 993779
rect 633615 993776 633681 993779
rect 140367 993774 633681 993776
rect 140367 993718 140372 993774
rect 140428 993718 633620 993774
rect 633676 993718 633681 993774
rect 140367 993716 633681 993718
rect 140367 993713 140433 993716
rect 633615 993713 633681 993716
rect 62031 993628 62097 993631
rect 83439 993628 83505 993631
rect 92943 993628 93009 993631
rect 62031 993626 93009 993628
rect 62031 993570 62036 993626
rect 62092 993570 83444 993626
rect 83500 993570 92948 993626
rect 93004 993570 93009 993626
rect 62031 993568 93009 993570
rect 62031 993565 62097 993568
rect 83439 993565 83505 993568
rect 92943 993565 93009 993568
rect 279279 993628 279345 993631
rect 288399 993628 288465 993631
rect 294778 993628 294784 993630
rect 279279 993626 294784 993628
rect 279279 993570 279284 993626
rect 279340 993570 288404 993626
rect 288460 993570 294784 993626
rect 279279 993568 294784 993570
rect 279279 993565 279345 993568
rect 288399 993565 288465 993568
rect 294778 993566 294784 993568
rect 294848 993566 294854 993630
rect 390159 993628 390225 993631
rect 469455 993628 469521 993631
rect 390159 993626 469521 993628
rect 390159 993570 390164 993626
rect 390220 993570 469460 993626
rect 469516 993570 469521 993626
rect 390159 993568 469521 993570
rect 390159 993565 390225 993568
rect 469455 993565 469521 993568
rect 294778 992086 294784 992150
rect 294848 992148 294854 992150
rect 390159 992148 390225 992151
rect 294848 992146 390225 992148
rect 294848 992090 390164 992146
rect 390220 992090 390225 992146
rect 294848 992088 390225 992090
rect 294848 992086 294854 992088
rect 390159 992085 390225 992088
rect 181455 985488 181521 985491
rect 187311 985488 187377 985491
rect 181455 985486 187377 985488
rect 181455 985430 181460 985486
rect 181516 985430 187316 985486
rect 187372 985430 187377 985486
rect 181455 985428 187377 985430
rect 181455 985425 181521 985428
rect 187311 985425 187377 985428
rect 655119 974388 655185 974391
rect 650208 974386 655185 974388
rect 650208 974330 655124 974386
rect 655180 974330 655185 974386
rect 650208 974328 655185 974330
rect 655119 974325 655185 974328
rect 59535 973056 59601 973059
rect 59535 973054 64416 973056
rect 59535 972998 59540 973054
rect 59596 972998 64416 973054
rect 59535 972996 64416 972998
rect 59535 972993 59601 972996
rect 40570 968702 40576 968766
rect 40640 968764 40646 968766
rect 41775 968764 41841 968767
rect 40640 968762 41841 968764
rect 40640 968706 41780 968762
rect 41836 968706 41841 968762
rect 40640 968704 41841 968706
rect 40640 968702 40646 968704
rect 41775 968701 41841 968704
rect 673935 967580 674001 967583
rect 675514 967580 675520 967582
rect 673935 967578 675520 967580
rect 673935 967522 673940 967578
rect 673996 967522 675520 967578
rect 673935 967520 675520 967522
rect 673935 967517 674001 967520
rect 675514 967518 675520 967520
rect 675584 967518 675590 967582
rect 41775 967138 41841 967139
rect 41722 967136 41728 967138
rect 41684 967076 41728 967136
rect 41792 967134 41841 967138
rect 41836 967078 41841 967134
rect 41722 967074 41728 967076
rect 41792 967074 41841 967078
rect 41775 967073 41841 967074
rect 674554 965594 674560 965658
rect 674624 965656 674630 965658
rect 675087 965656 675153 965659
rect 674624 965654 675153 965656
rect 674624 965598 675092 965654
rect 675148 965598 675153 965654
rect 674624 965596 675153 965598
rect 674624 965594 674630 965596
rect 675087 965593 675153 965596
rect 675759 965656 675825 965659
rect 675898 965656 675904 965658
rect 675759 965654 675904 965656
rect 675759 965598 675764 965654
rect 675820 965598 675904 965654
rect 675759 965596 675904 965598
rect 675759 965593 675825 965596
rect 675898 965594 675904 965596
rect 675968 965594 675974 965658
rect 40378 965002 40384 965066
rect 40448 965064 40454 965066
rect 41775 965064 41841 965067
rect 40448 965062 41841 965064
rect 40448 965006 41780 965062
rect 41836 965006 41841 965062
rect 40448 965004 41841 965006
rect 40448 965002 40454 965004
rect 41775 965001 41841 965004
rect 674746 964854 674752 964918
rect 674816 964916 674822 964918
rect 675087 964916 675153 964919
rect 674816 964914 675153 964916
rect 674816 964858 675092 964914
rect 675148 964858 675153 964914
rect 674816 964856 675153 964858
rect 674816 964854 674822 964856
rect 675087 964853 675153 964856
rect 40762 963966 40768 964030
rect 40832 964028 40838 964030
rect 41775 964028 41841 964031
rect 40832 964026 41841 964028
rect 40832 963970 41780 964026
rect 41836 963970 41841 964026
rect 40832 963968 41841 963970
rect 40832 963966 40838 963968
rect 41775 963965 41841 963968
rect 40954 963374 40960 963438
rect 41024 963436 41030 963438
rect 41775 963436 41841 963439
rect 41024 963434 41841 963436
rect 41024 963378 41780 963434
rect 41836 963378 41841 963434
rect 41024 963376 41841 963378
rect 41024 963374 41030 963376
rect 41775 963373 41841 963376
rect 41146 962782 41152 962846
rect 41216 962844 41222 962846
rect 41775 962844 41841 962847
rect 41216 962842 41841 962844
rect 41216 962786 41780 962842
rect 41836 962786 41841 962842
rect 41216 962784 41841 962786
rect 41216 962782 41222 962784
rect 41775 962781 41841 962784
rect 674938 962782 674944 962846
rect 675008 962844 675014 962846
rect 675087 962844 675153 962847
rect 675008 962842 675153 962844
rect 675008 962786 675092 962842
rect 675148 962786 675153 962842
rect 675008 962784 675153 962786
rect 675008 962782 675014 962784
rect 675087 962781 675153 962784
rect 655215 962696 655281 962699
rect 650208 962694 655281 962696
rect 650208 962638 655220 962694
rect 655276 962638 655281 962694
rect 650208 962636 655281 962638
rect 655215 962633 655281 962636
rect 674362 962486 674368 962550
rect 674432 962548 674438 962550
rect 675183 962548 675249 962551
rect 674432 962546 675249 962548
rect 674432 962490 675188 962546
rect 675244 962490 675249 962546
rect 674432 962488 675249 962490
rect 674432 962486 674438 962488
rect 675183 962485 675249 962488
rect 41530 962190 41536 962254
rect 41600 962252 41606 962254
rect 41871 962252 41937 962255
rect 41600 962250 41937 962252
rect 41600 962194 41876 962250
rect 41932 962194 41937 962250
rect 41600 962192 41937 962194
rect 41600 962190 41606 962192
rect 41871 962189 41937 962192
rect 42351 962252 42417 962255
rect 42874 962252 42880 962254
rect 42351 962250 42880 962252
rect 42351 962194 42356 962250
rect 42412 962194 42880 962250
rect 42351 962192 42880 962194
rect 42351 962189 42417 962192
rect 42874 962190 42880 962192
rect 42944 962252 42950 962254
rect 61839 962252 61905 962255
rect 675375 962254 675441 962255
rect 675322 962252 675328 962254
rect 42944 962250 61905 962252
rect 42944 962194 61844 962250
rect 61900 962194 61905 962250
rect 42944 962192 61905 962194
rect 675284 962192 675328 962252
rect 675392 962250 675441 962254
rect 675436 962194 675441 962250
rect 42944 962190 42950 962192
rect 61839 962189 61905 962192
rect 675322 962190 675328 962192
rect 675392 962190 675441 962194
rect 675375 962189 675441 962190
rect 43066 962104 43072 962106
rect 42114 962044 43072 962104
rect 42114 961811 42174 962044
rect 43066 962042 43072 962044
rect 43136 962104 43142 962106
rect 62031 962104 62097 962107
rect 43136 962102 62097 962104
rect 43136 962046 62036 962102
rect 62092 962046 62097 962102
rect 43136 962044 62097 962046
rect 43136 962042 43142 962044
rect 62031 962041 62097 962044
rect 42063 961806 42174 961811
rect 42063 961750 42068 961806
rect 42124 961750 42174 961806
rect 42063 961748 42174 961750
rect 42063 961745 42129 961748
rect 675759 961512 675825 961515
rect 676666 961512 676672 961514
rect 675759 961510 676672 961512
rect 675759 961454 675764 961510
rect 675820 961454 676672 961510
rect 675759 961452 676672 961454
rect 675759 961449 675825 961452
rect 676666 961450 676672 961452
rect 676736 961450 676742 961514
rect 675471 961070 675537 961071
rect 675471 961068 675520 961070
rect 675428 961066 675520 961068
rect 675428 961010 675476 961066
rect 675428 961008 675520 961010
rect 675471 961006 675520 961008
rect 675584 961006 675590 961070
rect 675471 961005 675537 961006
rect 675663 960182 675729 960183
rect 675663 960180 675712 960182
rect 675620 960178 675712 960180
rect 675620 960122 675668 960178
rect 675620 960120 675712 960122
rect 675663 960118 675712 960120
rect 675776 960118 675782 960182
rect 675663 960117 675729 960118
rect 41338 959674 41344 959738
rect 41408 959736 41414 959738
rect 41775 959736 41841 959739
rect 41408 959734 41841 959736
rect 41408 959678 41780 959734
rect 41836 959678 41841 959734
rect 41408 959676 41841 959678
rect 41408 959674 41414 959676
rect 41775 959673 41841 959676
rect 41871 959146 41937 959147
rect 41871 959142 41920 959146
rect 41984 959144 41990 959146
rect 41871 959086 41876 959142
rect 41871 959082 41920 959086
rect 41984 959084 42028 959144
rect 41984 959082 41990 959084
rect 41871 959081 41937 959082
rect 59343 958700 59409 958703
rect 59343 958698 64416 958700
rect 59343 958642 59348 958698
rect 59404 958642 64416 958698
rect 59343 958640 64416 958642
rect 59343 958637 59409 958640
rect 42063 958406 42129 958407
rect 42063 958402 42112 958406
rect 42176 958404 42182 958406
rect 42063 958346 42068 958402
rect 42063 958342 42112 958346
rect 42176 958344 42220 958404
rect 42176 958342 42182 958344
rect 42063 958341 42129 958342
rect 42159 957812 42225 957815
rect 42298 957812 42304 957814
rect 42159 957810 42304 957812
rect 42159 957754 42164 957810
rect 42220 957754 42304 957810
rect 42159 957752 42304 957754
rect 42159 957749 42225 957752
rect 42298 957750 42304 957752
rect 42368 957750 42374 957814
rect 675759 957664 675825 957667
rect 676474 957664 676480 957666
rect 675759 957662 676480 957664
rect 675759 957606 675764 957662
rect 675820 957606 676480 957662
rect 675759 957604 676480 957606
rect 675759 957601 675825 957604
rect 676474 957602 676480 957604
rect 676544 957602 676550 957666
rect 42159 956184 42225 956187
rect 42490 956184 42496 956186
rect 42159 956182 42496 956184
rect 42159 956126 42164 956182
rect 42220 956126 42496 956182
rect 42159 956124 42496 956126
rect 42159 956121 42225 956124
rect 42490 956122 42496 956124
rect 42560 956122 42566 956186
rect 675130 955974 675136 956038
rect 675200 956036 675206 956038
rect 675471 956036 675537 956039
rect 675200 956034 675537 956036
rect 675200 955978 675476 956034
rect 675532 955978 675537 956034
rect 675200 955976 675537 955978
rect 675200 955974 675206 955976
rect 675471 955973 675537 955976
rect 675087 953520 675153 953523
rect 677050 953520 677056 953522
rect 675087 953518 677056 953520
rect 675087 953462 675092 953518
rect 675148 953462 677056 953518
rect 675087 953460 677056 953462
rect 675087 953457 675153 953460
rect 677050 953458 677056 953460
rect 677120 953458 677126 953522
rect 675183 953372 675249 953375
rect 676858 953372 676864 953374
rect 675183 953370 676864 953372
rect 675183 953314 675188 953370
rect 675244 953314 676864 953370
rect 675183 953312 676864 953314
rect 675183 953309 675249 953312
rect 676858 953310 676864 953312
rect 676928 953310 676934 953374
rect 654351 951004 654417 951007
rect 650208 951002 654417 951004
rect 650208 950946 654356 951002
rect 654412 950946 654417 951002
rect 650208 950944 654417 950946
rect 654351 950941 654417 950944
rect 674754 945383 674814 945942
rect 674703 945378 674814 945383
rect 674703 945322 674708 945378
rect 674764 945322 674814 945378
rect 674703 945320 674814 945322
rect 674703 945317 674769 945320
rect 674754 944791 674814 945054
rect 674703 944786 674814 944791
rect 674703 944730 674708 944786
rect 674764 944730 674814 944786
rect 674703 944728 674814 944730
rect 674703 944725 674769 944728
rect 59535 944344 59601 944347
rect 59535 944342 64416 944344
rect 59535 944286 59540 944342
rect 59596 944286 64416 944342
rect 59535 944284 64416 944286
rect 59535 944281 59601 944284
rect 674754 943755 674814 944240
rect 674703 943750 674814 943755
rect 674703 943694 674708 943750
rect 674764 943694 674814 943750
rect 674703 943692 674814 943694
rect 674703 943689 674769 943692
rect 674607 943160 674673 943163
rect 674754 943160 674814 943426
rect 674607 943158 674814 943160
rect 674607 943102 674612 943158
rect 674668 943102 674814 943158
rect 674607 943100 674814 943102
rect 674607 943097 674673 943100
rect 674415 942642 674481 942645
rect 674415 942640 674784 942642
rect 674415 942584 674420 942640
rect 674476 942584 674784 942640
rect 674415 942582 674784 942584
rect 674415 942579 674481 942582
rect 673839 941976 673905 941979
rect 673839 941974 674784 941976
rect 673839 941918 673844 941974
rect 673900 941918 674784 941974
rect 673839 941916 674784 941918
rect 673839 941913 673905 941916
rect 674746 940878 674752 940942
rect 674816 940878 674822 940942
rect 674754 940318 674814 940878
rect 674946 940647 675006 941132
rect 674895 940642 675006 940647
rect 674895 940586 674900 940642
rect 674956 940586 675006 940642
rect 674895 940584 675006 940586
rect 674895 940581 674961 940584
rect 674031 939608 674097 939611
rect 674031 939606 674814 939608
rect 674031 939550 674036 939606
rect 674092 939550 674814 939606
rect 674031 939548 674814 939550
rect 674031 939545 674097 939548
rect 674754 939504 674814 939548
rect 653775 939312 653841 939315
rect 650208 939310 653841 939312
rect 650208 939254 653780 939310
rect 653836 939254 653841 939310
rect 650208 939252 653841 939254
rect 653775 939249 653841 939252
rect 674554 938806 674560 938870
rect 674624 938868 674630 938870
rect 674624 938808 674814 938868
rect 674624 938806 674630 938808
rect 674754 938690 674814 938808
rect 674938 938362 674944 938426
rect 675008 938362 675014 938426
rect 674946 937802 675006 938362
rect 673935 937240 674001 937243
rect 673935 937238 674784 937240
rect 673935 937182 673940 937238
rect 673996 937182 674784 937238
rect 673935 937180 674784 937182
rect 673935 937177 674001 937180
rect 674127 936352 674193 936355
rect 674127 936350 674784 936352
rect 674127 936294 674132 936350
rect 674188 936294 674784 936350
rect 674127 936292 674784 936294
rect 674127 936289 674193 936292
rect 675898 935846 675904 935910
rect 675968 935846 675974 935910
rect 675906 935582 675966 935846
rect 674362 934662 674368 934726
rect 674432 934724 674438 934726
rect 674432 934664 674784 934724
rect 674432 934662 674438 934664
rect 675322 934514 675328 934578
rect 675392 934514 675398 934578
rect 675330 933954 675390 934514
rect 675130 933626 675136 933690
rect 675200 933626 675206 933690
rect 675138 933066 675198 933626
rect 676474 932590 676480 932654
rect 676544 932590 676550 932654
rect 676482 932474 676542 932590
rect 676666 931850 676672 931914
rect 676736 931850 676742 931914
rect 676674 931586 676734 931850
rect 677050 931406 677056 931470
rect 677120 931406 677126 931470
rect 677058 930846 677118 931406
rect 676858 930222 676864 930286
rect 676928 930222 676934 930286
rect 59535 929988 59601 929991
rect 59535 929986 64416 929988
rect 59535 929930 59540 929986
rect 59596 929930 64416 929986
rect 676866 929958 676926 930222
rect 59535 929928 64416 929930
rect 59535 929925 59601 929928
rect 679746 928659 679806 929144
rect 679746 928654 679857 928659
rect 679746 928598 679796 928654
rect 679852 928598 679857 928654
rect 679746 928596 679857 928598
rect 679791 928593 679857 928596
rect 679791 928064 679857 928067
rect 679746 928062 679857 928064
rect 679746 928006 679796 928062
rect 679852 928006 679857 928062
rect 679746 928001 679857 928006
rect 679746 927664 679806 928001
rect 654447 927472 654513 927475
rect 650208 927470 654513 927472
rect 650208 927414 654452 927470
rect 654508 927414 654513 927470
rect 650208 927412 654513 927414
rect 654447 927409 654513 927412
rect 654447 915780 654513 915783
rect 650208 915778 654513 915780
rect 650208 915722 654452 915778
rect 654508 915722 654513 915778
rect 650208 915720 654513 915722
rect 654447 915717 654513 915720
rect 59535 915484 59601 915487
rect 59535 915482 64416 915484
rect 59535 915426 59540 915482
rect 59596 915426 64416 915482
rect 59535 915424 64416 915426
rect 59535 915421 59601 915424
rect 42639 908084 42705 908087
rect 42336 908082 42705 908084
rect 42336 908026 42644 908082
rect 42700 908026 42705 908082
rect 42336 908024 42705 908026
rect 42639 908021 42705 908024
rect 42255 907492 42321 907495
rect 42255 907490 42366 907492
rect 42255 907434 42260 907490
rect 42316 907434 42366 907490
rect 42255 907429 42366 907434
rect 42306 907314 42366 907429
rect 42874 907134 42880 907198
rect 42944 907196 42950 907198
rect 43119 907196 43185 907199
rect 42944 907194 43185 907196
rect 42944 907138 43124 907194
rect 43180 907138 43185 907194
rect 42944 907136 43185 907138
rect 42944 907134 42950 907136
rect 43119 907133 43185 907136
rect 42351 906752 42417 906755
rect 42306 906750 42417 906752
rect 42306 906694 42356 906750
rect 42412 906694 42417 906750
rect 42306 906689 42417 906694
rect 42306 906426 42366 906689
rect 40386 905423 40446 905686
rect 40335 905418 40446 905423
rect 40335 905362 40340 905418
rect 40396 905362 40446 905418
rect 40335 905360 40446 905362
rect 40335 905357 40401 905360
rect 42639 904828 42705 904831
rect 42336 904826 42705 904828
rect 42336 904770 42644 904826
rect 42700 904770 42705 904826
rect 42336 904768 42705 904770
rect 42639 904765 42705 904768
rect 43215 904236 43281 904239
rect 44751 904236 44817 904239
rect 42306 904234 44817 904236
rect 42306 904178 43220 904234
rect 43276 904178 44756 904234
rect 44812 904178 44817 904234
rect 42306 904176 44817 904178
rect 42306 904132 42366 904176
rect 43215 904173 43281 904176
rect 44751 904173 44817 904176
rect 654447 904088 654513 904091
rect 650208 904086 654513 904088
rect 650208 904030 654452 904086
rect 654508 904030 654513 904086
rect 650208 904028 654513 904030
rect 654447 904025 654513 904028
rect 42682 903348 42688 903350
rect 42336 903288 42688 903348
rect 42682 903286 42688 903288
rect 42752 903348 42758 903350
rect 44559 903348 44625 903351
rect 42752 903346 44625 903348
rect 42752 903290 44564 903346
rect 44620 903290 44625 903346
rect 42752 903288 44625 903290
rect 42752 903286 42758 903288
rect 44559 903285 44625 903288
rect 42490 903052 42496 903054
rect 42306 902992 42496 903052
rect 42306 902504 42366 902992
rect 42490 902990 42496 902992
rect 42560 902990 42566 903054
rect 41722 902250 41728 902314
rect 41792 902250 41798 902314
rect 41730 901690 41790 902250
rect 43215 901572 43281 901575
rect 40002 901570 43281 901572
rect 40002 901514 43220 901570
rect 43276 901514 43281 901570
rect 40002 901512 43281 901514
rect 40002 901427 40062 901512
rect 43215 901509 43281 901512
rect 40002 901422 40113 901427
rect 40002 901366 40052 901422
rect 40108 901366 40113 901422
rect 40002 901364 40113 901366
rect 40047 901361 40113 901364
rect 59535 901276 59601 901279
rect 59535 901274 64416 901276
rect 59535 901218 59540 901274
rect 59596 901218 64416 901274
rect 59535 901216 64416 901218
rect 59535 901213 59601 901216
rect 43023 901128 43089 901131
rect 42306 901126 43089 901128
rect 42306 901070 43028 901126
rect 43084 901070 43089 901126
rect 42306 901068 43089 901070
rect 42306 900876 42366 901068
rect 43023 901065 43089 901068
rect 42298 900622 42304 900686
rect 42368 900622 42374 900686
rect 42306 900062 42366 900622
rect 41530 899734 41536 899798
rect 41600 899734 41606 899798
rect 41538 899322 41598 899734
rect 40570 899142 40576 899206
rect 40640 899142 40646 899206
rect 40578 898582 40638 899142
rect 42927 897724 42993 897727
rect 42336 897722 42993 897724
rect 42336 897666 42932 897722
rect 42988 897666 42993 897722
rect 42336 897664 42993 897666
rect 42927 897661 42993 897664
rect 42106 897514 42112 897578
rect 42176 897514 42182 897578
rect 42114 896954 42174 897514
rect 41914 896626 41920 896690
rect 41984 896626 41990 896690
rect 41922 896066 41982 896626
rect 40378 895590 40384 895654
rect 40448 895590 40454 895654
rect 40386 895326 40446 895590
rect 40954 894998 40960 895062
rect 41024 894998 41030 895062
rect 40962 894586 41022 894998
rect 41338 894406 41344 894470
rect 41408 894406 41414 894470
rect 41346 893846 41406 894406
rect 41146 893518 41152 893582
rect 41216 893518 41222 893582
rect 41154 892958 41214 893518
rect 650031 892840 650097 892843
rect 649986 892838 650097 892840
rect 649986 892782 650036 892838
rect 650092 892782 650097 892838
rect 649986 892777 650097 892782
rect 40762 892482 40768 892546
rect 40832 892544 40838 892546
rect 40832 892484 41022 892544
rect 40832 892482 40838 892484
rect 40962 892218 41022 892484
rect 649986 892366 650046 892777
rect 42306 891215 42366 891330
rect 42306 891210 42417 891215
rect 42306 891154 42356 891210
rect 42412 891154 42417 891210
rect 42306 891152 42417 891154
rect 42351 891149 42417 891152
rect 42306 889735 42366 889850
rect 42306 889730 42417 889735
rect 42306 889674 42356 889730
rect 42412 889674 42417 889730
rect 42306 889672 42417 889674
rect 42351 889669 42417 889672
rect 43119 887364 43185 887367
rect 42882 887362 43185 887364
rect 42882 887306 43124 887362
rect 43180 887306 43185 887362
rect 42882 887304 43185 887306
rect 42882 887218 42942 887304
rect 43119 887301 43185 887304
rect 42874 887154 42880 887218
rect 42944 887154 42950 887218
rect 59535 886772 59601 886775
rect 59535 886770 64416 886772
rect 59535 886714 59540 886770
rect 59596 886714 64416 886770
rect 59535 886712 64416 886714
rect 59535 886709 59601 886712
rect 654447 880556 654513 880559
rect 650208 880554 654513 880556
rect 650208 880498 654452 880554
rect 654508 880498 654513 880554
rect 650208 880496 654513 880498
rect 654447 880493 654513 880496
rect 674362 876350 674368 876414
rect 674432 876412 674438 876414
rect 675087 876412 675153 876415
rect 674432 876410 675153 876412
rect 674432 876354 675092 876410
rect 675148 876354 675153 876410
rect 674432 876352 675153 876354
rect 674432 876350 674438 876352
rect 675087 876349 675153 876352
rect 675759 876412 675825 876415
rect 676666 876412 676672 876414
rect 675759 876410 676672 876412
rect 675759 876354 675764 876410
rect 675820 876354 676672 876410
rect 675759 876352 676672 876354
rect 675759 876349 675825 876352
rect 676666 876350 676672 876352
rect 676736 876350 676742 876414
rect 674746 876202 674752 876266
rect 674816 876264 674822 876266
rect 675087 876264 675153 876267
rect 674816 876262 675153 876264
rect 674816 876206 675092 876262
rect 675148 876206 675153 876262
rect 674816 876204 675153 876206
rect 674816 876202 674822 876204
rect 675087 876201 675153 876204
rect 675279 875820 675345 875823
rect 675706 875820 675712 875822
rect 675279 875818 675712 875820
rect 675279 875762 675284 875818
rect 675340 875762 675712 875818
rect 675279 875760 675712 875762
rect 675279 875757 675345 875760
rect 675706 875758 675712 875760
rect 675776 875758 675782 875822
rect 674938 873982 674944 874046
rect 675008 874044 675014 874046
rect 675471 874044 675537 874047
rect 675008 874042 675537 874044
rect 675008 873986 675476 874042
rect 675532 873986 675537 874042
rect 675008 873984 675537 873986
rect 675008 873982 675014 873984
rect 675471 873981 675537 873984
rect 674554 873390 674560 873454
rect 674624 873452 674630 873454
rect 675375 873452 675441 873455
rect 674624 873450 675441 873452
rect 674624 873394 675380 873450
rect 675436 873394 675441 873450
rect 674624 873392 675441 873394
rect 674624 873390 674630 873392
rect 675375 873389 675441 873392
rect 674170 872798 674176 872862
rect 674240 872860 674246 872862
rect 675375 872860 675441 872863
rect 674240 872858 675441 872860
rect 674240 872802 675380 872858
rect 675436 872802 675441 872858
rect 674240 872800 675441 872802
rect 674240 872798 674246 872800
rect 675375 872797 675441 872800
rect 58959 872416 59025 872419
rect 675567 872418 675633 872419
rect 58959 872414 64416 872416
rect 58959 872358 58964 872414
rect 59020 872358 64416 872414
rect 58959 872356 64416 872358
rect 58959 872353 59025 872356
rect 675514 872354 675520 872418
rect 675584 872416 675633 872418
rect 675584 872414 675676 872416
rect 675628 872358 675676 872414
rect 675584 872356 675676 872358
rect 675584 872354 675633 872356
rect 675567 872353 675633 872354
rect 675375 869902 675441 869903
rect 675322 869900 675328 869902
rect 675284 869840 675328 869900
rect 675392 869898 675441 869902
rect 675436 869842 675441 869898
rect 675322 869838 675328 869840
rect 675392 869838 675441 869842
rect 675375 869837 675441 869838
rect 654447 868864 654513 868867
rect 650208 868862 654513 868864
rect 650208 868806 654452 868862
rect 654508 868806 654513 868862
rect 650208 868804 654513 868806
rect 654447 868801 654513 868804
rect 675130 866878 675136 866942
rect 675200 866940 675206 866942
rect 675375 866940 675441 866943
rect 675200 866938 675441 866940
rect 675200 866882 675380 866938
rect 675436 866882 675441 866938
rect 675200 866880 675441 866882
rect 675200 866878 675206 866880
rect 675375 866877 675441 866880
rect 42298 866434 42304 866498
rect 42368 866496 42374 866498
rect 42874 866496 42880 866498
rect 42368 866436 42880 866496
rect 42368 866434 42374 866436
rect 42874 866434 42880 866436
rect 42944 866434 42950 866498
rect 675471 864722 675537 864723
rect 675471 864718 675520 864722
rect 675584 864720 675590 864722
rect 675471 864662 675476 864718
rect 675471 864658 675520 864662
rect 675584 864660 675628 864720
rect 675584 864658 675590 864660
rect 675471 864657 675537 864658
rect 42682 864214 42688 864278
rect 42752 864214 42758 864278
rect 42690 864130 42750 864214
rect 42682 864066 42688 864130
rect 42752 864066 42758 864130
rect 675663 862946 675729 862947
rect 675663 862942 675712 862946
rect 675776 862944 675782 862946
rect 675663 862886 675668 862942
rect 675663 862882 675712 862886
rect 675776 862884 675820 862944
rect 675776 862882 675782 862884
rect 675663 862881 675729 862882
rect 42490 858146 42496 858210
rect 42560 858146 42566 858210
rect 42498 858060 42558 858146
rect 43258 858060 43264 858062
rect 42498 858000 43264 858060
rect 43258 857998 43264 858000
rect 43328 857998 43334 858062
rect 59535 858060 59601 858063
rect 59535 858058 64416 858060
rect 59535 858002 59540 858058
rect 59596 858002 64416 858058
rect 59535 858000 64416 858002
rect 59535 857997 59601 858000
rect 654447 857172 654513 857175
rect 650208 857170 654513 857172
rect 650208 857114 654452 857170
rect 654508 857114 654513 857170
rect 650208 857112 654513 857114
rect 654447 857109 654513 857112
rect 40815 852732 40881 852735
rect 42682 852732 42688 852734
rect 40815 852730 42688 852732
rect 40815 852674 40820 852730
rect 40876 852674 42688 852730
rect 40815 852672 42688 852674
rect 40815 852669 40881 852672
rect 42682 852670 42688 852672
rect 42752 852670 42758 852734
rect 649551 846072 649617 846075
rect 649551 846070 649662 846072
rect 649551 846014 649556 846070
rect 649612 846014 649662 846070
rect 649551 846009 649662 846014
rect 649602 845450 649662 846009
rect 59535 843704 59601 843707
rect 59535 843702 64416 843704
rect 59535 843646 59540 843702
rect 59596 843646 64416 843702
rect 59535 843644 64416 843646
rect 59535 843641 59601 843644
rect 39994 842606 40000 842670
rect 40064 842668 40070 842670
rect 40143 842668 40209 842671
rect 40064 842666 40209 842668
rect 40064 842610 40148 842666
rect 40204 842610 40209 842666
rect 40064 842608 40209 842610
rect 40064 842606 40070 842608
rect 40143 842605 40209 842608
rect 43066 840978 43072 841042
rect 43136 840978 43142 841042
rect 43074 840746 43134 840978
rect 43066 840682 43072 840746
rect 43136 840682 43142 840746
rect 654447 833640 654513 833643
rect 650208 833638 654513 833640
rect 650208 833582 654452 833638
rect 654508 833582 654513 833638
rect 650208 833580 654513 833582
rect 654447 833577 654513 833580
rect 42874 830914 42880 830978
rect 42944 830976 42950 830978
rect 43258 830976 43264 830978
rect 42944 830916 43264 830976
rect 42944 830914 42950 830916
rect 43258 830914 43264 830916
rect 43328 830914 43334 830978
rect 58191 829496 58257 829499
rect 58191 829494 64416 829496
rect 58191 829438 58196 829494
rect 58252 829438 64416 829494
rect 58191 829436 64416 829438
rect 58191 829433 58257 829436
rect 39951 827574 40017 827575
rect 39951 827570 40000 827574
rect 40064 827572 40070 827574
rect 39951 827514 39956 827570
rect 39951 827510 40000 827514
rect 40064 827512 40108 827572
rect 40064 827510 40070 827512
rect 39951 827509 40017 827510
rect 42351 823872 42417 823875
rect 42306 823870 42417 823872
rect 42306 823814 42356 823870
rect 42412 823814 42417 823870
rect 42306 823809 42417 823814
rect 42306 823694 42366 823809
rect 42306 822688 42366 822880
rect 42447 822688 42513 822691
rect 42306 822686 42513 822688
rect 42306 822630 42452 822686
rect 42508 822630 42513 822686
rect 42306 822628 42513 822630
rect 42447 822625 42513 822628
rect 42351 822244 42417 822247
rect 42306 822242 42417 822244
rect 42306 822186 42356 822242
rect 42412 822186 42417 822242
rect 42306 822181 42417 822186
rect 42306 822066 42366 822181
rect 654447 821948 654513 821951
rect 650208 821946 654513 821948
rect 650208 821890 654452 821946
rect 654508 821890 654513 821946
rect 650208 821888 654513 821890
rect 654447 821885 654513 821888
rect 43215 821208 43281 821211
rect 42336 821206 43281 821208
rect 42336 821150 43220 821206
rect 43276 821150 43281 821206
rect 42336 821148 43281 821150
rect 43215 821145 43281 821148
rect 40335 820764 40401 820767
rect 40335 820762 40446 820764
rect 40335 820706 40340 820762
rect 40396 820706 40446 820762
rect 40335 820701 40446 820706
rect 40386 820438 40446 820701
rect 40194 819435 40254 819698
rect 40815 819580 40881 819583
rect 40143 819430 40254 819435
rect 40143 819374 40148 819430
rect 40204 819374 40254 819430
rect 40143 819372 40254 819374
rect 40770 819578 40881 819580
rect 40770 819522 40820 819578
rect 40876 819522 40881 819578
rect 40770 819517 40881 819522
rect 40143 819369 40209 819372
rect 40770 818398 40830 819517
rect 40762 818334 40768 818398
rect 40832 818334 40838 818398
rect 42306 817955 42366 818070
rect 42306 817950 42417 817955
rect 42306 817894 42356 817950
rect 42412 817894 42417 817950
rect 42306 817892 42417 817894
rect 42351 817889 42417 817892
rect 40194 816771 40254 817330
rect 40194 816766 40305 816771
rect 40194 816710 40244 816766
rect 40300 816710 40305 816766
rect 40194 816708 40305 816710
rect 40239 816705 40305 816708
rect 37314 815883 37374 816442
rect 37263 815878 37374 815883
rect 37263 815822 37268 815878
rect 37324 815822 37374 815878
rect 37263 815820 37374 815822
rect 37263 815817 37329 815820
rect 42306 815288 42366 815702
rect 42447 815288 42513 815291
rect 42306 815286 42513 815288
rect 42306 815230 42452 815286
rect 42508 815230 42513 815286
rect 42306 815228 42513 815230
rect 42447 815225 42513 815228
rect 59535 814992 59601 814995
rect 59535 814990 64416 814992
rect 41922 814403 41982 814962
rect 59535 814934 59540 814990
rect 59596 814934 64416 814990
rect 59535 814932 64416 814934
rect 59535 814929 59601 814932
rect 41922 814398 42033 814403
rect 41922 814342 41972 814398
rect 42028 814342 42033 814398
rect 41922 814340 42033 814342
rect 41967 814337 42033 814340
rect 41922 813663 41982 814222
rect 41871 813658 41982 813663
rect 41871 813602 41876 813658
rect 41932 813602 41982 813658
rect 41871 813600 41982 813602
rect 41871 813597 41937 813600
rect 37314 812775 37374 813334
rect 37314 812770 37425 812775
rect 37314 812714 37364 812770
rect 37420 812714 37425 812770
rect 37314 812712 37425 812714
rect 37359 812709 37425 812712
rect 42306 812328 42366 812520
rect 43119 812328 43185 812331
rect 42306 812326 43185 812328
rect 42306 812270 43124 812326
rect 43180 812270 43185 812326
rect 42306 812268 43185 812270
rect 43119 812265 43185 812268
rect 41730 811147 41790 811706
rect 41679 811142 41790 811147
rect 41679 811086 41684 811142
rect 41740 811086 41790 811142
rect 41679 811084 41790 811086
rect 41679 811081 41745 811084
rect 42306 810404 42366 810892
rect 43119 810404 43185 810407
rect 42306 810402 43185 810404
rect 42306 810346 43124 810402
rect 43180 810346 43185 810402
rect 42306 810344 43185 810346
rect 43119 810341 43185 810344
rect 654447 810256 654513 810259
rect 650208 810254 654513 810256
rect 41730 809667 41790 810226
rect 650208 810198 654452 810254
rect 654508 810198 654513 810254
rect 650208 810196 654513 810198
rect 654447 810193 654513 810196
rect 41730 809662 41841 809667
rect 41730 809606 41780 809662
rect 41836 809606 41841 809662
rect 41730 809604 41841 809606
rect 41775 809601 41841 809604
rect 42114 809223 42174 809412
rect 42063 809218 42174 809223
rect 42063 809162 42068 809218
rect 42124 809162 42174 809218
rect 42063 809160 42174 809162
rect 42063 809157 42129 809160
rect 42114 808335 42174 808598
rect 42114 808330 42225 808335
rect 42114 808274 42164 808330
rect 42220 808274 42225 808330
rect 42114 808272 42225 808274
rect 42159 808269 42225 808272
rect 42306 807296 42366 807784
rect 42927 807296 42993 807299
rect 42306 807294 42993 807296
rect 42306 807238 42932 807294
rect 42988 807238 42993 807294
rect 42306 807236 42993 807238
rect 42927 807233 42993 807236
rect 42306 806408 42366 806970
rect 42306 806348 42750 806408
rect 42690 805964 42750 806348
rect 42306 805904 42750 805964
rect 42306 805227 42366 805904
rect 42255 805222 42366 805227
rect 42255 805166 42260 805222
rect 42316 805166 42366 805222
rect 42255 805164 42366 805166
rect 42255 805161 42321 805164
rect 37263 802116 37329 802119
rect 41338 802116 41344 802118
rect 37263 802114 41344 802116
rect 37263 802058 37268 802114
rect 37324 802058 41344 802114
rect 37263 802056 41344 802058
rect 37263 802053 37329 802056
rect 41338 802054 41344 802056
rect 41408 802054 41414 802118
rect 37359 801968 37425 801971
rect 41530 801968 41536 801970
rect 37359 801966 41536 801968
rect 37359 801910 37364 801966
rect 37420 801910 41536 801966
rect 37359 801908 41536 801910
rect 37359 801905 37425 801908
rect 41530 801906 41536 801908
rect 41600 801906 41606 801970
rect 59535 800636 59601 800639
rect 59535 800634 64416 800636
rect 59535 800578 59540 800634
rect 59596 800578 64416 800634
rect 59535 800576 64416 800578
rect 59535 800573 59601 800576
rect 41679 800488 41745 800491
rect 42682 800488 42688 800490
rect 41679 800486 42688 800488
rect 41679 800430 41684 800486
rect 41740 800430 42688 800486
rect 41679 800428 42688 800430
rect 41679 800425 41745 800428
rect 42682 800426 42688 800428
rect 42752 800426 42758 800490
rect 41775 800342 41841 800343
rect 41722 800340 41728 800342
rect 41684 800280 41728 800340
rect 41792 800338 41841 800342
rect 41836 800282 41841 800338
rect 41722 800278 41728 800280
rect 41792 800278 41841 800282
rect 41775 800277 41841 800278
rect 42063 800342 42129 800343
rect 42063 800338 42112 800342
rect 42176 800340 42182 800342
rect 42063 800282 42068 800338
rect 42063 800278 42112 800282
rect 42176 800280 42220 800340
rect 42176 800278 42182 800280
rect 42063 800277 42129 800278
rect 42255 800046 42321 800047
rect 42255 800042 42304 800046
rect 42368 800044 42374 800046
rect 42255 799986 42260 800042
rect 42255 799982 42304 799986
rect 42368 799984 42412 800044
rect 42368 799982 42374 799984
rect 42255 799981 42321 799982
rect 649935 799156 650001 799159
rect 649935 799154 650046 799156
rect 649935 799098 649940 799154
rect 649996 799098 650046 799154
rect 649935 799093 650046 799098
rect 649986 798534 650046 799093
rect 42298 797910 42304 797974
rect 42368 797972 42374 797974
rect 42447 797972 42513 797975
rect 42368 797970 42513 797972
rect 42368 797914 42452 797970
rect 42508 797914 42513 797970
rect 42368 797912 42513 797914
rect 42368 797910 42374 797912
rect 42447 797909 42513 797912
rect 42735 794866 42801 794867
rect 42682 794802 42688 794866
rect 42752 794864 42801 794866
rect 42752 794862 42844 794864
rect 42796 794806 42844 794862
rect 42752 794804 42844 794806
rect 42752 794802 42801 794804
rect 42735 794801 42801 794802
rect 41775 794274 41841 794275
rect 41722 794210 41728 794274
rect 41792 794272 41841 794274
rect 41792 794270 41884 794272
rect 41836 794214 41884 794270
rect 41792 794212 41884 794214
rect 41792 794210 41841 794212
rect 41775 794209 41841 794210
rect 41722 794062 41728 794126
rect 41792 794124 41798 794126
rect 43066 794124 43072 794126
rect 41792 794064 43072 794124
rect 41792 794062 41798 794064
rect 43066 794062 43072 794064
rect 43136 794062 43142 794126
rect 42106 792138 42112 792202
rect 42176 792200 42182 792202
rect 42255 792200 42321 792203
rect 42176 792198 42321 792200
rect 42176 792142 42260 792198
rect 42316 792142 42321 792198
rect 42176 792140 42321 792142
rect 42176 792138 42182 792140
rect 42255 792137 42321 792140
rect 42735 792052 42801 792055
rect 43119 792052 43185 792055
rect 42735 792050 43185 792052
rect 42735 791994 42740 792050
rect 42796 791994 43124 792050
rect 43180 791994 43185 792050
rect 42735 791992 43185 791994
rect 42735 791989 42801 791992
rect 43119 791989 43185 791992
rect 41530 791842 41536 791906
rect 41600 791904 41606 791906
rect 42447 791904 42513 791907
rect 41600 791902 42513 791904
rect 41600 791846 42452 791902
rect 42508 791846 42513 791902
rect 41600 791844 42513 791846
rect 41600 791842 41606 791844
rect 42447 791841 42513 791844
rect 41338 791694 41344 791758
rect 41408 791756 41414 791758
rect 42735 791756 42801 791759
rect 41408 791754 42801 791756
rect 41408 791698 42740 791754
rect 42796 791698 42801 791754
rect 41408 791696 42801 791698
rect 41408 791694 41414 791696
rect 42735 791693 42801 791696
rect 41775 791166 41841 791167
rect 41722 791102 41728 791166
rect 41792 791164 41841 791166
rect 41792 791162 41884 791164
rect 41836 791106 41884 791162
rect 41792 791104 41884 791106
rect 41792 791102 41841 791104
rect 41775 791101 41841 791102
rect 41914 790954 41920 791018
rect 41984 791016 41990 791018
rect 42159 791016 42225 791019
rect 42490 791016 42496 791018
rect 41984 791014 42496 791016
rect 41984 790958 42164 791014
rect 42220 790958 42496 791014
rect 41984 790956 42496 790958
rect 41984 790954 41990 790956
rect 42159 790953 42225 790956
rect 42490 790954 42496 790956
rect 42560 790954 42566 791018
rect 675759 787908 675825 787911
rect 676282 787908 676288 787910
rect 675759 787906 676288 787908
rect 675759 787850 675764 787906
rect 675820 787850 676288 787906
rect 675759 787848 676288 787850
rect 675759 787845 675825 787848
rect 676282 787846 676288 787848
rect 676352 787846 676358 787910
rect 673978 787402 673984 787466
rect 674048 787464 674054 787466
rect 675471 787464 675537 787467
rect 674048 787462 675537 787464
rect 674048 787406 675476 787462
rect 675532 787406 675537 787462
rect 674048 787404 675537 787406
rect 674048 787402 674054 787404
rect 675471 787401 675537 787404
rect 654447 786724 654513 786727
rect 650208 786722 654513 786724
rect 650208 786666 654452 786722
rect 654508 786666 654513 786722
rect 650208 786664 654513 786666
rect 654447 786661 654513 786664
rect 675759 786724 675825 786727
rect 675898 786724 675904 786726
rect 675759 786722 675904 786724
rect 675759 786666 675764 786722
rect 675820 786666 675904 786722
rect 675759 786664 675904 786666
rect 675759 786661 675825 786664
rect 675898 786662 675904 786664
rect 675968 786662 675974 786726
rect 58959 786280 59025 786283
rect 58959 786278 64416 786280
rect 58959 786222 58964 786278
rect 59020 786222 64416 786278
rect 58959 786220 64416 786222
rect 58959 786217 59025 786220
rect 675759 784208 675825 784211
rect 676090 784208 676096 784210
rect 675759 784206 676096 784208
rect 675759 784150 675764 784206
rect 675820 784150 676096 784206
rect 675759 784148 676096 784150
rect 675759 784145 675825 784148
rect 676090 784146 676096 784148
rect 676160 784146 676166 784210
rect 675759 781988 675825 781991
rect 676474 781988 676480 781990
rect 675759 781986 676480 781988
rect 675759 781930 675764 781986
rect 675820 781930 676480 781986
rect 675759 781928 676480 781930
rect 675759 781925 675825 781928
rect 676474 781926 676480 781928
rect 676544 781926 676550 781990
rect 42735 780508 42801 780511
rect 42336 780506 42801 780508
rect 42336 780450 42740 780506
rect 42796 780450 42801 780506
rect 42336 780448 42801 780450
rect 42735 780445 42801 780448
rect 674223 780508 674289 780511
rect 677050 780508 677056 780510
rect 674223 780506 677056 780508
rect 674223 780450 674228 780506
rect 674284 780450 677056 780506
rect 674223 780448 677056 780450
rect 674223 780445 674289 780448
rect 677050 780446 677056 780448
rect 677120 780446 677126 780510
rect 42447 779916 42513 779919
rect 42306 779914 42513 779916
rect 42306 779858 42452 779914
rect 42508 779858 42513 779914
rect 42306 779856 42513 779858
rect 42306 779664 42366 779856
rect 42447 779853 42513 779856
rect 42735 778880 42801 778883
rect 42336 778878 42801 778880
rect 42336 778822 42740 778878
rect 42796 778822 42801 778878
rect 42336 778820 42801 778822
rect 42735 778817 42801 778820
rect 42306 777992 42366 778036
rect 43407 777992 43473 777995
rect 42306 777990 43473 777992
rect 42306 777934 43412 777990
rect 43468 777934 43473 777990
rect 42306 777932 43473 777934
rect 43407 777929 43473 777932
rect 674991 777548 675057 777551
rect 677050 777548 677056 777550
rect 674991 777546 677056 777548
rect 674991 777490 674996 777546
rect 675052 777490 677056 777546
rect 674991 777488 677056 777490
rect 674991 777485 675057 777488
rect 677050 777486 677056 777488
rect 677120 777486 677126 777550
rect 674799 777400 674865 777403
rect 676858 777400 676864 777402
rect 674799 777398 676864 777400
rect 674799 777342 674804 777398
rect 674860 777342 676864 777398
rect 674799 777340 676864 777342
rect 674799 777337 674865 777340
rect 676858 777338 676864 777340
rect 676928 777338 676934 777402
rect 43215 777252 43281 777255
rect 42336 777250 43281 777252
rect 42336 777194 43220 777250
rect 43276 777194 43281 777250
rect 42336 777192 43281 777194
rect 43215 777189 43281 777192
rect 43215 776512 43281 776515
rect 42336 776510 43281 776512
rect 42336 776454 43220 776510
rect 43276 776454 43281 776510
rect 42336 776452 43281 776454
rect 43215 776449 43281 776452
rect 40770 775182 40830 775742
rect 40762 775118 40768 775182
rect 40832 775118 40838 775182
rect 654447 775032 654513 775035
rect 650208 775030 654513 775032
rect 650208 774974 654452 775030
rect 654508 774974 654513 775030
rect 650208 774972 654513 774974
rect 654447 774969 654513 774972
rect 42831 774884 42897 774887
rect 42336 774882 42897 774884
rect 42336 774826 42836 774882
rect 42892 774826 42897 774882
rect 42336 774824 42897 774826
rect 42831 774821 42897 774824
rect 38850 773555 38910 774114
rect 38799 773550 38910 773555
rect 38799 773494 38804 773550
rect 38860 773494 38910 773550
rect 38799 773492 38910 773494
rect 38799 773489 38865 773492
rect 35970 772667 36030 773226
rect 676858 773046 676864 773110
rect 676928 773108 676934 773110
rect 677818 773108 677824 773110
rect 676928 773048 677824 773108
rect 676928 773046 676934 773048
rect 677818 773046 677824 773048
rect 677888 773046 677894 773110
rect 676858 772898 676864 772962
rect 676928 772960 676934 772962
rect 677242 772960 677248 772962
rect 676928 772900 677248 772960
rect 676928 772898 676934 772900
rect 677242 772898 677248 772900
rect 677312 772898 677318 772962
rect 35919 772662 36030 772667
rect 35919 772606 35924 772662
rect 35980 772606 36030 772662
rect 35919 772604 36030 772606
rect 674319 772664 674385 772667
rect 677242 772664 677248 772666
rect 674319 772662 677248 772664
rect 674319 772606 674324 772662
rect 674380 772606 677248 772662
rect 674319 772604 677248 772606
rect 35919 772601 35985 772604
rect 674319 772601 674385 772604
rect 677242 772602 677248 772604
rect 677312 772602 677318 772666
rect 42927 772516 42993 772519
rect 42336 772514 42993 772516
rect 42336 772458 42932 772514
rect 42988 772458 42993 772514
rect 42336 772456 42993 772458
rect 42927 772453 42993 772456
rect 59535 771924 59601 771927
rect 59535 771922 64416 771924
rect 59535 771866 59540 771922
rect 59596 771866 64416 771922
rect 59535 771864 64416 771866
rect 59535 771861 59601 771864
rect 41922 771187 41982 771746
rect 41922 771182 42033 771187
rect 41922 771126 41972 771182
rect 42028 771126 42033 771182
rect 41922 771124 42033 771126
rect 41967 771121 42033 771124
rect 41730 770447 41790 771006
rect 41730 770442 41841 770447
rect 41730 770386 41780 770442
rect 41836 770386 41841 770442
rect 41730 770384 41841 770386
rect 41775 770381 41841 770384
rect 37314 769559 37374 770118
rect 37314 769554 37425 769559
rect 37314 769498 37364 769554
rect 37420 769498 37425 769554
rect 37314 769496 37425 769498
rect 37359 769493 37425 769496
rect 42306 769112 42366 769378
rect 42447 769112 42513 769115
rect 42306 769110 42513 769112
rect 42306 769054 42452 769110
rect 42508 769054 42513 769110
rect 42306 769052 42513 769054
rect 42447 769049 42513 769052
rect 41922 767931 41982 768490
rect 41871 767926 41982 767931
rect 41871 767870 41876 767926
rect 41932 767870 41982 767926
rect 41871 767868 41982 767870
rect 41871 767865 41937 767868
rect 43119 767780 43185 767783
rect 42336 767778 43185 767780
rect 42336 767722 43124 767778
rect 43180 767722 43185 767778
rect 42336 767720 43185 767722
rect 43119 767717 43185 767720
rect 674703 767780 674769 767783
rect 674703 767778 674814 767780
rect 674703 767722 674708 767778
rect 674764 767722 674814 767778
rect 674703 767717 674814 767722
rect 674754 767454 674814 767717
rect 42927 767040 42993 767043
rect 42336 767038 42993 767040
rect 42336 766982 42932 767038
rect 42988 766982 42993 767038
rect 42336 766980 42993 766982
rect 42927 766977 42993 766980
rect 674703 766892 674769 766895
rect 674703 766890 674814 766892
rect 674703 766834 674708 766890
rect 674764 766834 674814 766890
rect 674703 766829 674814 766834
rect 674754 766714 674814 766829
rect 42114 766007 42174 766196
rect 42114 766002 42225 766007
rect 42114 765946 42164 766002
rect 42220 765946 42225 766002
rect 42114 765944 42225 765946
rect 42159 765941 42225 765944
rect 674319 765856 674385 765859
rect 674319 765854 674784 765856
rect 674319 765798 674324 765854
rect 674380 765798 674784 765854
rect 674319 765796 674784 765798
rect 674319 765793 674385 765796
rect 42114 765267 42174 765382
rect 42063 765262 42174 765267
rect 42063 765206 42068 765262
rect 42124 765206 42174 765262
rect 42063 765204 42174 765206
rect 674703 765264 674769 765267
rect 674703 765262 674814 765264
rect 674703 765206 674708 765262
rect 674764 765206 674814 765262
rect 42063 765201 42129 765204
rect 674703 765201 674814 765206
rect 674754 765086 674814 765201
rect 42735 764598 42801 764601
rect 42336 764596 42801 764598
rect 42336 764540 42740 764596
rect 42796 764540 42801 764596
rect 42336 764538 42801 764540
rect 42735 764535 42801 764538
rect 674754 764083 674814 764198
rect 674703 764078 674814 764083
rect 674703 764022 674708 764078
rect 674764 764022 674814 764078
rect 674703 764020 674814 764022
rect 674703 764017 674769 764020
rect 42306 763194 42366 763754
rect 674754 763343 674814 763532
rect 654447 763340 654513 763343
rect 650208 763338 654513 763340
rect 650208 763282 654452 763338
rect 654508 763282 654513 763338
rect 650208 763280 654513 763282
rect 654447 763277 654513 763280
rect 674703 763338 674814 763343
rect 674703 763282 674708 763338
rect 674764 763282 674814 763338
rect 674703 763280 674814 763282
rect 674703 763277 674769 763280
rect 42298 763130 42304 763194
rect 42368 763130 42374 763194
rect 42298 762686 42304 762750
rect 42368 762686 42374 762750
rect 42306 762304 42366 762686
rect 674754 762603 674814 762718
rect 674703 762598 674814 762603
rect 674703 762542 674708 762598
rect 674764 762542 674814 762598
rect 674703 762540 674814 762542
rect 674703 762537 674769 762540
rect 674746 762390 674752 762454
rect 674816 762390 674822 762454
rect 44847 762304 44913 762307
rect 42306 762302 44913 762304
rect 42306 762274 44852 762302
rect 42336 762246 44852 762274
rect 44908 762246 44913 762302
rect 42336 762244 44913 762246
rect 44847 762241 44913 762244
rect 674754 761904 674814 762390
rect 42106 761798 42112 761862
rect 42176 761860 42182 761862
rect 43215 761860 43281 761863
rect 42176 761858 43281 761860
rect 42176 761802 43220 761858
rect 43276 761802 43281 761858
rect 42176 761800 43281 761802
rect 42176 761798 42182 761800
rect 43215 761797 43281 761800
rect 675514 761650 675520 761714
rect 675584 761650 675590 761714
rect 675522 761090 675582 761650
rect 674362 760244 674368 760308
rect 674432 760306 674438 760308
rect 674432 760246 674784 760306
rect 674432 760244 674438 760246
rect 35919 760232 35985 760235
rect 40954 760232 40960 760234
rect 35919 760230 40960 760232
rect 35919 760174 35924 760230
rect 35980 760174 40960 760230
rect 35919 760172 40960 760174
rect 35919 760169 35985 760172
rect 40954 760170 40960 760172
rect 41024 760170 41030 760234
rect 674938 760022 674944 760086
rect 675008 760022 675014 760086
rect 37359 759640 37425 759643
rect 40378 759640 40384 759642
rect 37359 759638 40384 759640
rect 37359 759582 37364 759638
rect 37420 759582 40384 759638
rect 37359 759580 40384 759582
rect 37359 759577 37425 759580
rect 40378 759578 40384 759580
rect 40448 759578 40454 759642
rect 674946 759462 675006 760022
rect 675322 759134 675328 759198
rect 675392 759134 675398 759198
rect 675330 758722 675390 759134
rect 38799 758604 38865 758607
rect 41146 758604 41152 758606
rect 38799 758602 41152 758604
rect 38799 758546 38804 758602
rect 38860 758546 41152 758602
rect 38799 758544 41152 758546
rect 38799 758541 38865 758544
rect 41146 758542 41152 758544
rect 41216 758542 41222 758606
rect 675706 758542 675712 758606
rect 675776 758542 675782 758606
rect 675714 757982 675774 758542
rect 58191 757568 58257 757571
rect 58191 757566 64416 757568
rect 58191 757510 58196 757566
rect 58252 757510 64416 757566
rect 58191 757508 64416 757510
rect 58191 757505 58257 757508
rect 676666 757358 676672 757422
rect 676736 757358 676742 757422
rect 42159 757124 42225 757127
rect 42298 757124 42304 757126
rect 42159 757122 42304 757124
rect 42159 757066 42164 757122
rect 42220 757066 42304 757122
rect 42159 757064 42304 757066
rect 42159 757061 42225 757064
rect 42298 757062 42304 757064
rect 42368 757062 42374 757126
rect 676674 757094 676734 757358
rect 674554 756914 674560 756978
rect 674624 756976 674630 756978
rect 674624 756916 674814 756976
rect 674624 756914 674630 756916
rect 674754 756354 674814 756916
rect 674170 755434 674176 755498
rect 674240 755496 674246 755498
rect 674240 755436 674784 755496
rect 674240 755434 674246 755436
rect 675130 755286 675136 755350
rect 675200 755286 675206 755350
rect 41146 754842 41152 754906
rect 41216 754904 41222 754906
rect 41871 754904 41937 754907
rect 41216 754902 41937 754904
rect 41216 754846 41876 754902
rect 41932 754846 41937 754902
rect 41216 754844 41937 754846
rect 41216 754842 41222 754844
rect 41871 754841 41937 754844
rect 675138 754726 675198 755286
rect 677242 754398 677248 754462
rect 677312 754398 677318 754462
rect 42298 754250 42304 754314
rect 42368 754312 42374 754314
rect 42447 754312 42513 754315
rect 42368 754310 42513 754312
rect 42368 754254 42452 754310
rect 42508 754254 42513 754310
rect 42368 754252 42513 754254
rect 42368 754250 42374 754252
rect 42447 754249 42513 754252
rect 677250 753986 677310 754398
rect 676858 753806 676864 753870
rect 676928 753806 676934 753870
rect 676866 753246 676926 753806
rect 677818 752918 677824 752982
rect 677888 752918 677894 752982
rect 677826 752358 677886 752918
rect 649839 752092 649905 752095
rect 649794 752090 649905 752092
rect 649794 752034 649844 752090
rect 649900 752034 649905 752090
rect 649794 752029 649905 752034
rect 42682 751882 42688 751946
rect 42752 751944 42758 751946
rect 42831 751944 42897 751947
rect 42752 751942 42897 751944
rect 42752 751886 42836 751942
rect 42892 751886 42897 751942
rect 42752 751884 42897 751886
rect 42752 751882 42758 751884
rect 42831 751881 42897 751884
rect 42735 751650 42801 751651
rect 42682 751586 42688 751650
rect 42752 751648 42801 751650
rect 42752 751646 42844 751648
rect 42796 751590 42844 751646
rect 649794 751618 649854 752029
rect 673647 751648 673713 751651
rect 673647 751646 674784 751648
rect 42752 751588 42844 751590
rect 673647 751590 673652 751646
rect 673708 751590 674784 751646
rect 673647 751588 674784 751590
rect 42752 751586 42801 751588
rect 42735 751585 42801 751586
rect 673647 751585 673713 751588
rect 679746 750171 679806 750730
rect 679746 750166 679857 750171
rect 679746 750110 679796 750166
rect 679852 750110 679857 750166
rect 679746 750108 679857 750110
rect 679791 750105 679857 750108
rect 679791 749576 679857 749579
rect 679746 749574 679857 749576
rect 679746 749518 679796 749574
rect 679852 749518 679857 749574
rect 679746 749513 679857 749518
rect 679746 749250 679806 749513
rect 41775 748690 41841 748691
rect 41722 748626 41728 748690
rect 41792 748688 41841 748690
rect 41792 748686 41884 748688
rect 41836 748630 41884 748686
rect 41792 748628 41884 748630
rect 41792 748626 41841 748628
rect 41775 748625 41841 748626
rect 41967 747358 42033 747359
rect 41914 747294 41920 747358
rect 41984 747356 42033 747358
rect 41984 747354 42076 747356
rect 42028 747298 42076 747354
rect 41984 747296 42076 747298
rect 41984 747294 42033 747296
rect 41967 747293 42033 747294
rect 40378 747146 40384 747210
rect 40448 747208 40454 747210
rect 42831 747208 42897 747211
rect 40448 747206 42897 747208
rect 40448 747150 42836 747206
rect 42892 747150 42897 747206
rect 40448 747148 42897 747150
rect 40448 747146 40454 747148
rect 42831 747145 42897 747148
rect 40954 746850 40960 746914
rect 41024 746912 41030 746914
rect 42927 746912 42993 746915
rect 41024 746910 42993 746912
rect 41024 746854 42932 746910
rect 42988 746854 42993 746910
rect 41024 746852 42993 746854
rect 41024 746850 41030 746852
rect 42927 746849 42993 746852
rect 674362 743298 674368 743362
rect 674432 743360 674438 743362
rect 675087 743360 675153 743363
rect 674432 743358 675153 743360
rect 674432 743302 675092 743358
rect 675148 743302 675153 743358
rect 674432 743300 675153 743302
rect 674432 743298 674438 743300
rect 675087 743297 675153 743300
rect 58575 743212 58641 743215
rect 58575 743210 64416 743212
rect 58575 743154 58580 743210
rect 58636 743154 64416 743210
rect 58575 743152 64416 743154
rect 58575 743149 58641 743152
rect 675759 741732 675825 741735
rect 676666 741732 676672 741734
rect 675759 741730 676672 741732
rect 675759 741674 675764 741730
rect 675820 741674 676672 741730
rect 675759 741672 676672 741674
rect 675759 741669 675825 741672
rect 676666 741670 676672 741672
rect 676736 741670 676742 741734
rect 674170 741374 674176 741438
rect 674240 741436 674246 741438
rect 675087 741436 675153 741439
rect 674240 741434 675153 741436
rect 674240 741378 675092 741434
rect 675148 741378 675153 741434
rect 674240 741376 675153 741378
rect 674240 741374 674246 741376
rect 675087 741373 675153 741376
rect 675471 740402 675537 740403
rect 675471 740398 675520 740402
rect 675584 740400 675590 740402
rect 675471 740342 675476 740398
rect 675471 740338 675520 740342
rect 675584 740340 675628 740400
rect 675584 740338 675590 740340
rect 675471 740337 675537 740338
rect 654447 739808 654513 739811
rect 650208 739806 654513 739808
rect 650208 739750 654452 739806
rect 654508 739750 654513 739806
rect 650208 739748 654513 739750
rect 654447 739745 654513 739748
rect 674746 739302 674752 739366
rect 674816 739364 674822 739366
rect 675471 739364 675537 739367
rect 674816 739362 675537 739364
rect 674816 739306 675476 739362
rect 675532 739306 675537 739362
rect 674816 739304 675537 739306
rect 674816 739302 674822 739304
rect 675471 739301 675537 739304
rect 675375 738626 675441 738627
rect 675322 738624 675328 738626
rect 675284 738564 675328 738624
rect 675392 738622 675441 738626
rect 675436 738566 675441 738622
rect 675322 738562 675328 738564
rect 675392 738562 675441 738566
rect 675375 738561 675441 738562
rect 42639 737292 42705 737295
rect 42336 737290 42705 737292
rect 42336 737234 42644 737290
rect 42700 737234 42705 737290
rect 42336 737232 42705 737234
rect 42639 737229 42705 737232
rect 42351 736700 42417 736703
rect 42306 736698 42417 736700
rect 42306 736642 42356 736698
rect 42412 736642 42417 736698
rect 42306 736637 42417 736642
rect 675759 736700 675825 736703
rect 676474 736700 676480 736702
rect 675759 736698 676480 736700
rect 675759 736642 675764 736698
rect 675820 736642 676480 736698
rect 675759 736640 676480 736642
rect 675759 736637 675825 736640
rect 676474 736638 676480 736640
rect 676544 736638 676550 736702
rect 42306 736522 42366 736637
rect 42306 735519 42366 735634
rect 42306 735514 42417 735519
rect 42306 735458 42356 735514
rect 42412 735458 42417 735514
rect 42306 735456 42417 735458
rect 42351 735453 42417 735456
rect 43215 734924 43281 734927
rect 42336 734922 43281 734924
rect 42336 734866 43220 734922
rect 43276 734866 43281 734922
rect 42336 734864 43281 734866
rect 43215 734861 43281 734864
rect 675663 734482 675729 734483
rect 675663 734478 675712 734482
rect 675776 734480 675782 734482
rect 675663 734422 675668 734478
rect 675663 734418 675712 734422
rect 675776 734420 675820 734480
rect 675776 734418 675782 734420
rect 675663 734417 675729 734418
rect 43407 734036 43473 734039
rect 42336 734034 43473 734036
rect 42336 733978 43412 734034
rect 43468 733978 43473 734034
rect 42336 733976 43473 733978
rect 43407 733973 43473 733976
rect 41722 733826 41728 733890
rect 41792 733826 41798 733890
rect 41730 733370 41790 733826
rect 40608 733340 41790 733370
rect 40578 733310 41760 733340
rect 40578 733150 40638 733310
rect 40570 733086 40576 733150
rect 40640 733086 40646 733150
rect 40762 733086 40768 733150
rect 40832 733086 40838 733150
rect 40770 732556 40830 733086
rect 675183 732556 675249 732559
rect 676858 732556 676864 732558
rect 40770 732526 41184 732556
rect 675183 732554 676864 732556
rect 40800 732496 41214 732526
rect 41154 732262 41214 732496
rect 675183 732498 675188 732554
rect 675244 732498 676864 732554
rect 675183 732496 676864 732498
rect 675183 732493 675249 732496
rect 676858 732494 676864 732496
rect 676928 732494 676934 732558
rect 41146 732198 41152 732262
rect 41216 732198 41222 732262
rect 42306 731668 42366 731712
rect 42927 731668 42993 731671
rect 42306 731666 42993 731668
rect 42306 731610 42932 731666
rect 42988 731610 42993 731666
rect 42306 731608 42993 731610
rect 42927 731605 42993 731608
rect 40194 730339 40254 730898
rect 40194 730334 40305 730339
rect 40194 730278 40244 730334
rect 40300 730278 40305 730334
rect 40194 730276 40305 730278
rect 40239 730273 40305 730276
rect 41346 729598 41406 730084
rect 41338 729534 41344 729598
rect 41408 729534 41414 729598
rect 41538 728859 41598 729270
rect 41538 728854 41649 728859
rect 41538 728798 41588 728854
rect 41644 728798 41649 728854
rect 41538 728796 41649 728798
rect 41583 728793 41649 728796
rect 59535 728856 59601 728859
rect 59535 728854 64416 728856
rect 59535 728798 59540 728854
rect 59596 728798 64416 728854
rect 59535 728796 64416 728798
rect 59535 728793 59601 728796
rect 41730 727971 41790 728530
rect 655119 728116 655185 728119
rect 650208 728114 655185 728116
rect 650208 728058 655124 728114
rect 655180 728058 655185 728114
rect 650208 728056 655185 728058
rect 655119 728053 655185 728056
rect 41730 727966 41841 727971
rect 41730 727910 41780 727966
rect 41836 727910 41841 727966
rect 41730 727908 41841 727910
rect 41775 727905 41841 727908
rect 41538 727231 41598 727790
rect 41487 727226 41598 727231
rect 41487 727170 41492 727226
rect 41548 727170 41598 727226
rect 41487 727168 41598 727170
rect 41487 727165 41553 727168
rect 40962 726342 41022 726902
rect 40954 726278 40960 726342
rect 41024 726278 41030 726342
rect 41730 725899 41790 726162
rect 41679 725894 41790 725899
rect 41679 725838 41684 725894
rect 41740 725838 41790 725894
rect 41679 725836 41790 725838
rect 41679 725833 41745 725836
rect 42114 724715 42174 725274
rect 42063 724710 42174 724715
rect 42063 724654 42068 724710
rect 42124 724654 42174 724710
rect 42063 724652 42174 724654
rect 42063 724649 42129 724652
rect 42114 724123 42174 724534
rect 42114 724118 42225 724123
rect 42114 724062 42164 724118
rect 42220 724062 42225 724118
rect 42114 724060 42225 724062
rect 42159 724057 42225 724060
rect 41922 723235 41982 723794
rect 41922 723230 42033 723235
rect 41922 723174 41972 723230
rect 42028 723174 42033 723230
rect 41922 723172 42033 723174
rect 41967 723169 42033 723172
rect 43023 723084 43089 723087
rect 42336 723082 43089 723084
rect 42336 723026 43028 723082
rect 43084 723026 43089 723082
rect 42336 723024 43089 723026
rect 43023 723021 43089 723024
rect 674319 722492 674385 722495
rect 674319 722490 674784 722492
rect 674319 722434 674324 722490
rect 674380 722434 674784 722490
rect 674319 722432 674784 722434
rect 674319 722429 674385 722432
rect 42306 721604 42366 722166
rect 674799 721900 674865 721903
rect 674754 721898 674865 721900
rect 674754 721842 674804 721898
rect 674860 721842 674865 721898
rect 674754 721837 674865 721842
rect 674754 721722 674814 721837
rect 42490 721604 42496 721606
rect 42306 721544 42496 721604
rect 42490 721542 42496 721544
rect 42560 721542 42566 721606
rect 43066 721456 43072 721458
rect 42336 721396 43072 721456
rect 43066 721394 43072 721396
rect 43136 721394 43142 721458
rect 674319 720864 674385 720867
rect 674319 720862 674784 720864
rect 674319 720806 674324 720862
rect 674380 720806 674784 720862
rect 674319 720804 674784 720806
rect 674319 720801 674385 720804
rect 42306 719979 42366 720538
rect 674799 720272 674865 720275
rect 674754 720270 674865 720272
rect 674754 720214 674804 720270
rect 674860 720214 674865 720270
rect 674754 720209 674865 720214
rect 674754 720094 674814 720209
rect 42255 719974 42366 719979
rect 42255 719918 42260 719974
rect 42316 719918 42366 719974
rect 42255 719916 42366 719918
rect 42255 719913 42321 719916
rect 674754 719091 674814 719206
rect 674754 719086 674865 719091
rect 42306 718795 42366 719058
rect 674754 719030 674804 719086
rect 674860 719030 674865 719086
rect 674754 719028 674865 719030
rect 674799 719025 674865 719028
rect 42255 718790 42366 718795
rect 42255 718734 42260 718790
rect 42316 718734 42366 718790
rect 42255 718732 42366 718734
rect 42255 718729 42321 718732
rect 679746 718055 679806 718540
rect 679695 718050 679806 718055
rect 679695 717994 679700 718050
rect 679756 717994 679806 718050
rect 679695 717992 679806 717994
rect 679695 717989 679761 717992
rect 674511 717904 674577 717907
rect 674511 717902 674814 717904
rect 674511 717846 674516 717902
rect 674572 717846 674814 717902
rect 674511 717844 674814 717846
rect 674511 717841 674577 717844
rect 674754 717726 674814 717844
rect 675898 717065 675904 717129
rect 675968 717065 675974 717129
rect 675906 716912 675966 717065
rect 654447 716276 654513 716279
rect 650208 716274 654513 716276
rect 650208 716218 654452 716274
rect 654508 716218 654513 716274
rect 650208 716216 654513 716218
rect 654447 716213 654513 716216
rect 675087 716276 675153 716279
rect 675087 716274 675198 716276
rect 675087 716218 675092 716274
rect 675148 716218 675198 716274
rect 675087 716213 675198 716218
rect 41775 716130 41841 716131
rect 41722 716066 41728 716130
rect 41792 716128 41841 716130
rect 41792 716126 41884 716128
rect 41836 716070 41884 716126
rect 675138 716098 675198 716213
rect 41792 716068 41884 716070
rect 41792 716066 41841 716068
rect 41775 716065 41841 716066
rect 676282 715770 676288 715834
rect 676352 715770 676358 715834
rect 676290 715284 676350 715770
rect 674415 714500 674481 714503
rect 674415 714498 674784 714500
rect 674415 714442 674420 714498
rect 674476 714442 674784 714498
rect 674415 714440 674784 714442
rect 674415 714437 674481 714440
rect 59535 714352 59601 714355
rect 59535 714350 64416 714352
rect 59535 714294 59540 714350
rect 59596 714294 64416 714350
rect 59535 714292 64416 714294
rect 59535 714289 59601 714292
rect 41871 714056 41937 714059
rect 42106 714056 42112 714058
rect 41871 714054 42112 714056
rect 41871 713998 41876 714054
rect 41932 713998 42112 714054
rect 41871 713996 42112 713998
rect 41871 713993 41937 713996
rect 42106 713994 42112 713996
rect 42176 713994 42182 714058
rect 42063 713908 42129 713911
rect 42298 713908 42304 713910
rect 42063 713906 42304 713908
rect 42063 713850 42068 713906
rect 42124 713850 42304 713906
rect 42063 713848 42304 713850
rect 42063 713845 42129 713848
rect 42298 713846 42304 713848
rect 42368 713846 42374 713910
rect 674319 713760 674385 713763
rect 674319 713758 674784 713760
rect 674319 713702 674324 713758
rect 674380 713702 674784 713758
rect 674319 713700 674784 713702
rect 674319 713697 674385 713700
rect 674223 713020 674289 713023
rect 674223 713018 674784 713020
rect 674223 712962 674228 713018
rect 674284 712962 674784 713018
rect 674223 712960 674784 712962
rect 674223 712957 674289 712960
rect 673978 712070 673984 712134
rect 674048 712132 674054 712134
rect 674048 712072 674784 712132
rect 674048 712070 674054 712072
rect 676090 711922 676096 711986
rect 676160 711922 676166 711986
rect 42927 711838 42993 711839
rect 42874 711836 42880 711838
rect 42836 711776 42880 711836
rect 42944 711834 42993 711838
rect 42988 711778 42993 711834
rect 42874 711774 42880 711776
rect 42944 711774 42993 711778
rect 42927 711773 42993 711774
rect 42063 711690 42129 711691
rect 42063 711688 42112 711690
rect 42020 711686 42112 711688
rect 42020 711630 42068 711686
rect 42020 711628 42112 711630
rect 42063 711626 42112 711628
rect 42176 711626 42182 711690
rect 42682 711626 42688 711690
rect 42752 711688 42758 711690
rect 43023 711688 43089 711691
rect 42752 711686 43089 711688
rect 42752 711630 43028 711686
rect 43084 711630 43089 711686
rect 42752 711628 43089 711630
rect 42752 711626 42758 711628
rect 42063 711625 42129 711626
rect 43023 711625 43089 711628
rect 41530 711330 41536 711394
rect 41600 711330 41606 711394
rect 676098 711362 676158 711922
rect 41538 711096 41598 711330
rect 42682 711182 42688 711246
rect 42752 711244 42758 711246
rect 43119 711244 43185 711247
rect 42752 711242 43185 711244
rect 42752 711186 43124 711242
rect 43180 711186 43185 711242
rect 42752 711184 43185 711186
rect 42752 711182 42758 711184
rect 43119 711181 43185 711184
rect 41722 711096 41728 711098
rect 41538 711036 41728 711096
rect 41722 711034 41728 711036
rect 41792 711034 41798 711098
rect 42298 711034 42304 711098
rect 42368 711096 42374 711098
rect 42831 711096 42897 711099
rect 42368 711094 42897 711096
rect 42368 711038 42836 711094
rect 42892 711038 42897 711094
rect 42368 711036 42897 711038
rect 42368 711034 42374 711036
rect 42831 711033 42897 711036
rect 674415 710504 674481 710507
rect 674415 710502 674784 710504
rect 674415 710446 674420 710502
rect 674476 710446 674784 710502
rect 674415 710444 674784 710446
rect 674415 710441 674481 710444
rect 674799 709912 674865 709915
rect 674754 709910 674865 709912
rect 674754 709854 674804 709910
rect 674860 709854 674865 709910
rect 674754 709849 674865 709854
rect 674754 709734 674814 709849
rect 674415 709024 674481 709027
rect 674415 709022 674784 709024
rect 674415 708966 674420 709022
rect 674476 708966 674784 709022
rect 674415 708964 674784 708966
rect 674415 708961 674481 708964
rect 42063 708580 42129 708583
rect 43066 708580 43072 708582
rect 42063 708578 43072 708580
rect 42063 708522 42068 708578
rect 42124 708522 43072 708578
rect 42063 708520 43072 708522
rect 42063 708517 42129 708520
rect 43066 708518 43072 708520
rect 43136 708518 43142 708582
rect 677050 708370 677056 708434
rect 677120 708370 677126 708434
rect 677058 708254 677118 708370
rect 42874 707778 42880 707842
rect 42944 707840 42950 707842
rect 43023 707840 43089 707843
rect 42944 707838 43089 707840
rect 42944 707782 43028 707838
rect 43084 707782 43089 707838
rect 42944 707780 43089 707782
rect 42944 707778 42950 707780
rect 43023 707777 43089 707780
rect 42159 707396 42225 707399
rect 42490 707396 42496 707398
rect 42159 707394 42496 707396
rect 42159 707338 42164 707394
rect 42220 707338 42496 707394
rect 42159 707336 42496 707338
rect 42159 707333 42225 707336
rect 42490 707334 42496 707336
rect 42560 707334 42566 707398
rect 674415 707396 674481 707399
rect 674415 707394 674784 707396
rect 674415 707338 674420 707394
rect 674476 707338 674784 707394
rect 674415 707336 674784 707338
rect 674415 707333 674481 707336
rect 674799 706804 674865 706807
rect 674754 706802 674865 706804
rect 674754 706746 674804 706802
rect 674860 706746 674865 706802
rect 674754 706741 674865 706746
rect 674754 706626 674814 706741
rect 41967 706510 42033 706511
rect 41914 706508 41920 706510
rect 41876 706448 41920 706508
rect 41984 706506 42033 706510
rect 42028 706450 42033 706506
rect 41914 706446 41920 706448
rect 41984 706446 42033 706450
rect 41967 706445 42033 706446
rect 650127 705324 650193 705327
rect 650127 705322 650238 705324
rect 650127 705266 650132 705322
rect 650188 705266 650238 705322
rect 650127 705261 650238 705266
rect 41722 704966 41728 705030
rect 41792 704966 41798 705030
rect 41730 704735 41790 704966
rect 41530 704670 41536 704734
rect 41600 704732 41606 704734
rect 41730 704732 41841 704735
rect 41600 704730 41841 704732
rect 41600 704674 41780 704730
rect 41836 704674 41841 704730
rect 650178 704702 650238 705261
rect 679746 705179 679806 705738
rect 679746 705174 679857 705179
rect 679746 705118 679796 705174
rect 679852 705118 679857 705174
rect 679746 705116 679857 705118
rect 679791 705113 679857 705116
rect 41600 704672 41841 704674
rect 41600 704670 41606 704672
rect 41775 704669 41841 704672
rect 679791 704584 679857 704587
rect 679746 704582 679857 704584
rect 679746 704526 679796 704582
rect 679852 704526 679857 704582
rect 679746 704521 679857 704526
rect 679746 704258 679806 704521
rect 42063 704142 42129 704143
rect 42063 704140 42112 704142
rect 42020 704138 42112 704140
rect 42020 704082 42068 704138
rect 42020 704080 42112 704082
rect 42063 704078 42112 704080
rect 42176 704078 42182 704142
rect 42063 704077 42129 704078
rect 41338 703634 41344 703698
rect 41408 703696 41414 703698
rect 42255 703696 42321 703699
rect 41408 703694 42321 703696
rect 41408 703638 42260 703694
rect 42316 703638 42321 703694
rect 41408 703636 42321 703638
rect 41408 703634 41414 703636
rect 42255 703633 42321 703636
rect 40954 703486 40960 703550
rect 41024 703548 41030 703550
rect 42831 703548 42897 703551
rect 41024 703546 42897 703548
rect 41024 703490 42836 703546
rect 42892 703490 42897 703546
rect 41024 703488 42897 703490
rect 41024 703486 41030 703488
rect 42831 703485 42897 703488
rect 42255 700884 42321 700887
rect 42255 700882 42366 700884
rect 42255 700826 42260 700882
rect 42316 700826 42366 700882
rect 42255 700821 42366 700826
rect 42306 700591 42366 700821
rect 42255 700586 42366 700591
rect 42255 700530 42260 700586
rect 42316 700530 42366 700586
rect 42255 700528 42366 700530
rect 42255 700525 42321 700528
rect 59535 700144 59601 700147
rect 59535 700142 64416 700144
rect 59535 700086 59540 700142
rect 59596 700086 64416 700142
rect 59535 700084 64416 700086
rect 59535 700081 59601 700084
rect 675130 697862 675136 697926
rect 675200 697924 675206 697926
rect 675375 697924 675441 697927
rect 675200 697922 675441 697924
rect 675200 697866 675380 697922
rect 675436 697866 675441 697922
rect 675200 697864 675441 697866
rect 675200 697862 675206 697864
rect 675375 697861 675441 697864
rect 673978 697270 673984 697334
rect 674048 697332 674054 697334
rect 675471 697332 675537 697335
rect 674048 697330 675537 697332
rect 674048 697274 675476 697330
rect 675532 697274 675537 697330
rect 674048 697272 675537 697274
rect 674048 697270 674054 697272
rect 675471 697269 675537 697272
rect 674938 696826 674944 696890
rect 675008 696888 675014 696890
rect 675375 696888 675441 696891
rect 675008 696886 675441 696888
rect 675008 696830 675380 696886
rect 675436 696830 675441 696886
rect 675008 696828 675441 696830
rect 675008 696826 675014 696828
rect 675375 696825 675441 696828
rect 675759 694816 675825 694819
rect 676090 694816 676096 694818
rect 675759 694814 676096 694816
rect 675759 694758 675764 694814
rect 675820 694758 676096 694814
rect 675759 694756 676096 694758
rect 675759 694753 675825 694756
rect 676090 694754 676096 694756
rect 676160 694754 676166 694818
rect 674554 694606 674560 694670
rect 674624 694668 674630 694670
rect 675279 694668 675345 694671
rect 674624 694666 675345 694668
rect 674624 694610 675284 694666
rect 675340 694610 675345 694666
rect 674624 694608 675345 694610
rect 674624 694606 674630 694608
rect 675279 694605 675345 694608
rect 42639 694076 42705 694079
rect 42336 694074 42705 694076
rect 42336 694018 42644 694074
rect 42700 694018 42705 694074
rect 42336 694016 42705 694018
rect 42639 694013 42705 694016
rect 42351 693484 42417 693487
rect 42306 693482 42417 693484
rect 42306 693426 42356 693482
rect 42412 693426 42417 693482
rect 42306 693421 42417 693426
rect 675759 693484 675825 693487
rect 675898 693484 675904 693486
rect 675759 693482 675904 693484
rect 675759 693426 675764 693482
rect 675820 693426 675904 693482
rect 675759 693424 675904 693426
rect 675759 693421 675825 693424
rect 675898 693422 675904 693424
rect 675968 693422 675974 693486
rect 42306 693306 42366 693421
rect 654831 692892 654897 692895
rect 650208 692890 654897 692892
rect 650208 692834 654836 692890
rect 654892 692834 654897 692890
rect 650208 692832 654897 692834
rect 654831 692829 654897 692832
rect 41391 692744 41457 692747
rect 41530 692744 41536 692746
rect 41391 692742 41536 692744
rect 41391 692686 41396 692742
rect 41452 692686 41536 692742
rect 41391 692684 41536 692686
rect 41391 692681 41457 692684
rect 41530 692682 41536 692684
rect 41600 692682 41606 692746
rect 42639 692448 42705 692451
rect 42336 692446 42705 692448
rect 42336 692390 42644 692446
rect 42700 692390 42705 692446
rect 42336 692388 42705 692390
rect 42639 692385 42705 692388
rect 43407 691708 43473 691711
rect 42336 691706 43473 691708
rect 42336 691650 43412 691706
rect 43468 691650 43473 691706
rect 42336 691648 43473 691650
rect 43407 691645 43473 691648
rect 675759 691708 675825 691711
rect 676474 691708 676480 691710
rect 675759 691706 676480 691708
rect 675759 691650 675764 691706
rect 675820 691650 676480 691706
rect 675759 691648 676480 691650
rect 675759 691645 675825 691648
rect 676474 691646 676480 691648
rect 676544 691646 676550 691710
rect 43215 690820 43281 690823
rect 42336 690818 43281 690820
rect 42336 690762 43220 690818
rect 43276 690762 43281 690818
rect 42336 690760 43281 690762
rect 43215 690757 43281 690760
rect 40578 689638 40638 690198
rect 40570 689574 40576 689638
rect 40640 689574 40646 689638
rect 41146 689574 41152 689638
rect 41216 689574 41222 689638
rect 41154 689340 41214 689574
rect 674799 689340 674865 689343
rect 676666 689340 676672 689342
rect 41154 689310 42144 689340
rect 674799 689338 676672 689340
rect 41184 689280 42174 689310
rect 42114 688750 42174 689280
rect 674799 689282 674804 689338
rect 674860 689282 676672 689338
rect 674799 689280 676672 689282
rect 674799 689277 674865 689280
rect 676666 689278 676672 689280
rect 676736 689278 676742 689342
rect 675759 689192 675825 689195
rect 676666 689192 676672 689194
rect 675759 689190 676672 689192
rect 675759 689134 675764 689190
rect 675820 689134 676672 689190
rect 675759 689132 676672 689134
rect 675759 689129 675825 689132
rect 676666 689130 676672 689132
rect 676736 689130 676742 689194
rect 42106 688686 42112 688750
rect 42176 688686 42182 688750
rect 41538 688307 41598 688496
rect 41538 688302 41649 688307
rect 41538 688246 41588 688302
rect 41644 688246 41649 688302
rect 41538 688244 41649 688246
rect 41583 688241 41649 688244
rect 674895 688304 674961 688307
rect 677050 688304 677056 688306
rect 674895 688302 677056 688304
rect 674895 688246 674900 688302
rect 674956 688246 677056 688302
rect 674895 688244 677056 688246
rect 674895 688241 674961 688244
rect 677050 688242 677056 688244
rect 677120 688242 677126 688306
rect 40194 687123 40254 687682
rect 40194 687118 40305 687123
rect 40194 687062 40244 687118
rect 40300 687062 40305 687118
rect 40194 687060 40305 687062
rect 40239 687057 40305 687060
rect 41154 686382 41214 686868
rect 41146 686318 41152 686382
rect 41216 686318 41222 686382
rect 41730 685643 41790 686054
rect 41679 685638 41790 685643
rect 41679 685582 41684 685638
rect 41740 685582 41790 685638
rect 41679 685580 41790 685582
rect 58671 685640 58737 685643
rect 675087 685640 675153 685643
rect 677050 685640 677056 685642
rect 58671 685638 64416 685640
rect 58671 685582 58676 685638
rect 58732 685582 64416 685638
rect 58671 685580 64416 685582
rect 675087 685638 677056 685640
rect 675087 685582 675092 685638
rect 675148 685582 677056 685638
rect 675087 685580 677056 685582
rect 41679 685577 41745 685580
rect 58671 685577 58737 685580
rect 675087 685577 675153 685580
rect 677050 685578 677056 685580
rect 677120 685578 677126 685642
rect 42306 684900 42366 685388
rect 42490 684900 42496 684902
rect 42306 684840 42496 684900
rect 42490 684838 42496 684840
rect 42560 684838 42566 684902
rect 41730 684015 41790 684574
rect 41730 684010 41841 684015
rect 41730 683954 41780 684010
rect 41836 683954 41841 684010
rect 41730 683952 41841 683954
rect 41775 683949 41841 683952
rect 40962 683274 41022 683760
rect 40954 683210 40960 683274
rect 41024 683210 41030 683274
rect 42874 682976 42880 682978
rect 42336 682916 42880 682976
rect 42874 682914 42880 682916
rect 42944 682914 42950 682978
rect 41922 681499 41982 682058
rect 41871 681494 41982 681499
rect 41871 681438 41876 681494
rect 41932 681438 41982 681494
rect 41871 681436 41982 681438
rect 41871 681433 41937 681436
rect 41922 680907 41982 681318
rect 655311 681200 655377 681203
rect 650208 681198 655377 681200
rect 650208 681142 655316 681198
rect 655372 681142 655377 681198
rect 650208 681140 655377 681142
rect 655311 681137 655377 681140
rect 41922 680902 42033 680907
rect 41922 680846 41972 680902
rect 42028 680846 42033 680902
rect 41922 680844 42033 680846
rect 41967 680841 42033 680844
rect 42306 680019 42366 680578
rect 42255 680014 42366 680019
rect 42255 679958 42260 680014
rect 42316 679958 42366 680014
rect 42255 679956 42366 679958
rect 42255 679953 42321 679956
rect 43599 679868 43665 679871
rect 42336 679866 43665 679868
rect 42336 679810 43604 679866
rect 43660 679810 43665 679866
rect 42336 679808 43665 679810
rect 43599 679805 43665 679808
rect 674799 679720 674865 679723
rect 676282 679720 676288 679722
rect 674799 679718 676288 679720
rect 674799 679662 674804 679718
rect 674860 679662 676288 679718
rect 674799 679660 676288 679662
rect 674799 679657 674865 679660
rect 676282 679658 676288 679660
rect 676352 679658 676358 679722
rect 42306 678390 42366 678950
rect 42298 678326 42304 678390
rect 42368 678326 42374 678390
rect 43119 678240 43185 678243
rect 42336 678238 43185 678240
rect 42336 678182 43124 678238
rect 43180 678182 43185 678238
rect 42336 678180 43185 678182
rect 43119 678177 43185 678180
rect 674799 677500 674865 677503
rect 674754 677498 674865 677500
rect 674754 677442 674804 677498
rect 674860 677442 674865 677498
rect 674754 677437 674865 677442
rect 674754 677322 674814 677437
rect 42306 677207 42366 677322
rect 42306 677202 42417 677207
rect 42306 677146 42356 677202
rect 42412 677146 42417 677202
rect 42306 677144 42417 677146
rect 42351 677141 42417 677144
rect 674415 676464 674481 676467
rect 674415 676462 674784 676464
rect 674415 676406 674420 676462
rect 674476 676406 674784 676462
rect 674415 676404 674784 676406
rect 674415 676401 674481 676404
rect 674799 675872 674865 675875
rect 674754 675870 674865 675872
rect 42306 675727 42366 675842
rect 674754 675814 674804 675870
rect 674860 675814 674865 675870
rect 674754 675809 674865 675814
rect 42306 675722 42417 675727
rect 42306 675666 42356 675722
rect 42412 675666 42417 675722
rect 674754 675694 674814 675809
rect 42306 675664 42417 675666
rect 42351 675661 42417 675664
rect 41391 674838 41457 674839
rect 41338 674836 41344 674838
rect 41300 674776 41344 674836
rect 41408 674834 41457 674838
rect 41452 674778 41457 674834
rect 41338 674774 41344 674776
rect 41408 674774 41457 674778
rect 41391 674773 41457 674774
rect 674415 674836 674481 674839
rect 674415 674834 674784 674836
rect 674415 674778 674420 674834
rect 674476 674778 674784 674834
rect 674415 674776 674784 674778
rect 674415 674773 674481 674776
rect 674415 674096 674481 674099
rect 674415 674094 674784 674096
rect 674415 674038 674420 674094
rect 674476 674038 674784 674094
rect 674415 674036 674784 674038
rect 674415 674033 674481 674036
rect 674754 673211 674814 673326
rect 674754 673206 674865 673211
rect 674754 673150 674804 673206
rect 674860 673150 674865 673206
rect 674754 673148 674865 673150
rect 674799 673145 674865 673148
rect 675138 672323 675198 672512
rect 675087 672318 675198 672323
rect 675087 672262 675092 672318
rect 675148 672262 675198 672318
rect 675087 672260 675198 672262
rect 675087 672257 675153 672260
rect 676282 672258 676288 672322
rect 676352 672258 676358 672322
rect 676290 671698 676350 672258
rect 58383 671432 58449 671435
rect 58383 671430 64416 671432
rect 58383 671374 58388 671430
rect 58444 671374 64416 671430
rect 58383 671372 64416 671374
rect 58383 671369 58449 671372
rect 674703 671136 674769 671139
rect 674703 671134 674814 671136
rect 674703 671078 674708 671134
rect 674764 671078 674814 671134
rect 674703 671073 674814 671078
rect 41007 670988 41073 670991
rect 42639 670990 42705 670991
rect 43023 670990 43089 670991
rect 41722 670988 41728 670990
rect 41007 670986 41728 670988
rect 41007 670930 41012 670986
rect 41068 670930 41728 670986
rect 41007 670928 41728 670930
rect 41007 670925 41073 670928
rect 41722 670926 41728 670928
rect 41792 670926 41798 670990
rect 42639 670986 42688 670990
rect 42752 670988 42758 670990
rect 42639 670930 42644 670986
rect 42639 670926 42688 670930
rect 42752 670928 42796 670988
rect 43023 670986 43072 670990
rect 43136 670988 43142 670990
rect 43023 670930 43028 670986
rect 42752 670926 42758 670928
rect 43023 670926 43072 670930
rect 43136 670928 43180 670988
rect 43136 670926 43142 670928
rect 42639 670925 42705 670926
rect 43023 670925 43089 670926
rect 674754 670884 674814 671073
rect 674362 670038 674368 670102
rect 674432 670100 674438 670102
rect 674432 670040 674784 670100
rect 674432 670038 674438 670040
rect 675514 669742 675520 669806
rect 675584 669742 675590 669806
rect 654447 669360 654513 669363
rect 650208 669358 654513 669360
rect 650208 669302 654452 669358
rect 654508 669302 654513 669358
rect 650208 669300 654513 669302
rect 654447 669297 654513 669300
rect 675522 669256 675582 669742
rect 42543 668918 42609 668919
rect 42490 668854 42496 668918
rect 42560 668916 42609 668918
rect 42560 668914 42652 668916
rect 42604 668858 42652 668914
rect 42560 668856 42652 668858
rect 42560 668854 42609 668856
rect 42543 668853 42609 668854
rect 674127 668620 674193 668623
rect 674127 668618 674784 668620
rect 674127 668562 674132 668618
rect 674188 668562 674784 668618
rect 674127 668560 674784 668562
rect 674127 668557 674193 668560
rect 41775 668474 41841 668475
rect 41722 668472 41728 668474
rect 41684 668412 41728 668472
rect 41792 668470 41841 668474
rect 41836 668414 41841 668470
rect 41722 668410 41728 668412
rect 41792 668410 41841 668414
rect 41775 668409 41841 668410
rect 42298 668262 42304 668326
rect 42368 668324 42374 668326
rect 43119 668324 43185 668327
rect 42368 668322 43185 668324
rect 42368 668266 43124 668322
rect 43180 668266 43185 668322
rect 42368 668264 43185 668266
rect 42368 668262 42374 668264
rect 43119 668261 43185 668264
rect 674607 668028 674673 668031
rect 674607 668026 674814 668028
rect 674607 667970 674612 668026
rect 674668 667970 674814 668026
rect 674607 667968 674814 667970
rect 674607 667965 674673 667968
rect 674754 667776 674814 667968
rect 674170 666930 674176 666994
rect 674240 666992 674246 666994
rect 674240 666932 674784 666992
rect 674240 666930 674246 666932
rect 674746 666634 674752 666698
rect 674816 666634 674822 666698
rect 42927 666550 42993 666551
rect 42874 666486 42880 666550
rect 42944 666548 42993 666550
rect 42944 666546 43036 666548
rect 42988 666490 43036 666546
rect 42944 666488 43036 666490
rect 42944 666486 42993 666488
rect 42927 666485 42993 666486
rect 674754 666074 674814 666634
rect 675322 665894 675328 665958
rect 675392 665894 675398 665958
rect 41338 665746 41344 665810
rect 41408 665746 41414 665810
rect 41346 665662 41406 665746
rect 41338 665598 41344 665662
rect 41408 665598 41414 665662
rect 42159 665364 42225 665367
rect 43066 665364 43072 665366
rect 42159 665362 43072 665364
rect 42159 665306 42164 665362
rect 42220 665306 43072 665362
rect 42159 665304 43072 665306
rect 42159 665301 42225 665304
rect 43066 665302 43072 665304
rect 43136 665302 43142 665366
rect 675330 665334 675390 665894
rect 674991 664772 675057 664775
rect 674946 664770 675057 664772
rect 674946 664714 674996 664770
rect 675052 664714 675057 664770
rect 674946 664709 675057 664714
rect 674946 664446 675006 664709
rect 675706 664266 675712 664330
rect 675776 664266 675782 664330
rect 675714 663854 675774 664266
rect 677242 663526 677248 663590
rect 677312 663526 677318 663590
rect 42543 663440 42609 663443
rect 42682 663440 42688 663442
rect 42543 663438 42688 663440
rect 42543 663382 42548 663438
rect 42604 663382 42688 663438
rect 42543 663380 42688 663382
rect 42543 663377 42609 663380
rect 42682 663378 42688 663380
rect 42752 663378 42758 663442
rect 677250 662966 677310 663526
rect 676858 662342 676864 662406
rect 676928 662342 676934 662406
rect 676866 662226 676926 662342
rect 674703 661664 674769 661667
rect 674703 661662 674814 661664
rect 674703 661606 674708 661662
rect 674764 661606 674814 661662
rect 674703 661601 674814 661606
rect 41775 661370 41841 661371
rect 41338 661306 41344 661370
rect 41408 661368 41414 661370
rect 41722 661368 41728 661370
rect 41408 661308 41728 661368
rect 41792 661368 41841 661370
rect 41792 661366 41884 661368
rect 41836 661310 41884 661366
rect 674754 661338 674814 661601
rect 41408 661306 41414 661308
rect 41722 661306 41728 661308
rect 41792 661308 41884 661310
rect 41792 661306 41841 661308
rect 41775 661305 41841 661306
rect 41871 661074 41937 661075
rect 41871 661072 41920 661074
rect 41828 661070 41920 661072
rect 41828 661014 41876 661070
rect 41828 661012 41920 661014
rect 41871 661010 41920 661012
rect 41984 661010 41990 661074
rect 41871 661009 41937 661010
rect 40954 660862 40960 660926
rect 41024 660924 41030 660926
rect 42831 660924 42897 660927
rect 41024 660922 42897 660924
rect 41024 660866 42836 660922
rect 42892 660866 42897 660922
rect 41024 660864 42897 660866
rect 41024 660862 41030 660864
rect 42831 660861 42897 660864
rect 679746 660039 679806 660598
rect 679746 660034 679857 660039
rect 679746 659978 679796 660034
rect 679852 659978 679857 660034
rect 679746 659976 679857 659978
rect 679791 659973 679857 659976
rect 675706 659382 675712 659446
rect 675776 659444 675782 659446
rect 676666 659444 676672 659446
rect 675776 659384 676672 659444
rect 675776 659382 675782 659384
rect 676666 659382 676672 659384
rect 676736 659382 676742 659446
rect 675514 659234 675520 659298
rect 675584 659296 675590 659298
rect 676474 659296 676480 659298
rect 675584 659236 676480 659296
rect 675584 659234 675590 659236
rect 676474 659234 676480 659236
rect 676544 659234 676550 659298
rect 679791 659296 679857 659299
rect 679746 659294 679857 659296
rect 679746 659238 679796 659294
rect 679852 659238 679857 659294
rect 679746 659233 679857 659238
rect 679746 659118 679806 659233
rect 653775 658408 653841 658411
rect 650178 658406 653841 658408
rect 650178 658350 653780 658406
rect 653836 658350 653841 658406
rect 650178 658348 653841 658350
rect 650178 657786 650238 658348
rect 653775 658345 653841 658348
rect 59535 656928 59601 656931
rect 59535 656926 64416 656928
rect 59535 656870 59540 656926
rect 59596 656870 64416 656926
rect 59535 656868 64416 656870
rect 59535 656865 59601 656868
rect 41146 656126 41152 656190
rect 41216 656188 41222 656190
rect 41775 656188 41841 656191
rect 41216 656186 41841 656188
rect 41216 656130 41780 656186
rect 41836 656130 41841 656186
rect 41216 656128 41841 656130
rect 41216 656126 41222 656128
rect 41775 656125 41841 656128
rect 674991 652784 675057 652787
rect 675514 652784 675520 652786
rect 674991 652782 675520 652784
rect 674991 652726 674996 652782
rect 675052 652726 675520 652782
rect 674991 652724 675520 652726
rect 674991 652721 675057 652724
rect 675514 652722 675520 652724
rect 675584 652722 675590 652786
rect 675471 652638 675537 652639
rect 675471 652634 675520 652638
rect 675584 652636 675590 652638
rect 675471 652578 675476 652634
rect 675471 652574 675520 652578
rect 675584 652576 675628 652636
rect 675584 652574 675590 652576
rect 675471 652573 675537 652574
rect 674746 652130 674752 652194
rect 674816 652192 674822 652194
rect 675471 652192 675537 652195
rect 674816 652190 675537 652192
rect 674816 652134 675476 652190
rect 675532 652134 675537 652190
rect 674816 652132 675537 652134
rect 674816 652130 674822 652132
rect 675471 652129 675537 652132
rect 675279 651010 675345 651011
rect 675279 651006 675328 651010
rect 675392 651008 675398 651010
rect 675279 650950 675284 651006
rect 675279 650946 675328 650950
rect 675392 650948 675436 651008
rect 675392 650946 675398 650948
rect 675279 650945 675345 650946
rect 42831 650860 42897 650863
rect 42336 650858 42897 650860
rect 42336 650802 42836 650858
rect 42892 650802 42897 650858
rect 42336 650800 42897 650802
rect 42831 650797 42897 650800
rect 42306 649824 42366 650090
rect 42447 649824 42513 649827
rect 42306 649822 42513 649824
rect 42306 649766 42452 649822
rect 42508 649766 42513 649822
rect 42306 649764 42513 649766
rect 42447 649761 42513 649764
rect 675759 649676 675825 649679
rect 676282 649676 676288 649678
rect 675759 649674 676288 649676
rect 675759 649618 675764 649674
rect 675820 649618 676288 649674
rect 675759 649616 676288 649618
rect 675759 649613 675825 649616
rect 676282 649614 676288 649616
rect 676352 649614 676358 649678
rect 42447 649528 42513 649531
rect 42306 649526 42513 649528
rect 42306 649470 42452 649526
rect 42508 649470 42513 649526
rect 42306 649468 42513 649470
rect 42306 649202 42366 649468
rect 42447 649465 42513 649468
rect 43215 648492 43281 648495
rect 42336 648490 43281 648492
rect 42336 648434 43220 648490
rect 43276 648434 43281 648490
rect 42336 648432 43281 648434
rect 43215 648429 43281 648432
rect 673978 648430 673984 648494
rect 674048 648492 674054 648494
rect 676474 648492 676480 648494
rect 674048 648432 676480 648492
rect 674048 648430 674054 648432
rect 676474 648430 676480 648432
rect 676544 648430 676550 648494
rect 674170 648282 674176 648346
rect 674240 648344 674246 648346
rect 675183 648344 675249 648347
rect 674240 648342 675249 648344
rect 674240 648286 675188 648342
rect 675244 648286 675249 648342
rect 674240 648284 675249 648286
rect 674240 648282 674246 648284
rect 675183 648281 675249 648284
rect 43407 647604 43473 647607
rect 42336 647602 43473 647604
rect 42336 647546 43412 647602
rect 43468 647546 43473 647602
rect 42336 647544 43473 647546
rect 43407 647541 43473 647544
rect 40578 646422 40638 646982
rect 42106 646654 42112 646718
rect 42176 646654 42182 646718
rect 40570 646358 40576 646422
rect 40640 646358 40646 646422
rect 42114 646124 42174 646654
rect 43311 646124 43377 646127
rect 42114 646122 43377 646124
rect 42114 646094 43316 646122
rect 42144 646066 43316 646094
rect 43372 646066 43377 646122
rect 42144 646064 43377 646066
rect 43311 646061 43377 646064
rect 654447 645976 654513 645979
rect 650208 645974 654513 645976
rect 650208 645918 654452 645974
rect 654508 645918 654513 645974
rect 650208 645916 654513 645918
rect 654447 645913 654513 645916
rect 42543 645532 42609 645535
rect 42306 645530 42609 645532
rect 42306 645474 42548 645530
rect 42604 645474 42609 645530
rect 42306 645472 42609 645474
rect 42306 645354 42366 645472
rect 42543 645469 42609 645472
rect 674362 645470 674368 645534
rect 674432 645532 674438 645534
rect 675471 645532 675537 645535
rect 674432 645530 675537 645532
rect 674432 645474 675476 645530
rect 675532 645474 675537 645530
rect 674432 645472 675537 645474
rect 674432 645470 674438 645472
rect 675471 645469 675537 645472
rect 675898 645026 675904 645090
rect 675968 645026 675974 645090
rect 675906 644940 675966 645026
rect 676858 644940 676864 644942
rect 675906 644880 676864 644940
rect 676858 644878 676864 644880
rect 676928 644878 676934 644942
rect 40002 643907 40062 644466
rect 40002 643902 40113 643907
rect 40002 643846 40052 643902
rect 40108 643846 40113 643902
rect 40002 643844 40113 643846
rect 40047 643841 40113 643844
rect 40770 643166 40830 643726
rect 40762 643102 40768 643166
rect 40832 643102 40838 643166
rect 41730 642427 41790 642838
rect 59535 642720 59601 642723
rect 59535 642718 64416 642720
rect 59535 642662 59540 642718
rect 59596 642662 64416 642718
rect 59535 642660 64416 642662
rect 59535 642657 59601 642660
rect 41679 642422 41790 642427
rect 41679 642366 41684 642422
rect 41740 642366 41790 642422
rect 41679 642364 41790 642366
rect 41679 642361 41745 642364
rect 41538 641687 41598 642172
rect 674895 641980 674961 641983
rect 675130 641980 675136 641982
rect 674895 641978 675136 641980
rect 674895 641922 674900 641978
rect 674956 641922 675136 641978
rect 674895 641920 675136 641922
rect 674895 641917 674961 641920
rect 675130 641918 675136 641920
rect 675200 641918 675206 641982
rect 41487 641682 41598 641687
rect 41487 641626 41492 641682
rect 41548 641626 41598 641682
rect 41487 641624 41598 641626
rect 41487 641621 41553 641624
rect 41730 640799 41790 641358
rect 41730 640794 41841 640799
rect 41730 640738 41780 640794
rect 41836 640738 41841 640794
rect 41730 640736 41841 640738
rect 41775 640733 41841 640736
rect 675706 640734 675712 640798
rect 675776 640796 675782 640798
rect 676666 640796 676672 640798
rect 675776 640736 676672 640796
rect 675776 640734 675782 640736
rect 676666 640734 676672 640736
rect 676736 640734 676742 640798
rect 40962 640058 41022 640544
rect 675087 640500 675153 640503
rect 676474 640500 676480 640502
rect 675087 640498 676480 640500
rect 675087 640442 675092 640498
rect 675148 640442 676480 640498
rect 675087 640440 676480 640442
rect 675087 640437 675153 640440
rect 676474 640438 676480 640440
rect 676544 640438 676550 640502
rect 675759 640352 675825 640355
rect 676474 640352 676480 640354
rect 675759 640350 676480 640352
rect 675759 640294 675764 640350
rect 675820 640294 676480 640350
rect 675759 640292 676480 640294
rect 675759 640289 675825 640292
rect 676474 640290 676480 640292
rect 676544 640290 676550 640354
rect 40954 639994 40960 640058
rect 41024 639994 41030 640058
rect 674746 639846 674752 639910
rect 674816 639846 674822 639910
rect 41922 639467 41982 639730
rect 41871 639462 41982 639467
rect 41871 639406 41876 639462
rect 41932 639406 41982 639462
rect 41871 639404 41982 639406
rect 674754 639464 674814 639846
rect 674938 639464 674944 639466
rect 674754 639404 674944 639464
rect 41871 639401 41937 639404
rect 674938 639402 674944 639404
rect 675008 639402 675014 639466
rect 42306 638428 42366 638916
rect 675130 638514 675136 638578
rect 675200 638576 675206 638578
rect 675375 638576 675441 638579
rect 675200 638574 675441 638576
rect 675200 638518 675380 638574
rect 675436 638518 675441 638574
rect 675200 638516 675441 638518
rect 675200 638514 675206 638516
rect 675375 638513 675441 638516
rect 42927 638428 42993 638431
rect 42306 638426 42993 638428
rect 42306 638370 42932 638426
rect 42988 638370 42993 638426
rect 42306 638368 42993 638370
rect 42927 638365 42993 638368
rect 43119 638132 43185 638135
rect 42336 638130 43185 638132
rect 42336 638074 43124 638130
rect 43180 638074 43185 638130
rect 42336 638072 43185 638074
rect 43119 638069 43185 638072
rect 674362 637774 674368 637838
rect 674432 637836 674438 637838
rect 675183 637836 675249 637839
rect 674432 637834 675249 637836
rect 674432 637778 675188 637834
rect 675244 637778 675249 637834
rect 674432 637776 675249 637778
rect 674432 637774 674438 637776
rect 675183 637773 675249 637776
rect 42114 636803 42174 637362
rect 42063 636798 42174 636803
rect 42063 636742 42068 636798
rect 42124 636742 42174 636798
rect 42063 636740 42174 636742
rect 42063 636737 42129 636740
rect 41922 636359 41982 636622
rect 41922 636354 42033 636359
rect 41922 636298 41972 636354
rect 42028 636298 42033 636354
rect 41922 636296 42033 636298
rect 41967 636293 42033 636296
rect 42639 635912 42705 635915
rect 42874 635912 42880 635914
rect 42639 635910 42880 635912
rect 42639 635854 42644 635910
rect 42700 635854 42880 635910
rect 42639 635852 42880 635854
rect 42639 635849 42705 635852
rect 42874 635850 42880 635852
rect 42944 635850 42950 635914
rect 41538 635174 41598 635734
rect 41530 635110 41536 635174
rect 41600 635110 41606 635174
rect 676719 635024 676785 635027
rect 676858 635024 676864 635026
rect 676719 635022 676864 635024
rect 42306 634432 42366 634994
rect 676719 634966 676724 635022
rect 676780 634966 676864 635022
rect 676719 634964 676864 634966
rect 676719 634961 676785 634964
rect 676858 634962 676864 634964
rect 676928 634962 676934 635026
rect 42490 634432 42496 634434
rect 42306 634372 42496 634432
rect 42490 634370 42496 634372
rect 42560 634370 42566 634434
rect 655215 634284 655281 634287
rect 650208 634282 655281 634284
rect 650208 634226 655220 634282
rect 655276 634226 655281 634282
rect 650208 634224 655281 634226
rect 655215 634221 655281 634224
rect 42114 633547 42174 634106
rect 42114 633542 42225 633547
rect 42114 633486 42164 633542
rect 42220 633486 42225 633542
rect 42114 633484 42225 633486
rect 42159 633481 42225 633484
rect 676047 633250 676113 633251
rect 676047 633246 676096 633250
rect 676160 633248 676166 633250
rect 676047 633190 676052 633246
rect 676047 633186 676096 633190
rect 676160 633188 676204 633248
rect 676160 633186 676166 633188
rect 676047 633185 676113 633186
rect 42306 632511 42366 632626
rect 42255 632506 42366 632511
rect 42255 632450 42260 632506
rect 42316 632450 42366 632506
rect 42255 632448 42366 632450
rect 674703 632508 674769 632511
rect 674703 632506 674814 632508
rect 674703 632450 674708 632506
rect 674764 632450 674814 632506
rect 42255 632445 42321 632448
rect 674703 632445 674814 632450
rect 674754 632330 674814 632445
rect 674703 631768 674769 631771
rect 674703 631766 674814 631768
rect 674703 631710 674708 631766
rect 674764 631710 674814 631766
rect 674703 631705 674814 631710
rect 674754 631442 674814 631705
rect 674127 630732 674193 630735
rect 674127 630730 674784 630732
rect 674127 630674 674132 630730
rect 674188 630674 674784 630730
rect 674127 630672 674784 630674
rect 674127 630669 674193 630672
rect 674170 630374 674176 630438
rect 674240 630436 674246 630438
rect 676858 630436 676864 630438
rect 674240 630376 676864 630436
rect 674240 630374 674246 630376
rect 676858 630374 676864 630376
rect 676928 630374 676934 630438
rect 675183 630140 675249 630143
rect 676719 630142 676785 630143
rect 676090 630140 676096 630142
rect 675183 630138 676096 630140
rect 675183 630082 675188 630138
rect 675244 630082 676096 630138
rect 675183 630080 676096 630082
rect 675183 630077 675249 630080
rect 676090 630078 676096 630080
rect 676160 630078 676166 630142
rect 676666 630078 676672 630142
rect 676736 630140 676785 630142
rect 676736 630138 676828 630140
rect 676780 630082 676828 630138
rect 676736 630080 676828 630082
rect 676736 630078 676785 630080
rect 676719 630077 676785 630078
rect 673839 629844 673905 629847
rect 673839 629842 674784 629844
rect 673839 629786 673844 629842
rect 673900 629786 674784 629842
rect 673839 629784 674784 629786
rect 673839 629781 673905 629784
rect 673839 629104 673905 629107
rect 673839 629102 674784 629104
rect 673839 629046 673844 629102
rect 673900 629046 674784 629102
rect 673839 629044 674784 629046
rect 673839 629041 673905 629044
rect 670959 628364 671025 628367
rect 670959 628362 674784 628364
rect 670959 628306 670964 628362
rect 671020 628306 674784 628362
rect 670959 628304 674784 628306
rect 670959 628301 671025 628304
rect 58383 628216 58449 628219
rect 58383 628214 64416 628216
rect 58383 628158 58388 628214
rect 58444 628158 64416 628214
rect 58383 628156 64416 628158
rect 58383 628153 58449 628156
rect 41199 627772 41265 627775
rect 41338 627772 41344 627774
rect 41199 627770 41344 627772
rect 41199 627714 41204 627770
rect 41260 627714 41344 627770
rect 41199 627712 41344 627714
rect 41199 627709 41265 627712
rect 41338 627710 41344 627712
rect 41408 627710 41414 627774
rect 41967 627624 42033 627627
rect 42298 627624 42304 627626
rect 41967 627622 42304 627624
rect 41967 627566 41972 627622
rect 42028 627566 42304 627622
rect 41967 627564 42304 627566
rect 41967 627561 42033 627564
rect 42298 627562 42304 627564
rect 42368 627562 42374 627626
rect 41871 627476 41937 627479
rect 42106 627476 42112 627478
rect 41871 627474 42112 627476
rect 41871 627418 41876 627474
rect 41932 627418 42112 627474
rect 41871 627416 42112 627418
rect 41871 627413 41937 627416
rect 42106 627414 42112 627416
rect 42176 627414 42182 627478
rect 670863 627476 670929 627479
rect 674754 627476 674814 627520
rect 670863 627474 674814 627476
rect 670863 627418 670868 627474
rect 670924 627418 674814 627474
rect 670863 627416 674814 627418
rect 670863 627413 670929 627416
rect 674746 627266 674752 627330
rect 674816 627266 674822 627330
rect 674754 626706 674814 627266
rect 674511 626144 674577 626147
rect 674511 626142 674814 626144
rect 674511 626086 674516 626142
rect 674572 626086 674814 626142
rect 674511 626084 674814 626086
rect 674511 626081 674577 626084
rect 674754 625892 674814 626084
rect 674895 625700 674961 625703
rect 674895 625698 675006 625700
rect 674895 625642 674900 625698
rect 674956 625642 675006 625698
rect 674895 625637 675006 625642
rect 41338 625194 41344 625258
rect 41408 625256 41414 625258
rect 42159 625256 42225 625259
rect 41408 625254 42225 625256
rect 41408 625198 42164 625254
rect 42220 625198 42225 625254
rect 41408 625196 42225 625198
rect 41408 625194 41414 625196
rect 42159 625193 42225 625196
rect 674946 625078 675006 625637
rect 674031 624962 674097 624963
rect 673978 624960 673984 624962
rect 673940 624900 673984 624960
rect 674048 624958 674097 624962
rect 674092 624902 674097 624958
rect 673978 624898 673984 624900
rect 674048 624898 674097 624902
rect 674031 624897 674097 624898
rect 676047 624812 676113 624815
rect 676047 624810 676158 624812
rect 676047 624754 676052 624810
rect 676108 624754 676158 624810
rect 676047 624749 676158 624754
rect 42106 624454 42112 624518
rect 42176 624516 42182 624518
rect 42447 624516 42513 624519
rect 42176 624514 42513 624516
rect 42176 624458 42452 624514
rect 42508 624458 42513 624514
rect 42176 624456 42513 624458
rect 42176 624454 42182 624456
rect 42447 624453 42513 624456
rect 41530 624306 41536 624370
rect 41600 624368 41606 624370
rect 42106 624368 42112 624370
rect 41600 624308 42112 624368
rect 41600 624306 41606 624308
rect 42106 624306 42112 624308
rect 42176 624306 42182 624370
rect 676098 624264 676158 624749
rect 674319 623628 674385 623631
rect 674319 623626 674784 623628
rect 674319 623570 674324 623626
rect 674380 623570 674784 623626
rect 674319 623568 674784 623570
rect 674319 623565 674385 623568
rect 674415 622740 674481 622743
rect 674415 622738 674784 622740
rect 674415 622682 674420 622738
rect 674476 622682 674784 622738
rect 674415 622680 674784 622682
rect 674415 622677 674481 622680
rect 654447 622444 654513 622447
rect 650208 622442 654513 622444
rect 650208 622386 654452 622442
rect 654508 622386 654513 622442
rect 650208 622384 654513 622386
rect 654447 622381 654513 622384
rect 42159 622148 42225 622151
rect 42490 622148 42496 622150
rect 42159 622146 42496 622148
rect 42159 622090 42164 622146
rect 42220 622090 42496 622146
rect 42159 622088 42496 622090
rect 42159 622085 42225 622088
rect 42490 622086 42496 622088
rect 42560 622086 42566 622150
rect 675087 622148 675153 622151
rect 675087 622146 675774 622148
rect 675087 622090 675092 622146
rect 675148 622090 675774 622146
rect 675087 622088 675774 622090
rect 675087 622085 675153 622088
rect 675714 621970 675774 622088
rect 674554 621642 674560 621706
rect 674624 621704 674630 621706
rect 674624 621644 674814 621704
rect 674624 621642 674630 621644
rect 674754 621082 674814 621644
rect 42063 620966 42129 620967
rect 42063 620964 42112 620966
rect 42020 620962 42112 620964
rect 42020 620906 42068 620962
rect 42020 620904 42112 620906
rect 42063 620902 42112 620904
rect 42176 620902 42182 620966
rect 676666 620902 676672 620966
rect 676736 620902 676742 620966
rect 42063 620901 42129 620902
rect 42298 620754 42304 620818
rect 42368 620816 42374 620818
rect 42447 620816 42513 620819
rect 42368 620814 42513 620816
rect 42368 620758 42452 620814
rect 42508 620758 42513 620814
rect 42368 620756 42513 620758
rect 42368 620754 42374 620756
rect 42447 620753 42513 620756
rect 676674 620342 676734 620902
rect 674223 619484 674289 619487
rect 674223 619482 674784 619484
rect 674223 619426 674228 619482
rect 674284 619426 674784 619482
rect 674223 619424 674784 619426
rect 674223 619421 674289 619424
rect 41775 619190 41841 619191
rect 41722 619126 41728 619190
rect 41792 619188 41841 619190
rect 41792 619186 41884 619188
rect 41836 619130 41884 619186
rect 41792 619128 41884 619130
rect 41792 619126 41841 619128
rect 41775 619125 41841 619126
rect 674170 618830 674176 618894
rect 674240 618892 674246 618894
rect 674240 618832 674784 618892
rect 674240 618830 674246 618832
rect 41871 618302 41937 618303
rect 42831 618302 42897 618303
rect 41871 618300 41920 618302
rect 41828 618298 41920 618300
rect 41828 618242 41876 618298
rect 41828 618240 41920 618242
rect 41871 618238 41920 618240
rect 41984 618238 41990 618302
rect 42831 618300 42880 618302
rect 42788 618298 42880 618300
rect 42788 618242 42836 618298
rect 42788 618240 42880 618242
rect 42831 618238 42880 618240
rect 42944 618238 42950 618302
rect 41871 618237 41937 618238
rect 42831 618237 42897 618238
rect 40762 618090 40768 618154
rect 40832 618152 40838 618154
rect 42735 618152 42801 618155
rect 40832 618150 42801 618152
rect 40832 618094 42740 618150
rect 42796 618094 42801 618150
rect 40832 618092 42801 618094
rect 40832 618090 40838 618092
rect 42735 618089 42801 618092
rect 673839 618004 673905 618007
rect 673839 618002 674784 618004
rect 673839 617946 673844 618002
rect 673900 617946 674784 618002
rect 673839 617944 674784 617946
rect 673839 617941 673905 617944
rect 677050 617794 677056 617858
rect 677120 617794 677126 617858
rect 40954 617646 40960 617710
rect 41024 617708 41030 617710
rect 42447 617708 42513 617711
rect 41024 617706 42513 617708
rect 41024 617650 42452 617706
rect 42508 617650 42513 617706
rect 41024 617648 42513 617650
rect 41024 617646 41030 617648
rect 42447 617645 42513 617648
rect 677058 617234 677118 617794
rect 673839 616376 673905 616379
rect 673839 616374 674784 616376
rect 673839 616318 673844 616374
rect 673900 616318 674784 616374
rect 673839 616316 674784 616318
rect 673839 616313 673905 616316
rect 679746 615047 679806 615606
rect 679695 615042 679806 615047
rect 679695 614986 679700 615042
rect 679756 614986 679806 615042
rect 679695 614984 679806 614986
rect 679695 614981 679761 614984
rect 679695 614452 679761 614455
rect 679695 614450 679806 614452
rect 679695 614394 679700 614450
rect 679756 614394 679806 614450
rect 679695 614389 679806 614394
rect 679746 614052 679806 614389
rect 58383 613860 58449 613863
rect 58383 613858 64416 613860
rect 58383 613802 58388 613858
rect 58444 613802 64416 613858
rect 58383 613800 64416 613802
rect 58383 613797 58449 613800
rect 654447 610752 654513 610755
rect 650208 610750 654513 610752
rect 650208 610694 654452 610750
rect 654508 610694 654513 610750
rect 650208 610692 654513 610694
rect 654447 610689 654513 610692
rect 674362 607730 674368 607794
rect 674432 607792 674438 607794
rect 675087 607792 675153 607795
rect 674432 607790 675153 607792
rect 674432 607734 675092 607790
rect 675148 607734 675153 607790
rect 674432 607732 675153 607734
rect 674432 607730 674438 607732
rect 675087 607729 675153 607732
rect 42735 607718 42801 607721
rect 42336 607716 42801 607718
rect 42336 607660 42740 607716
rect 42796 607660 42801 607716
rect 42336 607658 42801 607660
rect 42735 607655 42801 607658
rect 674554 607434 674560 607498
rect 674624 607496 674630 607498
rect 675087 607496 675153 607499
rect 674624 607494 675153 607496
rect 674624 607438 675092 607494
rect 675148 607438 675153 607494
rect 674624 607436 675153 607438
rect 674624 607434 674630 607436
rect 675087 607433 675153 607436
rect 42735 606904 42801 606907
rect 42336 606902 42801 606904
rect 42336 606846 42740 606902
rect 42796 606846 42801 606902
rect 42336 606844 42801 606846
rect 42735 606841 42801 606844
rect 675663 606462 675729 606463
rect 675663 606458 675712 606462
rect 675776 606460 675782 606462
rect 675663 606402 675668 606458
rect 675663 606398 675712 606402
rect 675776 606400 675820 606460
rect 675776 606398 675782 606400
rect 675663 606397 675729 606398
rect 42447 606312 42513 606315
rect 42306 606310 42513 606312
rect 42306 606254 42452 606310
rect 42508 606254 42513 606310
rect 42306 606252 42513 606254
rect 42306 606060 42366 606252
rect 42447 606249 42513 606252
rect 43503 605276 43569 605279
rect 42336 605274 43569 605276
rect 42336 605218 43508 605274
rect 43564 605218 43569 605274
rect 42336 605216 43569 605218
rect 43503 605213 43569 605216
rect 673978 604918 673984 604982
rect 674048 604980 674054 604982
rect 675087 604980 675153 604983
rect 674048 604978 675153 604980
rect 674048 604922 675092 604978
rect 675148 604922 675153 604978
rect 674048 604920 675153 604922
rect 674048 604918 674054 604920
rect 675087 604917 675153 604920
rect 674031 604832 674097 604835
rect 674170 604832 674176 604834
rect 674031 604830 674176 604832
rect 674031 604774 674036 604830
rect 674092 604774 674176 604830
rect 674031 604772 674176 604774
rect 674031 604769 674097 604772
rect 674170 604770 674176 604772
rect 674240 604770 674246 604834
rect 43215 604684 43281 604687
rect 42306 604682 43281 604684
rect 42306 604626 43220 604682
rect 43276 604626 43281 604682
rect 42306 604624 43281 604626
rect 42306 604432 42366 604624
rect 43215 604621 43281 604624
rect 40570 603882 40576 603946
rect 40640 603882 40646 603946
rect 40578 603796 40638 603882
rect 40578 603766 42144 603796
rect 40608 603736 42174 603766
rect 42114 603206 42174 603736
rect 42106 603142 42112 603206
rect 42176 603142 42182 603206
rect 43311 602908 43377 602911
rect 42336 602906 43377 602908
rect 42336 602850 43316 602906
rect 43372 602850 43377 602906
rect 42336 602848 43377 602850
rect 43311 602845 43377 602848
rect 42927 602168 42993 602171
rect 42336 602166 42993 602168
rect 42336 602110 42932 602166
rect 42988 602110 42993 602166
rect 42336 602108 42993 602110
rect 42927 602105 42993 602108
rect 40002 600691 40062 601250
rect 40002 600686 40113 600691
rect 40002 600630 40052 600686
rect 40108 600630 40113 600686
rect 40002 600628 40113 600630
rect 40047 600625 40113 600628
rect 40578 599950 40638 600510
rect 675759 600244 675825 600247
rect 675898 600244 675904 600246
rect 675759 600242 675904 600244
rect 675759 600186 675764 600242
rect 675820 600186 675904 600242
rect 675759 600184 675904 600186
rect 675759 600181 675825 600184
rect 675898 600182 675904 600184
rect 675968 600182 675974 600246
rect 40570 599886 40576 599950
rect 40640 599886 40646 599950
rect 43023 599652 43089 599655
rect 42336 599650 43089 599652
rect 42336 599594 43028 599650
rect 43084 599594 43089 599650
rect 42336 599592 43089 599594
rect 43023 599589 43089 599592
rect 59535 599504 59601 599507
rect 59535 599502 64416 599504
rect 59535 599446 59540 599502
rect 59596 599446 64416 599502
rect 59535 599444 64416 599446
rect 59535 599441 59601 599444
rect 654447 599356 654513 599359
rect 649986 599354 654513 599356
rect 649986 599298 654452 599354
rect 654508 599298 654513 599354
rect 649986 599296 654513 599298
rect 649986 599178 650046 599296
rect 654447 599293 654513 599296
rect 674938 599146 674944 599210
rect 675008 599208 675014 599210
rect 676090 599208 676096 599210
rect 675008 599148 676096 599208
rect 675008 599146 675014 599148
rect 676090 599146 676096 599148
rect 676160 599146 676166 599210
rect 41922 598471 41982 599030
rect 41871 598466 41982 598471
rect 41871 598410 41876 598466
rect 41932 598410 41982 598466
rect 41871 598408 41982 598410
rect 41871 598405 41937 598408
rect 41730 597583 41790 598142
rect 41730 597578 41841 597583
rect 41730 597522 41780 597578
rect 41836 597522 41841 597578
rect 41730 597520 41841 597522
rect 41775 597517 41841 597520
rect 40962 596842 41022 597402
rect 40954 596778 40960 596842
rect 41024 596778 41030 596842
rect 41922 596251 41982 596514
rect 41922 596246 42033 596251
rect 41922 596190 41972 596246
rect 42028 596190 42033 596246
rect 41922 596188 42033 596190
rect 41967 596185 42033 596188
rect 42114 595215 42174 595774
rect 675759 595360 675825 595363
rect 676666 595360 676672 595362
rect 675759 595358 676672 595360
rect 675759 595302 675764 595358
rect 675820 595302 676672 595358
rect 675759 595300 676672 595302
rect 675759 595297 675825 595300
rect 676666 595298 676672 595300
rect 676736 595298 676742 595362
rect 42063 595210 42174 595215
rect 42063 595154 42068 595210
rect 42124 595154 42174 595210
rect 42063 595152 42174 595154
rect 42063 595149 42129 595152
rect 42831 594916 42897 594919
rect 42336 594914 42897 594916
rect 42336 594858 42836 594914
rect 42892 594858 42897 594914
rect 42336 594856 42897 594858
rect 42831 594853 42897 594856
rect 42114 593735 42174 594220
rect 42114 593730 42225 593735
rect 42114 593674 42164 593730
rect 42220 593674 42225 593730
rect 42114 593672 42225 593674
rect 42159 593669 42225 593672
rect 43119 593436 43185 593439
rect 42336 593434 43185 593436
rect 42336 593378 43124 593434
rect 43180 593378 43185 593434
rect 42336 593376 43185 593378
rect 43119 593373 43185 593376
rect 675759 593436 675825 593439
rect 676090 593436 676096 593438
rect 675759 593434 676096 593436
rect 675759 593378 675764 593434
rect 675820 593378 676096 593434
rect 675759 593376 676096 593378
rect 675759 593373 675825 593376
rect 676090 593374 676096 593376
rect 676160 593374 676166 593438
rect 42306 592400 42366 592592
rect 42447 592400 42513 592403
rect 42306 592398 42513 592400
rect 42306 592342 42452 592398
rect 42508 592342 42513 592398
rect 42306 592340 42513 592342
rect 42447 592337 42513 592340
rect 42543 591956 42609 591959
rect 42306 591954 42609 591956
rect 42306 591898 42548 591954
rect 42604 591898 42609 591954
rect 42306 591896 42609 591898
rect 42306 591778 42366 591896
rect 42543 591893 42609 591896
rect 42306 590772 42366 590964
rect 42543 590772 42609 590775
rect 42306 590770 42609 590772
rect 42306 590714 42548 590770
rect 42604 590714 42609 590770
rect 42306 590712 42609 590714
rect 42543 590709 42609 590712
rect 42306 589292 42366 589410
rect 42543 589292 42609 589295
rect 42306 589290 42609 589292
rect 42306 589234 42548 589290
rect 42604 589234 42609 589290
rect 42306 589232 42609 589234
rect 42543 589229 42609 589232
rect 654447 587220 654513 587223
rect 650208 587218 654513 587220
rect 650208 587162 654452 587218
rect 654508 587162 654513 587218
rect 650208 587160 654513 587162
rect 654447 587157 654513 587160
rect 42927 586628 42993 586631
rect 43066 586628 43072 586630
rect 42927 586626 43072 586628
rect 42927 586570 42932 586626
rect 42988 586570 43072 586626
rect 42927 586568 43072 586570
rect 42927 586565 42993 586568
rect 43066 586566 43072 586568
rect 43136 586566 43142 586630
rect 674754 586483 674814 587042
rect 674703 586478 674814 586483
rect 674703 586422 674708 586478
rect 674764 586422 674814 586478
rect 674703 586420 674814 586422
rect 674703 586417 674769 586420
rect 674415 586332 674481 586335
rect 674415 586330 674784 586332
rect 674415 586274 674420 586330
rect 674476 586274 674784 586330
rect 674415 586272 674784 586274
rect 674415 586269 674481 586272
rect 674415 585444 674481 585447
rect 674415 585442 674784 585444
rect 674415 585386 674420 585442
rect 674476 585386 674784 585442
rect 674415 585384 674784 585386
rect 674415 585381 674481 585384
rect 59535 585296 59601 585299
rect 59535 585294 64416 585296
rect 59535 585238 59540 585294
rect 59596 585238 64416 585294
rect 59535 585236 64416 585238
rect 59535 585233 59601 585236
rect 42543 585002 42609 585003
rect 42490 585000 42496 585002
rect 42452 584940 42496 585000
rect 42560 584998 42609 585002
rect 42604 584942 42609 584998
rect 42490 584938 42496 584940
rect 42560 584938 42609 584942
rect 42543 584937 42609 584938
rect 674607 584852 674673 584855
rect 674607 584850 674814 584852
rect 674607 584794 674612 584850
rect 674668 584794 674814 584850
rect 674607 584792 674814 584794
rect 674607 584789 674673 584792
rect 674754 584674 674814 584792
rect 41338 584494 41344 584558
rect 41408 584556 41414 584558
rect 42063 584556 42129 584559
rect 41408 584554 42129 584556
rect 41408 584498 42068 584554
rect 42124 584498 42129 584554
rect 41408 584496 42129 584498
rect 41408 584494 41414 584496
rect 42063 584493 42129 584496
rect 42447 584554 42513 584559
rect 674223 584558 674289 584559
rect 673978 584556 673984 584558
rect 42447 584498 42452 584554
rect 42508 584498 42513 584554
rect 42447 584493 42513 584498
rect 673794 584496 673984 584556
rect 41530 584346 41536 584410
rect 41600 584408 41606 584410
rect 41871 584408 41937 584411
rect 41600 584406 41937 584408
rect 41600 584350 41876 584406
rect 41932 584350 41937 584406
rect 41600 584348 41937 584350
rect 41600 584346 41606 584348
rect 41871 584345 41937 584348
rect 42450 584263 42510 584493
rect 42927 584410 42993 584411
rect 42874 584408 42880 584410
rect 42836 584348 42880 584408
rect 42944 584406 42993 584410
rect 42988 584350 42993 584406
rect 42874 584346 42880 584348
rect 42944 584346 42993 584350
rect 42927 584345 42993 584346
rect 41967 584260 42033 584263
rect 42298 584260 42304 584262
rect 41967 584258 42304 584260
rect 41967 584202 41972 584258
rect 42028 584202 42304 584258
rect 41967 584200 42304 584202
rect 41967 584197 42033 584200
rect 42298 584198 42304 584200
rect 42368 584198 42374 584262
rect 42447 584258 42513 584263
rect 42447 584202 42452 584258
rect 42508 584202 42513 584258
rect 42447 584197 42513 584202
rect 673794 584112 673854 584496
rect 673978 584494 673984 584496
rect 674048 584494 674054 584558
rect 674170 584494 674176 584558
rect 674240 584556 674289 584558
rect 674240 584554 674332 584556
rect 674284 584498 674332 584554
rect 674240 584496 674332 584498
rect 674240 584494 674289 584496
rect 674223 584493 674289 584494
rect 673978 584112 673984 584114
rect 673794 584052 673984 584112
rect 673978 584050 673984 584052
rect 674048 584050 674054 584114
rect 674754 583671 674814 583786
rect 674703 583666 674814 583671
rect 674703 583610 674708 583666
rect 674764 583610 674814 583666
rect 674703 583608 674814 583610
rect 674703 583605 674769 583608
rect 674703 583372 674769 583375
rect 674703 583370 674814 583372
rect 674703 583314 674708 583370
rect 674764 583314 674814 583370
rect 674703 583309 674814 583314
rect 674754 583194 674814 583309
rect 679695 582928 679761 582931
rect 679695 582926 679806 582928
rect 679695 582870 679700 582926
rect 679756 582870 679806 582926
rect 679695 582865 679806 582870
rect 679746 582336 679806 582865
rect 676896 582306 679806 582336
rect 676866 582276 679776 582306
rect 676866 581894 676926 582276
rect 676858 581830 676864 581894
rect 676928 581830 676934 581894
rect 675322 581682 675328 581746
rect 675392 581682 675398 581746
rect 675330 581566 675390 581682
rect 42298 581238 42304 581302
rect 42368 581300 42374 581302
rect 42831 581300 42897 581303
rect 42368 581298 42897 581300
rect 42368 581242 42836 581298
rect 42892 581242 42897 581298
rect 42368 581240 42897 581242
rect 42368 581238 42374 581240
rect 42831 581237 42897 581240
rect 676474 581238 676480 581302
rect 676544 581238 676550 581302
rect 676482 580678 676542 581238
rect 675514 580350 675520 580414
rect 675584 580350 675590 580414
rect 675522 579864 675582 580350
rect 676282 579610 676288 579674
rect 676352 579610 676358 579674
rect 676290 579050 676350 579610
rect 42927 578342 42993 578343
rect 42874 578278 42880 578342
rect 42944 578340 42993 578342
rect 42944 578338 43036 578340
rect 42988 578282 43036 578338
rect 42944 578280 43036 578282
rect 42944 578278 42993 578280
rect 42927 578277 42993 578278
rect 674946 578194 675006 578384
rect 674938 578130 674944 578194
rect 675008 578130 675014 578194
rect 675130 578130 675136 578194
rect 675200 578130 675206 578194
rect 43023 577602 43089 577603
rect 43023 577600 43072 577602
rect 42980 577598 43072 577600
rect 42980 577542 43028 577598
rect 42980 577540 43072 577542
rect 43023 577538 43072 577540
rect 43136 577538 43142 577602
rect 675138 577570 675198 578130
rect 43023 577537 43089 577538
rect 674746 577242 674752 577306
rect 674816 577242 674822 577306
rect 41530 577094 41536 577158
rect 41600 577156 41606 577158
rect 41775 577156 41841 577159
rect 41600 577154 41841 577156
rect 41600 577098 41780 577154
rect 41836 577098 41841 577154
rect 41600 577096 41841 577098
rect 41600 577094 41606 577096
rect 41775 577093 41841 577096
rect 42447 577010 42513 577011
rect 42447 577008 42496 577010
rect 42404 577006 42496 577008
rect 42404 576950 42452 577006
rect 42404 576948 42496 576950
rect 42447 576946 42496 576948
rect 42560 576946 42566 577010
rect 42447 576945 42513 576946
rect 674754 576756 674814 577242
rect 674223 575972 674289 575975
rect 674223 575970 674784 575972
rect 674223 575914 674228 575970
rect 674284 575914 674784 575970
rect 674223 575912 674784 575914
rect 674223 575909 674289 575912
rect 654447 575528 654513 575531
rect 650208 575526 654513 575528
rect 650208 575470 654452 575526
rect 654508 575470 654513 575526
rect 650208 575468 654513 575470
rect 654447 575465 654513 575468
rect 674703 575380 674769 575383
rect 674703 575378 674814 575380
rect 674703 575322 674708 575378
rect 674764 575322 674814 575378
rect 674703 575317 674814 575322
rect 674754 575128 674814 575317
rect 41871 575086 41937 575087
rect 41871 575084 41920 575086
rect 41828 575082 41920 575084
rect 41828 575026 41876 575082
rect 41828 575024 41920 575026
rect 41871 575022 41920 575024
rect 41984 575022 41990 575086
rect 41871 575021 41937 575022
rect 41775 574938 41841 574939
rect 41722 574874 41728 574938
rect 41792 574936 41841 574938
rect 41792 574934 41884 574936
rect 41836 574878 41884 574934
rect 41792 574876 41884 574878
rect 41792 574874 41841 574876
rect 41775 574873 41841 574874
rect 674703 574492 674769 574495
rect 674703 574490 674814 574492
rect 674703 574434 674708 574490
rect 674764 574434 674814 574490
rect 674703 574429 674814 574434
rect 674754 574314 674814 574429
rect 40954 573986 40960 574050
rect 41024 574048 41030 574050
rect 42255 574048 42321 574051
rect 41024 574046 42321 574048
rect 41024 573990 42260 574046
rect 42316 573990 42321 574046
rect 41024 573988 42321 573990
rect 41024 573986 41030 573988
rect 42255 573985 42321 573988
rect 41338 573838 41344 573902
rect 41408 573900 41414 573902
rect 41775 573900 41841 573903
rect 41408 573898 41841 573900
rect 41408 573842 41780 573898
rect 41836 573842 41841 573898
rect 41408 573840 41841 573842
rect 41408 573838 41414 573840
rect 41775 573837 41841 573840
rect 674415 573604 674481 573607
rect 674415 573602 674784 573604
rect 674415 573546 674420 573602
rect 674476 573546 674784 573602
rect 674415 573544 674784 573546
rect 674415 573541 674481 573544
rect 40570 573246 40576 573310
rect 40640 573308 40646 573310
rect 42831 573308 42897 573311
rect 40640 573306 42897 573308
rect 40640 573250 42836 573306
rect 42892 573250 42897 573306
rect 40640 573248 42897 573250
rect 40640 573246 40646 573248
rect 42831 573245 42897 573248
rect 674703 573012 674769 573015
rect 674703 573010 674814 573012
rect 674703 572954 674708 573010
rect 674764 572954 674814 573010
rect 674703 572949 674814 572954
rect 674754 572834 674814 572949
rect 674415 571976 674481 571979
rect 674415 571974 674784 571976
rect 674415 571918 674420 571974
rect 674476 571918 674784 571974
rect 674415 571916 674784 571918
rect 674415 571913 674481 571916
rect 674703 571384 674769 571387
rect 674703 571382 674814 571384
rect 674703 571326 674708 571382
rect 674764 571326 674814 571382
rect 674703 571321 674814 571326
rect 674754 571206 674814 571321
rect 59535 570792 59601 570795
rect 59535 570790 64416 570792
rect 59535 570734 59540 570790
rect 59596 570734 64416 570790
rect 59535 570732 64416 570734
rect 59535 570729 59601 570732
rect 679746 569759 679806 570318
rect 679746 569754 679857 569759
rect 679746 569698 679796 569754
rect 679852 569698 679857 569754
rect 679746 569696 679857 569698
rect 679791 569693 679857 569696
rect 679791 569164 679857 569167
rect 679746 569162 679857 569164
rect 679746 569106 679796 569162
rect 679852 569106 679857 569162
rect 679746 569101 679857 569106
rect 679746 568838 679806 569101
rect 675514 567326 675520 567390
rect 675584 567388 675590 567390
rect 679983 567388 680049 567391
rect 675584 567386 680049 567388
rect 675584 567330 679988 567386
rect 680044 567330 680049 567386
rect 675584 567328 680049 567330
rect 675584 567326 675590 567328
rect 679983 567325 680049 567328
rect 34479 564724 34545 564727
rect 34434 564722 34545 564724
rect 34434 564666 34484 564722
rect 34540 564666 34545 564722
rect 34434 564661 34545 564666
rect 34434 564472 34494 564661
rect 43311 564576 43377 564579
rect 43599 564576 43665 564579
rect 43311 564574 43665 564576
rect 43311 564518 43316 564574
rect 43372 564518 43604 564574
rect 43660 564518 43665 564574
rect 43311 564516 43665 564518
rect 43311 564513 43377 564516
rect 43599 564513 43665 564516
rect 654447 563836 654513 563839
rect 650208 563834 654513 563836
rect 650208 563778 654452 563834
rect 654508 563778 654513 563834
rect 650208 563776 654513 563778
rect 654447 563773 654513 563776
rect 42306 563540 42366 563658
rect 42447 563540 42513 563543
rect 42306 563538 42513 563540
rect 42306 563482 42452 563538
rect 42508 563482 42513 563538
rect 42306 563480 42513 563482
rect 42447 563477 42513 563480
rect 42351 563096 42417 563099
rect 42306 563094 42417 563096
rect 42306 563038 42356 563094
rect 42412 563038 42417 563094
rect 42306 563033 42417 563038
rect 42306 562844 42366 563033
rect 674938 562886 674944 562950
rect 675008 562948 675014 562950
rect 675087 562948 675153 562951
rect 675008 562946 675153 562948
rect 675008 562890 675092 562946
rect 675148 562890 675153 562946
rect 675008 562888 675153 562890
rect 675008 562886 675014 562888
rect 675087 562885 675153 562888
rect 43215 562060 43281 562063
rect 42336 562058 43281 562060
rect 42336 562002 43220 562058
rect 43276 562002 43281 562058
rect 42336 562000 43281 562002
rect 43215 561997 43281 562000
rect 674170 561702 674176 561766
rect 674240 561764 674246 561766
rect 675087 561764 675153 561767
rect 674240 561762 675153 561764
rect 674240 561706 675092 561762
rect 675148 561706 675153 561762
rect 674240 561704 675153 561706
rect 674240 561702 674246 561704
rect 675087 561701 675153 561704
rect 43503 561616 43569 561619
rect 42306 561614 43569 561616
rect 42306 561558 43508 561614
rect 43564 561558 43569 561614
rect 42306 561556 43569 561558
rect 42306 561216 42366 561556
rect 43503 561553 43569 561556
rect 675130 561554 675136 561618
rect 675200 561616 675206 561618
rect 675279 561616 675345 561619
rect 675200 561614 675345 561616
rect 675200 561558 675284 561614
rect 675340 561558 675345 561614
rect 675200 561556 675345 561558
rect 675200 561554 675206 561556
rect 675279 561553 675345 561556
rect 42106 560962 42112 561026
rect 42176 560962 42182 561026
rect 42114 560580 42174 560962
rect 43791 560580 43857 560583
rect 42114 560578 43857 560580
rect 42114 560550 43796 560578
rect 42144 560522 43796 560550
rect 43852 560522 43857 560578
rect 42144 560520 43857 560522
rect 43791 560517 43857 560520
rect 43599 559840 43665 559843
rect 42306 559838 43665 559840
rect 42306 559782 43604 559838
rect 43660 559782 43665 559838
rect 42306 559780 43665 559782
rect 42306 559736 42366 559780
rect 43599 559777 43665 559780
rect 41730 558656 41790 558922
rect 674746 558890 674752 558954
rect 674816 558952 674822 558954
rect 675471 558952 675537 558955
rect 674816 558950 675537 558952
rect 674816 558894 675476 558950
rect 675532 558894 675537 558950
rect 674816 558892 675537 558894
rect 674816 558890 674822 558892
rect 675471 558889 675537 558892
rect 41967 558656 42033 558659
rect 41730 558654 42033 558656
rect 41730 558598 41972 558654
rect 42028 558598 42033 558654
rect 41730 558596 42033 558598
rect 41967 558593 42033 558596
rect 40194 557475 40254 558034
rect 675759 557768 675825 557771
rect 676282 557768 676288 557770
rect 675759 557766 676288 557768
rect 675759 557710 675764 557766
rect 675820 557710 676288 557766
rect 675759 557708 676288 557710
rect 675759 557705 675825 557708
rect 676282 557706 676288 557708
rect 676352 557706 676358 557770
rect 40143 557470 40254 557475
rect 40143 557414 40148 557470
rect 40204 557414 40254 557470
rect 40143 557412 40254 557414
rect 40143 557409 40209 557412
rect 40578 556734 40638 557294
rect 40570 556670 40576 556734
rect 40640 556670 40646 556734
rect 59535 556584 59601 556587
rect 59535 556582 64416 556584
rect 59535 556526 59540 556582
rect 59596 556526 64416 556582
rect 59535 556524 64416 556526
rect 59535 556521 59601 556524
rect 41730 555995 41790 556406
rect 41679 555990 41790 555995
rect 41679 555934 41684 555990
rect 41740 555934 41790 555990
rect 41679 555932 41790 555934
rect 41679 555929 41745 555932
rect 41922 555255 41982 555814
rect 41871 555250 41982 555255
rect 41871 555194 41876 555250
rect 41932 555194 41982 555250
rect 41871 555192 41982 555194
rect 41871 555189 41937 555192
rect 41730 554367 41790 554926
rect 41730 554362 41841 554367
rect 41730 554306 41780 554362
rect 41836 554306 41841 554362
rect 41730 554304 41841 554306
rect 41775 554301 41841 554304
rect 40962 553626 41022 554186
rect 40954 553562 40960 553626
rect 41024 553562 41030 553626
rect 42114 553035 42174 553298
rect 42063 553030 42174 553035
rect 42063 552974 42068 553030
rect 42124 552974 42174 553030
rect 42063 552972 42174 552974
rect 42063 552969 42129 552972
rect 42306 551999 42366 552558
rect 654447 552144 654513 552147
rect 650208 552142 654513 552144
rect 650208 552086 654452 552142
rect 654508 552086 654513 552142
rect 650208 552084 654513 552086
rect 654447 552081 654513 552084
rect 42306 551994 42417 551999
rect 42306 551938 42356 551994
rect 42412 551938 42417 551994
rect 42306 551936 42417 551938
rect 42351 551933 42417 551936
rect 42927 551700 42993 551703
rect 42336 551698 42993 551700
rect 42336 551642 42932 551698
rect 42988 551642 42993 551698
rect 42336 551640 42993 551642
rect 42927 551637 42993 551640
rect 42831 551108 42897 551111
rect 42336 551106 42897 551108
rect 42336 551050 42836 551106
rect 42892 551050 42897 551106
rect 42336 551048 42897 551050
rect 42831 551045 42897 551048
rect 42114 550075 42174 550190
rect 42114 550070 42225 550075
rect 42114 550014 42164 550070
rect 42220 550014 42225 550070
rect 42114 550012 42225 550014
rect 42159 550009 42225 550012
rect 42306 549332 42366 549376
rect 43023 549332 43089 549335
rect 42306 549330 43089 549332
rect 42306 549274 43028 549330
rect 43084 549274 43089 549330
rect 42306 549272 43089 549274
rect 43023 549269 43089 549272
rect 43119 548592 43185 548595
rect 42336 548590 43185 548592
rect 42336 548534 43124 548590
rect 43180 548534 43185 548590
rect 42336 548532 43185 548534
rect 43119 548529 43185 548532
rect 42306 547260 42366 547748
rect 42306 547200 42750 547260
rect 42690 546816 42750 547200
rect 676858 547050 676864 547114
rect 676928 547112 676934 547114
rect 679791 547112 679857 547115
rect 676928 547110 679857 547112
rect 676928 547054 679796 547110
rect 679852 547054 679857 547110
rect 676928 547052 679857 547054
rect 676928 547050 676934 547052
rect 679791 547049 679857 547052
rect 42306 546756 42750 546816
rect 42306 546298 42366 546756
rect 42639 546298 42705 546301
rect 42306 546296 42705 546298
rect 42306 546268 42644 546296
rect 42336 546240 42644 546268
rect 42700 546240 42705 546296
rect 42336 546238 42705 546240
rect 42639 546235 42705 546238
rect 59535 542228 59601 542231
rect 59535 542226 64416 542228
rect 59535 542170 59540 542226
rect 59596 542170 64416 542226
rect 59535 542168 64416 542170
rect 59535 542165 59601 542168
rect 674754 541639 674814 542050
rect 674703 541634 674814 541639
rect 674703 541578 674708 541634
rect 674764 541578 674814 541634
rect 674703 541576 674814 541578
rect 674703 541573 674769 541576
rect 41871 541340 41937 541343
rect 42682 541340 42688 541342
rect 41871 541338 42688 541340
rect 41871 541282 41876 541338
rect 41932 541282 42688 541338
rect 41871 541280 42688 541282
rect 41871 541277 41937 541280
rect 42682 541278 42688 541280
rect 42752 541278 42758 541342
rect 674415 541340 674481 541343
rect 674415 541338 674784 541340
rect 674415 541282 674420 541338
rect 674476 541282 674784 541338
rect 674415 541280 674784 541282
rect 674415 541277 674481 541280
rect 41967 541192 42033 541195
rect 42106 541192 42112 541194
rect 41967 541190 42112 541192
rect 41967 541134 41972 541190
rect 42028 541134 42112 541190
rect 41967 541132 42112 541134
rect 41967 541129 42033 541132
rect 42106 541130 42112 541132
rect 42176 541130 42182 541194
rect 42063 541044 42129 541047
rect 43066 541044 43072 541046
rect 42063 541042 43072 541044
rect 42063 540986 42068 541042
rect 42124 540986 43072 541042
rect 42063 540984 43072 540986
rect 42063 540981 42129 540984
rect 43066 540982 43072 540984
rect 43136 540982 43142 541046
rect 674703 540748 674769 540751
rect 674703 540746 674814 540748
rect 674703 540690 674708 540746
rect 674764 540690 674814 540746
rect 674703 540685 674814 540690
rect 674754 540422 674814 540685
rect 655119 540304 655185 540307
rect 650208 540302 655185 540304
rect 650208 540246 655124 540302
rect 655180 540246 655185 540302
rect 650208 540244 655185 540246
rect 655119 540241 655185 540244
rect 674703 539860 674769 539863
rect 674703 539858 674814 539860
rect 674703 539802 674708 539858
rect 674764 539802 674814 539858
rect 674703 539797 674814 539802
rect 674754 539682 674814 539797
rect 42063 538974 42129 538975
rect 42063 538972 42112 538974
rect 42020 538970 42112 538972
rect 42020 538914 42068 538970
rect 42020 538912 42112 538914
rect 42063 538910 42112 538912
rect 42176 538910 42182 538974
rect 42063 538909 42129 538910
rect 676674 538679 676734 538794
rect 42682 538614 42688 538678
rect 42752 538676 42758 538678
rect 42927 538676 42993 538679
rect 42752 538674 42993 538676
rect 42752 538618 42932 538674
rect 42988 538618 42993 538674
rect 42752 538616 42993 538618
rect 676674 538674 676785 538679
rect 676674 538618 676724 538674
rect 676780 538618 676785 538674
rect 676674 538616 676785 538618
rect 42752 538614 42758 538616
rect 42927 538613 42993 538616
rect 676719 538613 676785 538616
rect 675514 538380 675520 538382
rect 675330 538320 675520 538380
rect 675330 538158 675390 538320
rect 675514 538318 675520 538320
rect 675584 538318 675590 538382
rect 674784 538128 675390 538158
rect 674754 538098 675360 538128
rect 674754 537643 674814 538098
rect 674754 537638 674865 537643
rect 679791 537640 679857 537643
rect 674754 537582 674804 537638
rect 674860 537582 674865 537638
rect 674754 537580 674865 537582
rect 674799 537577 674865 537580
rect 679746 537638 679857 537640
rect 679746 537582 679796 537638
rect 679852 537582 679857 537638
rect 679746 537577 679857 537582
rect 679746 537314 679806 537577
rect 675706 536986 675712 537050
rect 675776 536986 675782 537050
rect 42831 536900 42897 536903
rect 43066 536900 43072 536902
rect 42831 536898 43072 536900
rect 42831 536842 42836 536898
rect 42892 536842 43072 536898
rect 42831 536840 43072 536842
rect 42831 536837 42897 536840
rect 43066 536838 43072 536840
rect 43136 536838 43142 536902
rect 675714 536500 675774 536986
rect 676666 536246 676672 536310
rect 676736 536246 676742 536310
rect 676674 535686 676734 536246
rect 674362 534840 674368 534904
rect 674432 534902 674438 534904
rect 674432 534842 674784 534902
rect 674432 534840 674438 534842
rect 673978 534026 673984 534090
rect 674048 534088 674054 534090
rect 674048 534028 674784 534088
rect 674048 534026 674054 534028
rect 675898 533730 675904 533794
rect 675968 533730 675974 533794
rect 675906 533392 675966 533730
rect 676090 532694 676096 532758
rect 676160 532694 676166 532758
rect 40954 532546 40960 532610
rect 41024 532608 41030 532610
rect 42639 532608 42705 532611
rect 41024 532606 42705 532608
rect 41024 532550 42644 532606
rect 42700 532550 42705 532606
rect 676098 532578 676158 532694
rect 41024 532548 42705 532550
rect 41024 532546 41030 532548
rect 42639 532545 42705 532548
rect 40570 532250 40576 532314
rect 40640 532312 40646 532314
rect 42735 532312 42801 532315
rect 40640 532310 42801 532312
rect 40640 532254 42740 532310
rect 42796 532254 42801 532310
rect 40640 532252 42801 532254
rect 40640 532250 40646 532252
rect 42735 532249 42801 532252
rect 674554 532250 674560 532314
rect 674624 532312 674630 532314
rect 674624 532252 674814 532312
rect 674624 532250 674630 532252
rect 41775 531722 41841 531723
rect 41722 531658 41728 531722
rect 41792 531720 41841 531722
rect 41792 531718 41884 531720
rect 41836 531662 41884 531718
rect 674754 531690 674814 532252
rect 41792 531660 41884 531662
rect 41792 531658 41841 531660
rect 41775 531657 41841 531658
rect 41871 531278 41937 531279
rect 41871 531276 41920 531278
rect 41828 531274 41920 531276
rect 41828 531218 41876 531274
rect 41828 531216 41920 531218
rect 41871 531214 41920 531216
rect 41984 531214 41990 531278
rect 41871 531213 41937 531214
rect 673839 530980 673905 530983
rect 673839 530978 674784 530980
rect 673839 530922 673844 530978
rect 673900 530922 674784 530978
rect 673839 530920 674784 530922
rect 673839 530917 673905 530920
rect 673839 530092 673905 530095
rect 673839 530090 674784 530092
rect 673839 530034 673844 530090
rect 673900 530034 674784 530090
rect 673839 530032 674784 530034
rect 673839 530029 673905 530032
rect 673839 529352 673905 529355
rect 673839 529350 674784 529352
rect 673839 529294 673844 529350
rect 673900 529294 674784 529350
rect 673839 529292 674784 529294
rect 673839 529289 673905 529292
rect 654447 528612 654513 528615
rect 650208 528610 654513 528612
rect 650208 528554 654452 528610
rect 654508 528554 654513 528610
rect 650208 528552 654513 528554
rect 654447 528549 654513 528552
rect 673743 528612 673809 528615
rect 673743 528610 674784 528612
rect 673743 528554 673748 528610
rect 673804 528554 674784 528610
rect 673743 528552 674784 528554
rect 673743 528549 673809 528552
rect 673839 527872 673905 527875
rect 673839 527870 674784 527872
rect 673839 527814 673844 527870
rect 673900 527814 674784 527870
rect 673839 527812 674784 527814
rect 673839 527809 673905 527812
rect 59439 527576 59505 527579
rect 59439 527574 64416 527576
rect 59439 527518 59444 527574
rect 59500 527518 64416 527574
rect 59439 527516 64416 527518
rect 59439 527513 59505 527516
rect 673743 526984 673809 526987
rect 673743 526982 674784 526984
rect 673743 526926 673748 526982
rect 673804 526926 674784 526982
rect 673743 526924 674784 526926
rect 673743 526921 673809 526924
rect 673839 526244 673905 526247
rect 673839 526242 674784 526244
rect 673839 526186 673844 526242
rect 673900 526186 674784 526242
rect 673839 526184 674784 526186
rect 673839 526181 673905 526184
rect 679746 524767 679806 525326
rect 679746 524762 679857 524767
rect 679746 524706 679796 524762
rect 679852 524706 679857 524762
rect 679746 524704 679857 524706
rect 679791 524701 679857 524704
rect 679791 524172 679857 524175
rect 679746 524170 679857 524172
rect 679746 524114 679796 524170
rect 679852 524114 679857 524170
rect 679746 524109 679857 524114
rect 679746 523846 679806 524109
rect 654447 516920 654513 516923
rect 650208 516918 654513 516920
rect 650208 516862 654452 516918
rect 654508 516862 654513 516918
rect 650208 516860 654513 516862
rect 654447 516857 654513 516860
rect 59535 513368 59601 513371
rect 59535 513366 64416 513368
rect 59535 513310 59540 513366
rect 59596 513310 64416 513366
rect 59535 513308 64416 513310
rect 59535 513305 59601 513308
rect 654447 505228 654513 505231
rect 650208 505226 654513 505228
rect 650208 505170 654452 505226
rect 654508 505170 654513 505226
rect 650208 505168 654513 505170
rect 654447 505165 654513 505168
rect 58095 499012 58161 499015
rect 58095 499010 64416 499012
rect 58095 498954 58100 499010
rect 58156 498954 64416 499010
rect 58095 498952 64416 498954
rect 58095 498949 58161 498952
rect 674754 497831 674814 498094
rect 674703 497826 674814 497831
rect 674703 497770 674708 497826
rect 674764 497770 674814 497826
rect 674703 497768 674814 497770
rect 674703 497765 674769 497768
rect 674415 497310 674481 497313
rect 674415 497308 674784 497310
rect 674415 497252 674420 497308
rect 674476 497252 674784 497308
rect 674415 497250 674784 497252
rect 674415 497247 674481 497250
rect 674415 496496 674481 496499
rect 674415 496494 674784 496496
rect 674415 496438 674420 496494
rect 674476 496438 674784 496494
rect 674415 496436 674784 496438
rect 674415 496433 674481 496436
rect 676719 495904 676785 495907
rect 676674 495902 676785 495904
rect 676674 495846 676724 495902
rect 676780 495846 676785 495902
rect 676674 495841 676785 495846
rect 676674 495578 676734 495841
rect 676674 494575 676734 494838
rect 676674 494570 676785 494575
rect 676674 494514 676724 494570
rect 676780 494514 676785 494570
rect 676674 494512 676785 494514
rect 676719 494509 676785 494512
rect 679695 494424 679761 494427
rect 679695 494422 679806 494424
rect 679695 494366 679700 494422
rect 679756 494366 679806 494422
rect 679695 494361 679806 494366
rect 679746 493536 679806 494361
rect 679887 493536 679953 493539
rect 679746 493534 679953 493536
rect 679746 493478 679892 493534
rect 679948 493478 679953 493534
rect 679746 493476 679953 493478
rect 679887 493473 679953 493476
rect 654447 493388 654513 493391
rect 650208 493386 654513 493388
rect 650208 493330 654452 493386
rect 654508 493330 654513 493386
rect 650208 493328 654513 493330
rect 654447 493325 654513 493328
rect 676674 493095 676734 493358
rect 676623 493090 676734 493095
rect 676623 493034 676628 493090
rect 676684 493034 676734 493090
rect 676623 493032 676734 493034
rect 676623 493029 676689 493032
rect 675130 492734 675136 492798
rect 675200 492734 675206 492798
rect 675138 492470 675198 492734
rect 674607 491908 674673 491911
rect 674607 491906 674814 491908
rect 674607 491850 674612 491906
rect 674668 491850 674814 491906
rect 674607 491848 674814 491850
rect 674607 491845 674673 491848
rect 674754 491730 674814 491848
rect 674938 491402 674944 491466
rect 675008 491402 675014 491466
rect 674946 490842 675006 491402
rect 674223 490132 674289 490135
rect 674223 490130 674784 490132
rect 674223 490074 674228 490130
rect 674284 490074 674784 490130
rect 674223 490072 674784 490074
rect 674223 490069 674289 490072
rect 674511 489688 674577 489691
rect 674511 489686 674814 489688
rect 674511 489630 674516 489686
rect 674572 489630 674814 489686
rect 674511 489628 674814 489630
rect 674511 489625 674577 489628
rect 674754 489362 674814 489628
rect 674895 488800 674961 488803
rect 674895 488798 675006 488800
rect 674895 488742 674900 488798
rect 674956 488742 675006 488798
rect 674895 488737 675006 488742
rect 674946 488622 675006 488737
rect 674170 487702 674176 487766
rect 674240 487764 674246 487766
rect 674240 487704 674784 487764
rect 674240 487702 674246 487704
rect 674746 487406 674752 487470
rect 674816 487406 674822 487470
rect 674754 486920 674814 487406
rect 674031 486136 674097 486139
rect 674031 486134 674784 486136
rect 674031 486078 674036 486134
rect 674092 486078 674784 486134
rect 674031 486076 674784 486078
rect 674031 486073 674097 486076
rect 674319 485322 674385 485325
rect 674319 485320 674784 485322
rect 674319 485264 674324 485320
rect 674380 485264 674784 485320
rect 674319 485262 674784 485264
rect 674319 485259 674385 485262
rect 674127 484656 674193 484659
rect 674127 484654 674784 484656
rect 674127 484598 674132 484654
rect 674188 484598 674784 484654
rect 674127 484596 674784 484598
rect 674127 484593 674193 484596
rect 59535 484508 59601 484511
rect 59535 484506 64416 484508
rect 59535 484450 59540 484506
rect 59596 484450 64416 484506
rect 59535 484448 64416 484450
rect 59535 484445 59601 484448
rect 676282 484002 676288 484066
rect 676352 484002 676358 484066
rect 676290 483812 676350 484002
rect 674991 483176 675057 483179
rect 674946 483174 675057 483176
rect 674946 483118 674996 483174
rect 675052 483118 675057 483174
rect 674946 483113 675057 483118
rect 674946 482998 675006 483113
rect 675087 482436 675153 482439
rect 675087 482434 675198 482436
rect 675087 482378 675092 482434
rect 675148 482378 675198 482434
rect 675087 482373 675198 482378
rect 675138 482184 675198 482373
rect 654447 481696 654513 481699
rect 650208 481694 654513 481696
rect 650208 481638 654452 481694
rect 654508 481638 654513 481694
rect 650208 481636 654513 481638
rect 654447 481633 654513 481636
rect 679746 480811 679806 481370
rect 679746 480806 679857 480811
rect 679746 480750 679796 480806
rect 679852 480750 679857 480806
rect 679746 480748 679857 480750
rect 679791 480745 679857 480748
rect 679791 480068 679857 480071
rect 679746 480066 679857 480068
rect 679746 480010 679796 480066
rect 679852 480010 679857 480066
rect 679746 480005 679857 480010
rect 679746 479890 679806 480005
rect 673978 475270 673984 475334
rect 674048 475332 674054 475334
rect 679887 475332 679953 475335
rect 674048 475330 679953 475332
rect 674048 475274 679892 475330
rect 679948 475274 679953 475330
rect 674048 475272 679953 475274
rect 674048 475270 674054 475272
rect 679887 475269 679953 475272
rect 59535 470300 59601 470303
rect 59535 470298 64416 470300
rect 59535 470242 59540 470298
rect 59596 470242 64416 470298
rect 59535 470240 64416 470242
rect 59535 470237 59601 470240
rect 654447 470004 654513 470007
rect 650208 470002 654513 470004
rect 650208 469946 654452 470002
rect 654508 469946 654513 470002
rect 650208 469944 654513 469946
rect 654447 469941 654513 469944
rect 654351 458312 654417 458315
rect 650208 458310 654417 458312
rect 650208 458254 654356 458310
rect 654412 458254 654417 458310
rect 650208 458252 654417 458254
rect 654351 458249 654417 458252
rect 59535 455796 59601 455799
rect 59535 455794 64416 455796
rect 59535 455738 59540 455794
rect 59596 455738 64416 455794
rect 59535 455736 64416 455738
rect 59535 455733 59601 455736
rect 654447 446472 654513 446475
rect 650208 446470 654513 446472
rect 650208 446414 654452 446470
rect 654508 446414 654513 446470
rect 650208 446412 654513 446414
rect 654447 446409 654513 446412
rect 59535 441440 59601 441443
rect 59535 441438 64416 441440
rect 59535 441382 59540 441438
rect 59596 441382 64416 441438
rect 59535 441380 64416 441382
rect 59535 441377 59601 441380
rect 42639 436926 42705 436929
rect 42336 436924 42705 436926
rect 42336 436868 42644 436924
rect 42700 436868 42705 436924
rect 42336 436866 42705 436868
rect 42639 436863 42705 436866
rect 42639 436112 42705 436115
rect 42336 436110 42705 436112
rect 42336 436054 42644 436110
rect 42700 436054 42705 436110
rect 42336 436052 42705 436054
rect 42639 436049 42705 436052
rect 42351 435520 42417 435523
rect 42306 435518 42417 435520
rect 42306 435462 42356 435518
rect 42412 435462 42417 435518
rect 42306 435457 42417 435462
rect 42306 435194 42366 435457
rect 654351 434780 654417 434783
rect 650208 434778 654417 434780
rect 650208 434722 654356 434778
rect 654412 434722 654417 434778
rect 650208 434720 654417 434722
rect 654351 434717 654417 434720
rect 43407 434484 43473 434487
rect 42336 434482 43473 434484
rect 42336 434426 43412 434482
rect 43468 434426 43473 434482
rect 42336 434424 43473 434426
rect 43407 434421 43473 434424
rect 43215 433596 43281 433599
rect 42336 433594 43281 433596
rect 42336 433538 43220 433594
rect 43276 433538 43281 433594
rect 42336 433536 43281 433538
rect 43215 433533 43281 433536
rect 43791 433004 43857 433007
rect 42144 433002 43857 433004
rect 42144 432974 43796 433002
rect 42114 432946 43796 432974
rect 43852 432946 43857 433002
rect 42114 432944 43857 432946
rect 42114 432710 42174 432944
rect 43791 432941 43857 432944
rect 42106 432646 42112 432710
rect 42176 432646 42182 432710
rect 43599 432116 43665 432119
rect 40608 432114 43665 432116
rect 40608 432086 43604 432114
rect 40578 432058 43604 432086
rect 43660 432058 43665 432114
rect 40578 432056 43665 432058
rect 40578 431970 40638 432056
rect 43599 432053 43665 432056
rect 40570 431906 40576 431970
rect 40640 431906 40646 431970
rect 40962 430786 41022 431346
rect 40954 430722 40960 430786
rect 41024 430722 41030 430786
rect 41922 429899 41982 430458
rect 41871 429894 41982 429899
rect 41871 429838 41876 429894
rect 41932 429838 41982 429894
rect 41871 429836 41982 429838
rect 41871 429833 41937 429836
rect 40770 429454 40830 429718
rect 40762 429390 40768 429454
rect 40832 429390 40838 429454
rect 41346 428418 41406 428830
rect 41338 428354 41344 428418
rect 41408 428354 41414 428418
rect 41538 427678 41598 428238
rect 41530 427614 41536 427678
rect 41600 427614 41606 427678
rect 41730 426791 41790 427350
rect 59343 427084 59409 427087
rect 59343 427082 64416 427084
rect 59343 427026 59348 427082
rect 59404 427026 64416 427082
rect 59343 427024 64416 427026
rect 59343 427021 59409 427024
rect 41730 426786 41841 426791
rect 41730 426730 41780 426786
rect 41836 426730 41841 426786
rect 41730 426728 41841 426730
rect 41775 426725 41841 426728
rect 41154 426346 41214 426536
rect 41146 426282 41152 426346
rect 41216 426282 41222 426346
rect 40386 425162 40446 425722
rect 40378 425098 40384 425162
rect 40448 425098 40454 425162
rect 42306 424420 42366 424908
rect 43119 424420 43185 424423
rect 42306 424418 43185 424420
rect 42306 424362 43124 424418
rect 43180 424362 43185 424418
rect 42306 424360 43185 424362
rect 43119 424357 43185 424360
rect 42735 424124 42801 424127
rect 42336 424122 42801 424124
rect 42336 424066 42740 424122
rect 42796 424066 42801 424122
rect 42336 424064 42801 424066
rect 42735 424061 42801 424064
rect 42114 423239 42174 423428
rect 42114 423234 42225 423239
rect 42114 423178 42164 423234
rect 42220 423178 42225 423234
rect 42114 423176 42225 423178
rect 42159 423173 42225 423176
rect 654447 423088 654513 423091
rect 650208 423086 654513 423088
rect 650208 423030 654452 423086
rect 654508 423030 654513 423086
rect 650208 423028 654513 423030
rect 654447 423025 654513 423028
rect 42927 422644 42993 422647
rect 42336 422642 42993 422644
rect 42336 422586 42932 422642
rect 42988 422586 42993 422642
rect 42336 422584 42993 422586
rect 42927 422581 42993 422584
rect 42306 421312 42366 421800
rect 43023 421312 43089 421315
rect 42306 421310 43089 421312
rect 42306 421254 43028 421310
rect 43084 421254 43089 421310
rect 42306 421252 43089 421254
rect 43023 421249 43089 421252
rect 42831 421016 42897 421019
rect 42336 421014 42897 421016
rect 42336 420958 42836 421014
rect 42892 420958 42897 421014
rect 42336 420956 42897 420958
rect 42831 420953 42897 420956
rect 42639 420128 42705 420131
rect 42336 420126 42705 420128
rect 42336 420070 42644 420126
rect 42700 420070 42705 420126
rect 42336 420068 42705 420070
rect 42639 420065 42705 420068
rect 41722 419030 41728 419094
rect 41792 419092 41798 419094
rect 42298 419092 42304 419094
rect 41792 419032 42304 419092
rect 41792 419030 41798 419032
rect 42298 419030 42304 419032
rect 42368 419030 42374 419094
rect 42639 418648 42705 418651
rect 42336 418646 42705 418648
rect 42336 418590 42644 418646
rect 42700 418590 42705 418646
rect 42336 418588 42705 418590
rect 42639 418585 42705 418588
rect 57807 412728 57873 412731
rect 57807 412726 64416 412728
rect 57807 412670 57812 412726
rect 57868 412670 64416 412726
rect 57807 412668 64416 412670
rect 57807 412665 57873 412668
rect 676623 411990 676689 411991
rect 676623 411986 676672 411990
rect 676736 411988 676742 411990
rect 676623 411930 676628 411986
rect 676623 411926 676672 411930
rect 676736 411928 676780 411988
rect 676736 411926 676742 411928
rect 676623 411925 676689 411926
rect 655023 411248 655089 411251
rect 650208 411246 655089 411248
rect 650208 411190 655028 411246
rect 655084 411190 655089 411246
rect 650208 411188 655089 411190
rect 655023 411185 655089 411188
rect 674415 409916 674481 409919
rect 674415 409914 674784 409916
rect 674415 409858 674420 409914
rect 674476 409858 674784 409914
rect 674415 409856 674784 409858
rect 674415 409853 674481 409856
rect 674703 409324 674769 409327
rect 674703 409322 674814 409324
rect 674703 409266 674708 409322
rect 674764 409266 674814 409322
rect 674703 409261 674814 409266
rect 674754 409072 674814 409261
rect 674703 408436 674769 408439
rect 674703 408434 674814 408436
rect 674703 408378 674708 408434
rect 674764 408378 674814 408434
rect 674703 408373 674814 408378
rect 674754 408258 674814 408373
rect 676719 407696 676785 407699
rect 676674 407694 676785 407696
rect 676674 407638 676724 407694
rect 676780 407638 676785 407694
rect 676674 407633 676785 407638
rect 676674 407444 676734 407633
rect 673839 406660 673905 406663
rect 673839 406658 674784 406660
rect 673839 406602 673844 406658
rect 673900 406602 674784 406658
rect 673839 406600 674784 406602
rect 673839 406597 673905 406600
rect 41530 406006 41536 406070
rect 41600 406068 41606 406070
rect 41775 406068 41841 406071
rect 41600 406066 41841 406068
rect 41600 406010 41780 406066
rect 41836 406010 41841 406066
rect 41600 406008 41841 406010
rect 41600 406006 41606 406008
rect 41775 406005 41841 406008
rect 673978 405858 673984 405922
rect 674048 405920 674054 405922
rect 674048 405860 674784 405920
rect 674048 405858 674054 405860
rect 675322 405266 675328 405330
rect 675392 405328 675398 405330
rect 676666 405328 676672 405330
rect 675392 405268 676672 405328
rect 675392 405266 675398 405268
rect 676666 405266 676672 405268
rect 676736 405266 676742 405330
rect 676674 405150 676734 405266
rect 41775 404294 41841 404295
rect 41722 404230 41728 404294
rect 41792 404292 41841 404294
rect 42298 404292 42304 404294
rect 41792 404290 42304 404292
rect 41836 404234 42304 404290
rect 41792 404232 42304 404234
rect 41792 404230 41841 404232
rect 42298 404230 42304 404232
rect 42368 404230 42374 404294
rect 41775 404229 41841 404230
rect 674946 404147 675006 404262
rect 674895 404142 675006 404147
rect 674895 404086 674900 404142
rect 674956 404086 675006 404142
rect 674895 404084 675006 404086
rect 674895 404081 674961 404084
rect 41530 403786 41536 403850
rect 41600 403848 41606 403850
rect 42063 403848 42129 403851
rect 42682 403848 42688 403850
rect 41600 403846 42688 403848
rect 41600 403790 42068 403846
rect 42124 403790 42688 403846
rect 41600 403788 42688 403790
rect 41600 403786 41606 403788
rect 42063 403785 42129 403788
rect 42682 403786 42688 403788
rect 42752 403786 42758 403850
rect 674170 403490 674176 403554
rect 674240 403552 674246 403554
rect 674240 403492 674784 403552
rect 674240 403490 674246 403492
rect 675330 402519 675390 402634
rect 40378 402454 40384 402518
rect 40448 402516 40454 402518
rect 41775 402516 41841 402519
rect 40448 402514 41841 402516
rect 40448 402458 41780 402514
rect 41836 402458 41841 402514
rect 40448 402456 41841 402458
rect 675330 402514 675441 402519
rect 675330 402458 675380 402514
rect 675436 402458 675441 402514
rect 675330 402456 675441 402458
rect 40448 402454 40454 402456
rect 41775 402453 41841 402456
rect 675375 402453 675441 402456
rect 41338 402010 41344 402074
rect 41408 402072 41414 402074
rect 41775 402072 41841 402075
rect 41408 402070 41841 402072
rect 41408 402014 41780 402070
rect 41836 402014 41841 402070
rect 41408 402012 41841 402014
rect 41408 402010 41414 402012
rect 41775 402009 41841 402012
rect 674127 401924 674193 401927
rect 674127 401922 674784 401924
rect 674127 401866 674132 401922
rect 674188 401866 674784 401922
rect 674127 401864 674784 401866
rect 674127 401861 674193 401864
rect 674554 400530 674560 400594
rect 674624 400592 674630 400594
rect 674754 400592 674814 401154
rect 674624 400532 674814 400592
rect 674624 400530 674630 400532
rect 674362 400382 674368 400446
rect 674432 400444 674438 400446
rect 674432 400384 674784 400444
rect 674432 400382 674438 400384
rect 40954 400086 40960 400150
rect 41024 400148 41030 400150
rect 41775 400148 41841 400151
rect 41024 400146 41841 400148
rect 41024 400090 41780 400146
rect 41836 400090 41841 400146
rect 41024 400088 41841 400090
rect 41024 400086 41030 400088
rect 41775 400085 41841 400088
rect 41146 399494 41152 399558
rect 41216 399556 41222 399558
rect 41775 399556 41841 399559
rect 654447 399556 654513 399559
rect 41216 399554 41841 399556
rect 41216 399498 41780 399554
rect 41836 399498 41841 399554
rect 41216 399496 41841 399498
rect 650208 399554 654513 399556
rect 650208 399498 654452 399554
rect 654508 399498 654513 399554
rect 650208 399496 654513 399498
rect 41216 399494 41222 399496
rect 41775 399493 41841 399496
rect 654447 399493 654513 399496
rect 675330 399411 675390 399526
rect 675279 399406 675390 399411
rect 675279 399350 675284 399406
rect 675340 399350 675390 399406
rect 675279 399348 675390 399350
rect 675279 399345 675345 399348
rect 40762 398754 40768 398818
rect 40832 398816 40838 398818
rect 41775 398816 41841 398819
rect 40832 398814 41841 398816
rect 40832 398758 41780 398814
rect 41836 398758 41841 398814
rect 40832 398756 41841 398758
rect 40832 398754 40838 398756
rect 41775 398753 41841 398756
rect 674607 398520 674673 398523
rect 674754 398520 674814 398786
rect 674607 398518 674814 398520
rect 674607 398462 674612 398518
rect 674668 398462 674814 398518
rect 674607 398460 674814 398462
rect 674607 398457 674673 398460
rect 59055 398372 59121 398375
rect 59055 398370 64416 398372
rect 59055 398314 59060 398370
rect 59116 398314 64416 398370
rect 59055 398312 64416 398314
rect 59055 398309 59121 398312
rect 674319 397928 674385 397931
rect 674319 397926 674784 397928
rect 674319 397870 674324 397926
rect 674380 397870 674784 397926
rect 674319 397868 674784 397870
rect 674319 397865 674385 397868
rect 674031 397188 674097 397191
rect 674031 397186 674784 397188
rect 674031 397130 674036 397186
rect 674092 397130 674784 397186
rect 674031 397128 674784 397130
rect 674031 397125 674097 397128
rect 674415 396448 674481 396451
rect 674415 396446 674784 396448
rect 674415 396390 674420 396446
rect 674476 396390 674784 396446
rect 674415 396388 674784 396390
rect 674415 396385 674481 396388
rect 674754 395415 674814 395604
rect 674754 395410 674865 395415
rect 674754 395354 674804 395410
rect 674860 395354 674865 395410
rect 674754 395352 674865 395354
rect 674799 395349 674865 395352
rect 674754 394527 674814 394790
rect 674703 394522 674814 394527
rect 674703 394466 674708 394522
rect 674764 394466 674814 394522
rect 674703 394464 674814 394466
rect 674703 394461 674769 394464
rect 42351 393932 42417 393935
rect 42306 393930 42417 393932
rect 42306 393874 42356 393930
rect 42412 393874 42417 393930
rect 42306 393869 42417 393874
rect 42306 393680 42366 393869
rect 674511 393784 674577 393787
rect 674754 393784 674814 393976
rect 674511 393782 674814 393784
rect 674511 393726 674516 393782
rect 674572 393726 674814 393782
rect 674511 393724 674814 393726
rect 674511 393721 674577 393724
rect 42351 393192 42417 393195
rect 42306 393190 42417 393192
rect 42306 393134 42356 393190
rect 42412 393134 42417 393190
rect 42306 393129 42417 393134
rect 42306 392866 42366 393129
rect 679746 392603 679806 393162
rect 679746 392598 679857 392603
rect 679746 392542 679796 392598
rect 679852 392542 679857 392598
rect 679746 392540 679857 392542
rect 679791 392537 679857 392540
rect 42351 392304 42417 392307
rect 42306 392302 42417 392304
rect 42306 392246 42356 392302
rect 42412 392246 42417 392302
rect 42306 392241 42417 392246
rect 42306 392052 42366 392241
rect 679791 392156 679857 392159
rect 679746 392154 679857 392156
rect 679746 392098 679796 392154
rect 679852 392098 679857 392154
rect 679746 392093 679857 392098
rect 679746 391682 679806 392093
rect 43215 391268 43281 391271
rect 42336 391266 43281 391268
rect 42336 391210 43220 391266
rect 43276 391210 43281 391266
rect 42336 391208 43281 391210
rect 43215 391205 43281 391208
rect 43311 390972 43377 390975
rect 42306 390970 43377 390972
rect 42306 390914 43316 390970
rect 43372 390914 43377 390970
rect 42306 390912 43377 390914
rect 42306 390424 42366 390912
rect 43311 390909 43377 390912
rect 42106 390170 42112 390234
rect 42176 390170 42182 390234
rect 42114 389788 42174 390170
rect 42114 389758 42336 389788
rect 42144 389728 42366 389758
rect 42306 389492 42366 389728
rect 42490 389492 42496 389494
rect 42306 389432 42496 389492
rect 42490 389430 42496 389432
rect 42560 389430 42566 389494
rect 40578 388606 40638 388870
rect 40570 388542 40576 388606
rect 40640 388542 40646 388606
rect 40962 387570 41022 388130
rect 653871 387864 653937 387867
rect 650208 387862 653937 387864
rect 650208 387806 653876 387862
rect 653932 387806 653937 387862
rect 650208 387804 653937 387806
rect 653871 387801 653937 387804
rect 40954 387506 40960 387570
rect 41024 387506 41030 387570
rect 42114 386683 42174 387242
rect 42063 386678 42174 386683
rect 42063 386622 42068 386678
rect 42124 386622 42174 386678
rect 42063 386620 42174 386622
rect 42063 386617 42129 386620
rect 40770 386090 40830 386502
rect 40762 386026 40768 386090
rect 40832 386026 40838 386090
rect 41346 385202 41406 385614
rect 41338 385138 41344 385202
rect 41408 385138 41414 385202
rect 41538 384462 41598 385022
rect 41530 384398 41536 384462
rect 41600 384398 41606 384462
rect 42306 383575 42366 384134
rect 59535 384016 59601 384019
rect 59535 384014 64416 384016
rect 59535 383958 59540 384014
rect 59596 383958 64416 384014
rect 59535 383956 64416 383958
rect 59535 383953 59601 383956
rect 42306 383570 42417 383575
rect 42306 383514 42356 383570
rect 42412 383514 42417 383570
rect 42306 383512 42417 383514
rect 42351 383509 42417 383512
rect 41154 383130 41214 383394
rect 41146 383066 41152 383130
rect 41216 383066 41222 383130
rect 42114 381946 42174 382506
rect 42106 381882 42112 381946
rect 42176 381882 42182 381946
rect 42831 381796 42897 381799
rect 42336 381794 42897 381796
rect 42336 381738 42836 381794
rect 42892 381738 42897 381794
rect 42336 381736 42897 381738
rect 42831 381733 42897 381736
rect 43023 380908 43089 380911
rect 42336 380906 43089 380908
rect 42336 380850 43028 380906
rect 43084 380850 43089 380906
rect 42336 380848 43089 380850
rect 43023 380845 43089 380848
rect 37314 380023 37374 380212
rect 37314 380018 37425 380023
rect 37314 379962 37364 380018
rect 37420 379962 37425 380018
rect 37314 379960 37425 379962
rect 37359 379957 37425 379960
rect 42306 378839 42366 379398
rect 42255 378834 42366 378839
rect 42255 378778 42260 378834
rect 42316 378778 42366 378834
rect 42255 378776 42366 378778
rect 42255 378773 42321 378776
rect 674554 378774 674560 378838
rect 674624 378836 674630 378838
rect 675471 378836 675537 378839
rect 674624 378834 675537 378836
rect 674624 378778 675476 378834
rect 675532 378778 675537 378834
rect 674624 378776 675537 378778
rect 674624 378774 674630 378776
rect 675471 378773 675537 378776
rect 42306 378540 42366 378584
rect 43119 378540 43185 378543
rect 42306 378538 43185 378540
rect 42306 378482 43124 378538
rect 43180 378482 43185 378538
rect 42306 378480 43185 378482
rect 43119 378477 43185 378480
rect 42735 377800 42801 377803
rect 42336 377798 42801 377800
rect 42336 377742 42740 377798
rect 42796 377742 42801 377798
rect 42336 377740 42801 377742
rect 42735 377737 42801 377740
rect 42114 376619 42174 376956
rect 42114 376614 42225 376619
rect 42114 376558 42164 376614
rect 42220 376558 42225 376614
rect 42114 376556 42225 376558
rect 42159 376553 42225 376556
rect 654159 376172 654225 376175
rect 650208 376170 654225 376172
rect 650208 376114 654164 376170
rect 654220 376114 654225 376170
rect 650208 376112 654225 376114
rect 654159 376109 654225 376112
rect 42114 375287 42174 375402
rect 42114 375282 42225 375287
rect 42114 375226 42164 375282
rect 42220 375226 42225 375282
rect 42114 375224 42225 375226
rect 42159 375221 42225 375224
rect 675087 374544 675153 374547
rect 675514 374544 675520 374546
rect 675087 374542 675520 374544
rect 675087 374486 675092 374542
rect 675148 374486 675520 374542
rect 675087 374484 675520 374486
rect 675087 374481 675153 374484
rect 675514 374482 675520 374484
rect 675584 374482 675590 374546
rect 674170 373890 674176 373954
rect 674240 373952 674246 373954
rect 675471 373952 675537 373955
rect 674240 373950 675537 373952
rect 674240 373894 675476 373950
rect 675532 373894 675537 373950
rect 674240 373892 675537 373894
rect 674240 373890 674246 373892
rect 675471 373889 675537 373892
rect 674362 371966 674368 372030
rect 674432 372028 674438 372030
rect 675375 372028 675441 372031
rect 674432 372026 675441 372028
rect 674432 371970 675380 372026
rect 675436 371970 675441 372026
rect 674432 371968 675441 371970
rect 674432 371966 674438 371968
rect 675375 371965 675441 371968
rect 675183 371584 675249 371587
rect 675706 371584 675712 371586
rect 675183 371582 675712 371584
rect 675183 371526 675188 371582
rect 675244 371526 675712 371582
rect 675183 371524 675712 371526
rect 675183 371521 675249 371524
rect 675706 371522 675712 371524
rect 675776 371522 675782 371586
rect 59535 369660 59601 369663
rect 59535 369658 64416 369660
rect 59535 369602 59540 369658
rect 59596 369602 64416 369658
rect 59535 369600 64416 369602
rect 59535 369597 59601 369600
rect 40570 368710 40576 368774
rect 40640 368772 40646 368774
rect 40640 368712 41790 368772
rect 40640 368710 40646 368712
rect 41730 368626 41790 368712
rect 42106 368710 42112 368774
rect 42176 368710 42182 368774
rect 41722 368562 41728 368626
rect 41792 368562 41798 368626
rect 42114 368478 42174 368710
rect 42106 368414 42112 368478
rect 42176 368414 42182 368478
rect 41914 368266 41920 368330
rect 41984 368328 41990 368330
rect 42298 368328 42304 368330
rect 41984 368268 42304 368328
rect 41984 368266 41990 368268
rect 42298 368266 42304 368268
rect 42368 368266 42374 368330
rect 674754 364483 674814 364672
rect 674703 364478 674814 364483
rect 674703 364422 674708 364478
rect 674764 364422 674814 364478
rect 674703 364420 674814 364422
rect 674703 364417 674769 364420
rect 654447 364332 654513 364335
rect 650208 364330 654513 364332
rect 650208 364274 654452 364330
rect 654508 364274 654513 364330
rect 650208 364272 654513 364274
rect 654447 364269 654513 364272
rect 674415 363888 674481 363891
rect 674415 363886 674784 363888
rect 674415 363830 674420 363886
rect 674476 363830 674784 363886
rect 674415 363828 674784 363830
rect 674415 363825 674481 363828
rect 674607 363296 674673 363299
rect 674607 363294 674814 363296
rect 674607 363238 674612 363294
rect 674668 363238 674814 363294
rect 674607 363236 674814 363238
rect 674607 363233 674673 363236
rect 41722 363148 41728 363150
rect 40386 363088 41728 363148
rect 40386 363002 40446 363088
rect 41722 363086 41728 363088
rect 41792 363086 41798 363150
rect 674754 363044 674814 363236
rect 40378 362938 40384 363002
rect 40448 362938 40454 363002
rect 41530 362790 41536 362854
rect 41600 362852 41606 362854
rect 41775 362852 41841 362855
rect 41600 362850 41841 362852
rect 41600 362794 41780 362850
rect 41836 362794 41841 362850
rect 41600 362792 41841 362794
rect 41600 362790 41606 362792
rect 41775 362789 41841 362792
rect 673839 362260 673905 362263
rect 673839 362258 674784 362260
rect 673839 362202 673844 362258
rect 673900 362202 674784 362258
rect 673839 362200 674784 362202
rect 673839 362197 673905 362200
rect 674170 361384 674176 361448
rect 674240 361446 674246 361448
rect 674240 361386 674784 361446
rect 674240 361384 674246 361386
rect 42063 360928 42129 360931
rect 42298 360928 42304 360930
rect 42063 360926 42304 360928
rect 42063 360870 42068 360926
rect 42124 360870 42304 360926
rect 42063 360868 42304 360870
rect 42063 360865 42129 360868
rect 42298 360866 42304 360868
rect 42368 360866 42374 360930
rect 673978 360718 673984 360782
rect 674048 360780 674054 360782
rect 674048 360750 679776 360780
rect 674048 360720 679806 360750
rect 674048 360718 674054 360720
rect 41775 360634 41841 360635
rect 41722 360570 41728 360634
rect 41792 360632 41841 360634
rect 42682 360632 42688 360634
rect 41792 360630 42688 360632
rect 41836 360574 42688 360630
rect 41792 360572 42688 360574
rect 41792 360570 41841 360572
rect 42682 360570 42688 360572
rect 42752 360570 42758 360634
rect 41775 360569 41841 360570
rect 675322 360126 675328 360190
rect 675392 360188 675398 360190
rect 675898 360188 675904 360190
rect 675392 360128 675904 360188
rect 675392 360126 675398 360128
rect 675898 360126 675904 360128
rect 675968 360126 675974 360190
rect 679746 360188 679806 360720
rect 679887 360188 679953 360191
rect 679746 360186 679953 360188
rect 679746 360130 679892 360186
rect 679948 360130 679953 360186
rect 679746 360128 679953 360130
rect 675330 359936 675390 360126
rect 679887 360125 679953 360128
rect 42063 359450 42129 359451
rect 42063 359446 42112 359450
rect 42176 359448 42182 359450
rect 42063 359390 42068 359446
rect 42063 359386 42112 359390
rect 42176 359388 42220 359448
rect 42176 359386 42182 359388
rect 42063 359385 42129 359386
rect 674031 359152 674097 359155
rect 674031 359150 674784 359152
rect 674031 359094 674036 359150
rect 674092 359094 674784 359150
rect 674031 359092 674784 359094
rect 674031 359089 674097 359092
rect 41338 358646 41344 358710
rect 41408 358708 41414 358710
rect 41775 358708 41841 358711
rect 41408 358706 41841 358708
rect 41408 358650 41780 358706
rect 41836 358650 41841 358706
rect 41408 358648 41841 358650
rect 41408 358646 41414 358648
rect 41775 358645 41841 358648
rect 674362 358202 674368 358266
rect 674432 358264 674438 358266
rect 674432 358204 674784 358264
rect 674432 358202 674438 358204
rect 674511 357228 674577 357231
rect 674754 357228 674814 357494
rect 674511 357226 674814 357228
rect 674511 357170 674516 357226
rect 674572 357170 674814 357226
rect 674511 357168 674814 357170
rect 674511 357165 674577 357168
rect 40954 356870 40960 356934
rect 41024 356932 41030 356934
rect 41871 356932 41937 356935
rect 41024 356930 41937 356932
rect 41024 356874 41876 356930
rect 41932 356874 41937 356930
rect 41024 356872 41937 356874
rect 41024 356870 41030 356872
rect 41871 356869 41937 356872
rect 675138 356491 675198 356606
rect 41146 356426 41152 356490
rect 41216 356488 41222 356490
rect 41775 356488 41841 356491
rect 41216 356486 41841 356488
rect 41216 356430 41780 356486
rect 41836 356430 41841 356486
rect 41216 356428 41841 356430
rect 675138 356486 675249 356491
rect 675138 356430 675188 356486
rect 675244 356430 675249 356486
rect 675138 356428 675249 356430
rect 41216 356426 41222 356428
rect 41775 356425 41841 356428
rect 675183 356425 675249 356428
rect 40762 355538 40768 355602
rect 40832 355600 40838 355602
rect 41775 355600 41841 355603
rect 40832 355598 41841 355600
rect 40832 355542 41780 355598
rect 41836 355542 41841 355598
rect 40832 355540 41841 355542
rect 40832 355538 40838 355540
rect 41775 355537 41841 355540
rect 674754 355454 674814 356014
rect 674746 355390 674752 355454
rect 674816 355390 674822 355454
rect 58959 355304 59025 355307
rect 58959 355302 64416 355304
rect 58959 355246 58964 355302
rect 59020 355246 64416 355302
rect 58959 355244 64416 355246
rect 58959 355241 59025 355244
rect 674554 354502 674560 354566
rect 674624 354564 674630 354566
rect 674754 354564 674814 355126
rect 674624 354504 674814 354564
rect 674624 354502 674630 354504
rect 675330 354123 675390 354386
rect 675279 354118 675390 354123
rect 675279 354062 675284 354118
rect 675340 354062 675390 354118
rect 675279 354060 675390 354062
rect 675279 354057 675345 354060
rect 675138 353383 675198 353498
rect 675087 353378 675198 353383
rect 675087 353322 675092 353378
rect 675148 353322 675198 353378
rect 675087 353320 675198 353322
rect 675087 353317 675153 353320
rect 674319 352788 674385 352791
rect 674319 352786 674784 352788
rect 674319 352730 674324 352786
rect 674380 352730 674784 352786
rect 674319 352728 674784 352730
rect 674319 352725 674385 352728
rect 655311 352640 655377 352643
rect 650208 352638 655377 352640
rect 650208 352582 655316 352638
rect 655372 352582 655377 352638
rect 650208 352580 655377 352582
rect 655311 352577 655377 352580
rect 675138 351458 675198 351870
rect 675130 351394 675136 351458
rect 675200 351394 675206 351458
rect 674223 351308 674289 351311
rect 674223 351306 674784 351308
rect 674223 351250 674228 351306
rect 674284 351250 674784 351306
rect 674223 351248 674784 351250
rect 674223 351245 674289 351248
rect 42351 350716 42417 350719
rect 42306 350714 42417 350716
rect 42306 350658 42356 350714
rect 42412 350658 42417 350714
rect 42306 350653 42417 350658
rect 42306 350538 42366 350653
rect 674946 350275 675006 350390
rect 674895 350270 675006 350275
rect 674895 350214 674900 350270
rect 674956 350214 675006 350270
rect 674895 350212 675006 350214
rect 674895 350209 674961 350212
rect 42639 349680 42705 349683
rect 42336 349678 42705 349680
rect 42336 349622 42644 349678
rect 42700 349622 42705 349678
rect 42336 349620 42705 349622
rect 42639 349617 42705 349620
rect 674754 349387 674814 349576
rect 674703 349382 674814 349387
rect 674703 349326 674708 349382
rect 674764 349326 674814 349382
rect 674703 349324 674814 349326
rect 674703 349321 674769 349324
rect 42351 349088 42417 349091
rect 42306 349086 42417 349088
rect 42306 349030 42356 349086
rect 42412 349030 42417 349086
rect 42306 349025 42417 349030
rect 42306 348910 42366 349025
rect 674946 348647 675006 348762
rect 674946 348642 675057 348647
rect 674946 348586 674996 348642
rect 675052 348586 675057 348642
rect 674946 348584 675057 348586
rect 674991 348581 675057 348584
rect 43311 348052 43377 348055
rect 42336 348050 43377 348052
rect 42336 347994 43316 348050
rect 43372 347994 43377 348050
rect 42336 347992 43377 347994
rect 43311 347989 43377 347992
rect 43215 347756 43281 347759
rect 42306 347754 43281 347756
rect 42306 347698 43220 347754
rect 43276 347698 43281 347754
rect 42306 347696 43281 347698
rect 42306 347208 42366 347696
rect 43215 347693 43281 347696
rect 679746 347463 679806 347948
rect 679746 347458 679857 347463
rect 679746 347402 679796 347458
rect 679852 347402 679857 347458
rect 679746 347400 679857 347402
rect 679791 347397 679857 347400
rect 42490 346868 42496 346870
rect 42306 346808 42496 346868
rect 42306 346572 42366 346808
rect 42490 346806 42496 346808
rect 42560 346806 42566 346870
rect 679791 346720 679857 346723
rect 42144 346542 42366 346572
rect 679746 346718 679857 346720
rect 679746 346662 679796 346718
rect 679852 346662 679857 346718
rect 679746 346657 679857 346662
rect 42114 346512 42336 346542
rect 42114 346130 42174 346512
rect 679746 346468 679806 346657
rect 42106 346066 42112 346130
rect 42176 346066 42182 346130
rect 41338 345918 41344 345982
rect 41408 345980 41414 345982
rect 42298 345980 42304 345982
rect 41408 345920 42304 345980
rect 41408 345918 41414 345920
rect 42298 345918 42304 345920
rect 42368 345918 42374 345982
rect 42306 345728 42366 345918
rect 674938 345474 674944 345538
rect 675008 345536 675014 345538
rect 679887 345536 679953 345539
rect 675008 345534 679953 345536
rect 675008 345478 679892 345534
rect 679948 345478 679953 345534
rect 675008 345476 679953 345478
rect 675008 345474 675014 345476
rect 679887 345473 679953 345476
rect 40770 344354 40830 344914
rect 40762 344290 40768 344354
rect 40832 344290 40838 344354
rect 42735 344130 42801 344133
rect 42336 344128 42801 344130
rect 42336 344072 42740 344128
rect 42796 344072 42801 344128
rect 42336 344070 42801 344072
rect 42735 344067 42801 344070
rect 40962 342874 41022 343286
rect 40954 342810 40960 342874
rect 41024 342810 41030 342874
rect 42490 342662 42496 342726
rect 42560 342724 42566 342726
rect 43066 342724 43072 342726
rect 42560 342664 43072 342724
rect 42560 342662 42566 342664
rect 43066 342662 43072 342664
rect 43136 342662 43142 342726
rect 41346 341986 41406 342472
rect 41338 341922 41344 341986
rect 41408 341922 41414 341986
rect 41538 341246 41598 341806
rect 41530 341182 41536 341246
rect 41600 341182 41606 341246
rect 59535 340948 59601 340951
rect 654159 340948 654225 340951
rect 59535 340946 64416 340948
rect 37314 340359 37374 340918
rect 59535 340890 59540 340946
rect 59596 340890 64416 340946
rect 59535 340888 64416 340890
rect 650208 340946 654225 340948
rect 650208 340890 654164 340946
rect 654220 340890 654225 340946
rect 650208 340888 654225 340890
rect 59535 340885 59601 340888
rect 654159 340885 654225 340888
rect 37263 340354 37374 340359
rect 37263 340298 37268 340354
rect 37324 340298 37374 340354
rect 37263 340296 37374 340298
rect 37263 340293 37329 340296
rect 41154 339914 41214 340178
rect 41146 339850 41152 339914
rect 41216 339850 41222 339914
rect 40386 338730 40446 339290
rect 40378 338666 40384 338730
rect 40448 338666 40454 338730
rect 43407 338580 43473 338583
rect 42336 338578 43473 338580
rect 42336 338522 43412 338578
rect 43468 338522 43473 338578
rect 42336 338520 43473 338522
rect 43407 338517 43473 338520
rect 37122 337251 37182 337662
rect 37122 337246 37233 337251
rect 37359 337248 37425 337251
rect 37122 337190 37172 337246
rect 37228 337190 37233 337246
rect 37122 337188 37233 337190
rect 37167 337185 37233 337188
rect 37314 337246 37425 337248
rect 37314 337190 37364 337246
rect 37420 337190 37425 337246
rect 37314 337185 37425 337190
rect 37314 337070 37374 337185
rect 41922 335622 41982 336182
rect 41914 335558 41920 335622
rect 41984 335558 41990 335622
rect 43119 335472 43185 335475
rect 42336 335470 43185 335472
rect 42336 335414 43124 335470
rect 43180 335414 43185 335470
rect 42336 335412 43185 335414
rect 43119 335409 43185 335412
rect 675471 335178 675537 335179
rect 675471 335174 675520 335178
rect 675584 335176 675590 335178
rect 675471 335118 675476 335174
rect 675471 335114 675520 335118
rect 675584 335116 675628 335176
rect 675584 335114 675590 335116
rect 675471 335113 675537 335114
rect 43023 334584 43089 334587
rect 42336 334582 43089 334584
rect 42336 334526 43028 334582
rect 43084 334526 43089 334582
rect 42336 334524 43089 334526
rect 43023 334521 43089 334524
rect 42306 333403 42366 333814
rect 675322 333782 675328 333846
rect 675392 333844 675398 333846
rect 675471 333844 675537 333847
rect 675392 333842 675537 333844
rect 675392 333786 675476 333842
rect 675532 333786 675537 333842
rect 675392 333784 675537 333786
rect 675392 333782 675398 333784
rect 675471 333781 675537 333784
rect 674746 333486 674752 333550
rect 674816 333548 674822 333550
rect 675375 333548 675441 333551
rect 674816 333546 675441 333548
rect 674816 333490 675380 333546
rect 675436 333490 675441 333546
rect 674816 333488 675441 333490
rect 674816 333486 674822 333488
rect 675375 333485 675441 333488
rect 42306 333398 42417 333403
rect 42306 333342 42356 333398
rect 42412 333342 42417 333398
rect 42306 333340 42417 333342
rect 42351 333337 42417 333340
rect 42306 332071 42366 332260
rect 42306 332066 42417 332071
rect 42306 332010 42356 332066
rect 42412 332010 42417 332066
rect 42306 332008 42417 332010
rect 42351 332005 42417 332008
rect 675130 330526 675136 330590
rect 675200 330588 675206 330590
rect 675471 330588 675537 330591
rect 675200 330586 675537 330588
rect 675200 330530 675476 330586
rect 675532 330530 675537 330586
rect 675200 330528 675537 330530
rect 675200 330526 675206 330528
rect 675471 330525 675537 330528
rect 675183 329552 675249 329555
rect 675514 329552 675520 329554
rect 675183 329550 675520 329552
rect 675183 329494 675188 329550
rect 675244 329494 675520 329550
rect 675183 329492 675520 329494
rect 675183 329489 675249 329492
rect 675514 329490 675520 329492
rect 675584 329490 675590 329554
rect 653967 329256 654033 329259
rect 650208 329254 654033 329256
rect 650208 329198 653972 329254
rect 654028 329198 654033 329254
rect 650208 329196 654033 329198
rect 653967 329193 654033 329196
rect 674362 328306 674368 328370
rect 674432 328368 674438 328370
rect 675375 328368 675441 328371
rect 674432 328366 675441 328368
rect 674432 328310 675380 328366
rect 675436 328310 675441 328366
rect 674432 328308 675441 328310
rect 674432 328306 674438 328308
rect 675375 328305 675441 328308
rect 674554 326826 674560 326890
rect 674624 326888 674630 326890
rect 675375 326888 675441 326891
rect 674624 326886 675441 326888
rect 674624 326830 675380 326886
rect 675436 326830 675441 326886
rect 674624 326828 675441 326830
rect 674624 326826 674630 326828
rect 675375 326825 675441 326828
rect 59535 326444 59601 326447
rect 59535 326442 64416 326444
rect 59535 326386 59540 326442
rect 59596 326386 64416 326442
rect 59535 326384 64416 326386
rect 59535 326381 59601 326384
rect 674703 319932 674769 319935
rect 674703 319930 674814 319932
rect 674703 319874 674708 319930
rect 674764 319874 674814 319930
rect 674703 319869 674814 319874
rect 41530 319722 41536 319786
rect 41600 319784 41606 319786
rect 41775 319784 41841 319787
rect 41600 319782 41841 319784
rect 41600 319726 41780 319782
rect 41836 319726 41841 319782
rect 41600 319724 41841 319726
rect 41600 319722 41606 319724
rect 41775 319721 41841 319724
rect 674754 319680 674814 319869
rect 674415 318896 674481 318899
rect 674415 318894 674784 318896
rect 674415 318838 674420 318894
rect 674476 318838 674784 318894
rect 674415 318836 674784 318838
rect 674415 318833 674481 318836
rect 41530 318686 41536 318750
rect 41600 318748 41606 318750
rect 42159 318748 42225 318751
rect 43066 318748 43072 318750
rect 41600 318746 43072 318748
rect 41600 318690 42164 318746
rect 42220 318690 43072 318746
rect 41600 318688 43072 318690
rect 41600 318686 41606 318688
rect 42159 318685 42225 318688
rect 43066 318686 43072 318688
rect 43136 318686 43142 318750
rect 674703 318304 674769 318307
rect 674703 318302 674814 318304
rect 674703 318246 674708 318302
rect 674764 318246 674814 318302
rect 674703 318241 674814 318246
rect 674754 318052 674814 318241
rect 41775 318010 41841 318011
rect 41722 317946 41728 318010
rect 41792 318008 41841 318010
rect 41792 318006 41884 318008
rect 41836 317950 41884 318006
rect 41792 317948 41884 317950
rect 41792 317946 41841 317948
rect 41775 317945 41841 317946
rect 41871 317418 41937 317419
rect 41871 317416 41920 317418
rect 41828 317414 41920 317416
rect 41828 317358 41876 317414
rect 41828 317356 41920 317358
rect 41871 317354 41920 317356
rect 41984 317354 41990 317418
rect 655119 317416 655185 317419
rect 650208 317414 655185 317416
rect 650208 317358 655124 317414
rect 655180 317358 655185 317414
rect 650208 317356 655185 317358
rect 41871 317353 41937 317354
rect 655119 317353 655185 317356
rect 674170 317206 674176 317270
rect 674240 317268 674246 317270
rect 674240 317208 674784 317268
rect 674240 317206 674246 317208
rect 674170 316392 674176 316456
rect 674240 316454 674246 316456
rect 674240 316394 674784 316454
rect 674240 316392 674246 316394
rect 40378 316022 40384 316086
rect 40448 316084 40454 316086
rect 41775 316084 41841 316087
rect 40448 316082 41841 316084
rect 40448 316026 41780 316082
rect 41836 316026 41841 316082
rect 40448 316024 41841 316026
rect 40448 316022 40454 316024
rect 41775 316021 41841 316024
rect 674938 315874 674944 315938
rect 675008 315874 675014 315938
rect 674362 315726 674368 315790
rect 674432 315788 674438 315790
rect 674946 315788 675006 315874
rect 674432 315758 675006 315788
rect 674432 315728 674976 315758
rect 674432 315726 674438 315728
rect 41338 315578 41344 315642
rect 41408 315640 41414 315642
rect 41775 315640 41841 315643
rect 41408 315638 41841 315640
rect 41408 315582 41780 315638
rect 41836 315582 41841 315638
rect 41408 315580 41841 315582
rect 41408 315578 41414 315580
rect 41775 315577 41841 315580
rect 675898 315134 675904 315198
rect 675968 315134 675974 315198
rect 673978 314838 673984 314902
rect 674048 314900 674054 314902
rect 675906 314900 675966 315134
rect 674048 314870 675966 314900
rect 674048 314840 675936 314870
rect 674048 314838 674054 314840
rect 677058 313867 677118 314130
rect 41722 313802 41728 313866
rect 41792 313864 41798 313866
rect 43066 313864 43072 313866
rect 41792 313804 43072 313864
rect 41792 313802 41798 313804
rect 43066 313802 43072 313804
rect 43136 313802 43142 313866
rect 677007 313862 677118 313867
rect 677007 313806 677012 313862
rect 677068 313806 677118 313862
rect 677007 313804 677118 313806
rect 677007 313801 677073 313804
rect 40762 313654 40768 313718
rect 40832 313716 40838 313718
rect 41775 313716 41841 313719
rect 40832 313714 41841 313716
rect 40832 313658 41780 313714
rect 41836 313658 41841 313714
rect 40832 313656 41841 313658
rect 40832 313654 40838 313656
rect 41775 313653 41841 313656
rect 41146 313210 41152 313274
rect 41216 313272 41222 313274
rect 41775 313272 41841 313275
rect 41216 313270 41841 313272
rect 41216 313214 41780 313270
rect 41836 313214 41841 313270
rect 41216 313212 41841 313214
rect 41216 313210 41222 313212
rect 41775 313209 41841 313212
rect 674754 312682 674814 313242
rect 674746 312618 674752 312682
rect 674816 312618 674822 312682
rect 674319 312532 674385 312535
rect 674319 312530 674784 312532
rect 674319 312474 674324 312530
rect 674380 312474 674784 312530
rect 674319 312472 674784 312474
rect 674319 312469 674385 312472
rect 40954 312322 40960 312386
rect 41024 312384 41030 312386
rect 41775 312384 41841 312387
rect 41024 312382 41841 312384
rect 41024 312326 41780 312382
rect 41836 312326 41841 312382
rect 41024 312324 41841 312326
rect 41024 312322 41030 312324
rect 41775 312321 41841 312324
rect 59535 312236 59601 312239
rect 59535 312234 64416 312236
rect 59535 312178 59540 312234
rect 59596 312178 64416 312234
rect 59535 312176 64416 312178
rect 59535 312173 59601 312176
rect 676866 311499 676926 311614
rect 676866 311494 676977 311499
rect 676866 311438 676916 311494
rect 676972 311438 676977 311494
rect 676866 311436 676977 311438
rect 676911 311433 676977 311436
rect 676866 310759 676926 311022
rect 676815 310754 676926 310759
rect 676815 310698 676820 310754
rect 676876 310698 676926 310754
rect 676815 310696 676926 310698
rect 676815 310693 676881 310696
rect 674554 309510 674560 309574
rect 674624 309572 674630 309574
rect 674754 309572 674814 310134
rect 674624 309512 674814 309572
rect 674624 309510 674630 309512
rect 674607 309128 674673 309131
rect 674754 309128 674814 309394
rect 674607 309126 674814 309128
rect 674607 309070 674612 309126
rect 674668 309070 674814 309126
rect 674607 309068 674814 309070
rect 674607 309065 674673 309068
rect 674415 308536 674481 308539
rect 674415 308534 674784 308536
rect 674415 308478 674420 308534
rect 674476 308478 674784 308534
rect 674415 308476 674784 308478
rect 674415 308473 674481 308476
rect 675138 307503 675198 307766
rect 42255 307500 42321 307503
rect 42255 307498 42366 307500
rect 42255 307442 42260 307498
rect 42316 307442 42366 307498
rect 42255 307437 42366 307442
rect 675087 307498 675198 307503
rect 675087 307442 675092 307498
rect 675148 307442 675198 307498
rect 675087 307440 675198 307442
rect 675087 307437 675153 307440
rect 42306 307322 42366 307437
rect 42255 306760 42321 306763
rect 42255 306758 42366 306760
rect 42255 306702 42260 306758
rect 42316 306702 42366 306758
rect 42255 306697 42366 306702
rect 42306 306434 42366 306697
rect 674946 306466 675006 306878
rect 674938 306402 674944 306466
rect 675008 306402 675014 306466
rect 673935 306168 674001 306171
rect 674754 306168 674814 306212
rect 673935 306166 674814 306168
rect 673935 306110 673940 306166
rect 673996 306110 674814 306166
rect 673935 306108 674814 306110
rect 673935 306105 674001 306108
rect 42831 305724 42897 305727
rect 655215 305724 655281 305727
rect 42336 305722 42897 305724
rect 42336 305666 42836 305722
rect 42892 305666 42897 305722
rect 42336 305664 42897 305666
rect 650208 305722 655281 305724
rect 650208 305666 655220 305722
rect 655276 305666 655281 305722
rect 650208 305664 655281 305666
rect 42831 305661 42897 305664
rect 655215 305661 655281 305664
rect 674946 305283 675006 305398
rect 674946 305278 675057 305283
rect 674946 305222 674996 305278
rect 675052 305222 675057 305278
rect 674946 305220 675057 305222
rect 674991 305217 675057 305220
rect 43407 304836 43473 304839
rect 42336 304834 43473 304836
rect 42336 304778 43412 304834
rect 43468 304778 43473 304834
rect 42336 304776 43473 304778
rect 43407 304773 43473 304776
rect 674031 304540 674097 304543
rect 674754 304540 674814 304584
rect 674031 304538 674814 304540
rect 674031 304482 674036 304538
rect 674092 304482 674814 304538
rect 674031 304480 674814 304482
rect 674031 304477 674097 304480
rect 43215 304096 43281 304099
rect 42336 304094 43281 304096
rect 42336 304038 43220 304094
rect 43276 304038 43281 304094
rect 42336 304036 43281 304038
rect 43215 304033 43281 304036
rect 674223 303800 674289 303803
rect 674223 303798 674784 303800
rect 674223 303742 674228 303798
rect 674284 303742 674784 303798
rect 674223 303740 674784 303742
rect 674223 303737 674289 303740
rect 42114 302766 42174 303326
rect 40570 302702 40576 302766
rect 40640 302702 40646 302766
rect 42106 302702 42112 302766
rect 42176 302702 42182 302766
rect 42298 302702 42304 302766
rect 42368 302702 42374 302766
rect 40578 302616 40638 302702
rect 42306 302616 42366 302702
rect 40578 302556 42366 302616
rect 40578 302512 40638 302556
rect 679746 302471 679806 302956
rect 679746 302466 679857 302471
rect 679746 302410 679796 302466
rect 679852 302410 679857 302466
rect 679746 302408 679857 302410
rect 679791 302405 679857 302408
rect 679791 301728 679857 301731
rect 679746 301726 679857 301728
rect 40962 301138 41022 301698
rect 679746 301670 679796 301726
rect 679852 301670 679857 301726
rect 679746 301665 679857 301670
rect 679746 301402 679806 301665
rect 40954 301074 40960 301138
rect 41024 301074 41030 301138
rect 40002 300399 40062 300884
rect 39951 300394 40062 300399
rect 39951 300338 39956 300394
rect 40012 300338 40062 300394
rect 39951 300336 40062 300338
rect 39951 300333 40017 300336
rect 40770 299658 40830 300070
rect 40762 299594 40768 299658
rect 40832 299594 40838 299658
rect 41346 298770 41406 299256
rect 41338 298706 41344 298770
rect 41408 298706 41414 298770
rect 41530 298706 41536 298770
rect 41600 298768 41606 298770
rect 42490 298768 42496 298770
rect 41600 298708 42496 298768
rect 41600 298706 41606 298708
rect 42490 298706 42496 298708
rect 42560 298706 42566 298770
rect 41538 298030 41598 298590
rect 41530 297966 41536 298030
rect 41600 297966 41606 298030
rect 41730 297291 41790 297776
rect 59535 297732 59601 297735
rect 59535 297730 64416 297732
rect 59535 297674 59540 297730
rect 59596 297674 64416 297730
rect 59535 297672 64416 297674
rect 59535 297669 59601 297672
rect 41730 297286 41841 297291
rect 41730 297230 41780 297286
rect 41836 297230 41841 297286
rect 41730 297228 41841 297230
rect 41775 297225 41841 297228
rect 41154 296698 41214 296962
rect 41146 296634 41152 296698
rect 41216 296634 41222 296698
rect 40386 295514 40446 296074
rect 40378 295450 40384 295514
rect 40448 295450 40454 295514
rect 42114 294775 42174 295334
rect 42114 294770 42225 294775
rect 42114 294714 42164 294770
rect 42220 294714 42225 294770
rect 42114 294712 42225 294714
rect 42159 294709 42225 294712
rect 37314 294035 37374 294446
rect 37314 294030 37425 294035
rect 655407 294032 655473 294035
rect 37314 293974 37364 294030
rect 37420 293974 37425 294030
rect 37314 293972 37425 293974
rect 650208 294030 655473 294032
rect 650208 293974 655412 294030
rect 655468 293974 655473 294030
rect 650208 293972 655473 293974
rect 37359 293969 37425 293972
rect 655407 293969 655473 293972
rect 43119 293884 43185 293887
rect 42336 293882 43185 293884
rect 42336 293826 43124 293882
rect 43180 293826 43185 293882
rect 42336 293824 43185 293826
rect 43119 293821 43185 293824
rect 42306 292407 42366 292966
rect 42255 292402 42366 292407
rect 42255 292346 42260 292402
rect 42316 292346 42366 292402
rect 42255 292344 42366 292346
rect 42255 292341 42321 292344
rect 42831 292256 42897 292259
rect 42336 292254 42897 292256
rect 42336 292198 42836 292254
rect 42892 292198 42897 292254
rect 42336 292196 42897 292198
rect 42831 292193 42897 292196
rect 42306 290924 42366 291338
rect 42543 290924 42609 290927
rect 42306 290922 42609 290924
rect 42306 290866 42548 290922
rect 42604 290866 42609 290922
rect 42306 290864 42609 290866
rect 42543 290861 42609 290864
rect 43215 290628 43281 290631
rect 42336 290626 43281 290628
rect 42336 290570 43220 290626
rect 43276 290570 43281 290626
rect 42336 290568 43281 290570
rect 43215 290565 43281 290568
rect 675471 290186 675537 290187
rect 675471 290182 675520 290186
rect 675584 290184 675590 290186
rect 675471 290126 675476 290182
rect 675471 290122 675520 290126
rect 675584 290124 675628 290184
rect 675584 290122 675590 290124
rect 675471 290121 675537 290122
rect 675375 289594 675441 289595
rect 675322 289592 675328 289594
rect 675284 289532 675328 289592
rect 675392 289590 675441 289594
rect 675436 289534 675441 289590
rect 675322 289530 675328 289532
rect 675392 289530 675441 289534
rect 675375 289529 675441 289530
rect 42639 289148 42705 289151
rect 42336 289146 42705 289148
rect 42336 289090 42644 289146
rect 42700 289090 42705 289146
rect 42336 289088 42705 289090
rect 42639 289085 42705 289088
rect 674938 285238 674944 285302
rect 675008 285300 675014 285302
rect 675471 285300 675537 285303
rect 675008 285298 675537 285300
rect 675008 285242 675476 285298
rect 675532 285242 675537 285298
rect 675008 285240 675537 285242
rect 675008 285238 675014 285240
rect 675471 285237 675537 285240
rect 42255 283674 42321 283675
rect 42255 283670 42304 283674
rect 42368 283672 42374 283674
rect 42255 283614 42260 283670
rect 42255 283610 42304 283614
rect 42368 283612 42412 283672
rect 42368 283610 42374 283612
rect 674746 283610 674752 283674
rect 674816 283672 674822 283674
rect 675375 283672 675441 283675
rect 674816 283670 675441 283672
rect 674816 283614 675380 283670
rect 675436 283614 675441 283670
rect 674816 283612 675441 283614
rect 674816 283610 674822 283612
rect 42255 283609 42321 283610
rect 675375 283609 675441 283612
rect 57615 283524 57681 283527
rect 57615 283522 64416 283524
rect 57615 283466 57620 283522
rect 57676 283466 64416 283522
rect 57615 283464 64416 283466
rect 57615 283461 57681 283464
rect 41914 282278 41920 282342
rect 41984 282340 41990 282342
rect 42490 282340 42496 282342
rect 41984 282280 42496 282340
rect 41984 282278 41990 282280
rect 42490 282278 42496 282280
rect 42560 282278 42566 282342
rect 653775 282340 653841 282343
rect 650208 282338 653841 282340
rect 650208 282282 653780 282338
rect 653836 282282 653841 282338
rect 650208 282280 653841 282282
rect 653775 282277 653841 282280
rect 674746 282278 674752 282342
rect 674816 282340 674822 282342
rect 674991 282340 675057 282343
rect 674816 282338 675057 282340
rect 674816 282282 674996 282338
rect 675052 282282 675057 282338
rect 674816 282280 675057 282282
rect 674816 282278 674822 282280
rect 674991 282277 675057 282280
rect 674554 281834 674560 281898
rect 674624 281896 674630 281898
rect 675375 281896 675441 281899
rect 674624 281894 675441 281896
rect 674624 281838 675380 281894
rect 675436 281838 675441 281894
rect 674624 281836 675441 281838
rect 674624 281834 674630 281836
rect 675375 281833 675441 281836
rect 42298 281538 42304 281602
rect 42368 281600 42374 281602
rect 42639 281600 42705 281603
rect 42368 281598 42705 281600
rect 42368 281542 42644 281598
rect 42700 281542 42705 281598
rect 42368 281540 42705 281542
rect 42368 281538 42374 281540
rect 42639 281537 42705 281540
rect 41530 276506 41536 276570
rect 41600 276568 41606 276570
rect 41775 276568 41841 276571
rect 41600 276566 41841 276568
rect 41600 276510 41780 276566
rect 41836 276510 41841 276566
rect 41600 276508 41841 276510
rect 41600 276506 41606 276508
rect 41775 276505 41841 276508
rect 674703 274940 674769 274943
rect 674703 274938 674814 274940
rect 674703 274882 674708 274938
rect 674764 274882 674814 274938
rect 674703 274877 674814 274882
rect 41967 274794 42033 274795
rect 41914 274730 41920 274794
rect 41984 274792 42033 274794
rect 46479 274792 46545 274795
rect 41984 274790 46545 274792
rect 42028 274734 46484 274790
rect 46540 274734 46545 274790
rect 41984 274732 46545 274734
rect 41984 274730 42033 274732
rect 41967 274729 42033 274730
rect 46479 274729 46545 274732
rect 674754 274688 674814 274877
rect 675183 274348 675249 274351
rect 673794 274346 675249 274348
rect 673794 274290 675188 274346
rect 675244 274290 675249 274346
rect 673794 274288 675249 274290
rect 41722 273990 41728 274054
rect 41792 274052 41798 274054
rect 41967 274052 42033 274055
rect 43066 274052 43072 274054
rect 41792 274050 43072 274052
rect 41792 273994 41972 274050
rect 42028 273994 43072 274050
rect 41792 273992 43072 273994
rect 41792 273990 41798 273992
rect 41967 273989 42033 273992
rect 43066 273990 43072 273992
rect 43136 274052 43142 274054
rect 46287 274052 46353 274055
rect 43136 274050 46353 274052
rect 43136 273994 46292 274050
rect 46348 273994 46353 274050
rect 43136 273992 46353 273994
rect 43136 273990 43142 273992
rect 46287 273989 46353 273992
rect 46479 274052 46545 274055
rect 673794 274052 673854 274288
rect 675183 274285 675249 274288
rect 46479 274050 673854 274052
rect 46479 273994 46484 274050
rect 46540 273994 673854 274050
rect 46479 273992 673854 273994
rect 674703 274052 674769 274055
rect 674703 274050 674814 274052
rect 674703 273994 674708 274050
rect 674764 273994 674814 274050
rect 46479 273989 46545 273992
rect 674703 273989 674814 273994
rect 287866 273842 287872 273906
rect 287936 273904 287942 273906
rect 410703 273904 410769 273907
rect 287936 273902 410769 273904
rect 287936 273846 410708 273902
rect 410764 273846 410769 273902
rect 674754 273874 674814 273989
rect 287936 273844 410769 273846
rect 287936 273842 287942 273844
rect 410703 273841 410769 273844
rect 276399 273756 276465 273759
rect 282159 273756 282225 273759
rect 276399 273754 282225 273756
rect 276399 273698 276404 273754
rect 276460 273698 282164 273754
rect 282220 273698 282225 273754
rect 276399 273696 282225 273698
rect 276399 273693 276465 273696
rect 282159 273693 282225 273696
rect 299439 273756 299505 273759
rect 302319 273756 302385 273759
rect 319695 273756 319761 273759
rect 299439 273754 302385 273756
rect 299439 273698 299444 273754
rect 299500 273698 302324 273754
rect 302380 273698 302385 273754
rect 299439 273696 302385 273698
rect 299439 273693 299505 273696
rect 302319 273693 302385 273696
rect 302850 273754 319761 273756
rect 302850 273698 319700 273754
rect 319756 273698 319761 273754
rect 302850 273696 319761 273698
rect 247887 273608 247953 273611
rect 146754 273548 168510 273608
rect 100911 273460 100977 273463
rect 100674 273458 100977 273460
rect 100674 273402 100916 273458
rect 100972 273402 100977 273458
rect 100674 273400 100977 273402
rect 46287 273312 46353 273315
rect 66159 273312 66225 273315
rect 46287 273310 60414 273312
rect 46287 273254 46292 273310
rect 46348 273254 60414 273310
rect 46287 273252 60414 273254
rect 46287 273249 46353 273252
rect 60354 273238 60414 273252
rect 60546 273310 66225 273312
rect 60546 273254 66164 273310
rect 66220 273254 66225 273310
rect 60546 273252 66225 273254
rect 60546 273238 60606 273252
rect 66159 273249 66225 273252
rect 80559 273312 80625 273315
rect 86223 273312 86289 273315
rect 80559 273310 86289 273312
rect 80559 273254 80564 273310
rect 80620 273254 86228 273310
rect 86284 273254 86289 273310
rect 80559 273252 86289 273254
rect 80559 273249 80625 273252
rect 86223 273249 86289 273252
rect 86415 273312 86481 273315
rect 100674 273312 100734 273400
rect 100911 273397 100977 273400
rect 120783 273460 120849 273463
rect 146754 273460 146814 273548
rect 120783 273458 146814 273460
rect 120783 273402 120788 273458
rect 120844 273402 146814 273458
rect 120783 273400 146814 273402
rect 120783 273397 120849 273400
rect 86415 273310 100734 273312
rect 86415 273254 86420 273310
rect 86476 273254 100734 273310
rect 86415 273252 100734 273254
rect 86415 273249 86481 273252
rect 60354 273178 60606 273238
rect 168450 273164 168510 273548
rect 246210 273606 247953 273608
rect 246210 273550 247892 273606
rect 247948 273550 247953 273606
rect 246210 273548 247953 273550
rect 181551 273460 181617 273463
rect 207279 273460 207345 273463
rect 246210 273460 246270 273548
rect 247887 273545 247953 273548
rect 181551 273458 207345 273460
rect 181551 273402 181556 273458
rect 181612 273402 207284 273458
rect 207340 273402 207345 273458
rect 181551 273400 207345 273402
rect 181551 273397 181617 273400
rect 207279 273397 207345 273400
rect 227586 273400 246270 273460
rect 302319 273460 302385 273463
rect 302850 273460 302910 273696
rect 319695 273693 319761 273696
rect 443535 273756 443601 273759
rect 460623 273756 460689 273759
rect 443535 273754 460689 273756
rect 443535 273698 443540 273754
rect 443596 273698 460628 273754
rect 460684 273698 460689 273754
rect 443535 273696 460689 273698
rect 443535 273693 443601 273696
rect 460623 273693 460689 273696
rect 339759 273608 339825 273611
rect 403119 273608 403185 273611
rect 665199 273608 665265 273611
rect 674746 273608 674752 273610
rect 339759 273606 339966 273608
rect 339759 273550 339764 273606
rect 339820 273550 339966 273606
rect 339759 273548 339966 273550
rect 339759 273545 339825 273548
rect 302319 273458 302910 273460
rect 302319 273402 302324 273458
rect 302380 273402 302910 273458
rect 302319 273400 302910 273402
rect 339906 273460 339966 273548
rect 390210 273606 403185 273608
rect 390210 273550 403124 273606
rect 403180 273550 403185 273606
rect 390210 273548 403185 273550
rect 348399 273460 348465 273463
rect 339906 273458 348465 273460
rect 339906 273402 348404 273458
rect 348460 273402 348465 273458
rect 339906 273400 348465 273402
rect 208431 273312 208497 273315
rect 227586 273312 227646 273400
rect 302319 273397 302385 273400
rect 348399 273397 348465 273400
rect 348591 273460 348657 273463
rect 348591 273458 367230 273460
rect 348591 273402 348596 273458
rect 348652 273402 367230 273458
rect 348591 273400 367230 273402
rect 348591 273397 348657 273400
rect 208431 273310 227646 273312
rect 208431 273254 208436 273310
rect 208492 273254 227646 273310
rect 208431 273252 227646 273254
rect 247887 273312 247953 273315
rect 256335 273312 256401 273315
rect 247887 273310 256401 273312
rect 247887 273254 247892 273310
rect 247948 273254 256340 273310
rect 256396 273254 256401 273310
rect 247887 273252 256401 273254
rect 208431 273249 208497 273252
rect 247887 273249 247953 273252
rect 256335 273249 256401 273252
rect 181551 273164 181617 273167
rect 168450 273162 181617 273164
rect 168450 273106 181556 273162
rect 181612 273106 181617 273162
rect 168450 273104 181617 273106
rect 367170 273164 367230 273400
rect 390210 273312 390270 273548
rect 403119 273545 403185 273548
rect 508290 273548 509886 273608
rect 429231 273460 429297 273463
rect 437775 273460 437841 273463
rect 429231 273458 437841 273460
rect 429231 273402 429236 273458
rect 429292 273402 437780 273458
rect 437836 273402 437841 273458
rect 429231 273400 437841 273402
rect 429231 273397 429297 273400
rect 437775 273397 437841 273400
rect 460623 273460 460689 273463
rect 508290 273460 508350 273548
rect 460623 273458 508350 273460
rect 460623 273402 460628 273458
rect 460684 273402 508350 273458
rect 460623 273400 508350 273402
rect 509826 273460 509886 273548
rect 665199 273606 674752 273608
rect 665199 273550 665204 273606
rect 665260 273550 674752 273606
rect 665199 273548 674752 273550
rect 665199 273545 665265 273548
rect 674746 273546 674752 273548
rect 674816 273546 674822 273610
rect 674938 273546 674944 273610
rect 675008 273608 675014 273610
rect 675183 273608 675249 273611
rect 675008 273606 675249 273608
rect 675008 273550 675188 273606
rect 675244 273550 675249 273606
rect 675008 273548 675249 273550
rect 675008 273546 675014 273548
rect 675183 273545 675249 273548
rect 529839 273460 529905 273463
rect 509826 273458 529905 273460
rect 509826 273402 529844 273458
rect 529900 273402 529905 273458
rect 509826 273400 529905 273402
rect 460623 273397 460689 273400
rect 529839 273397 529905 273400
rect 550146 273400 570366 273460
rect 368706 273252 390270 273312
rect 410415 273312 410481 273315
rect 429039 273312 429105 273315
rect 410415 273310 429105 273312
rect 410415 273254 410420 273310
rect 410476 273254 429044 273310
rect 429100 273254 429105 273310
rect 410415 273252 429105 273254
rect 368706 273164 368766 273252
rect 410415 273249 410481 273252
rect 429039 273249 429105 273252
rect 530031 273312 530097 273315
rect 550146 273312 550206 273400
rect 530031 273310 550206 273312
rect 530031 273254 530036 273310
rect 530092 273254 550206 273310
rect 530031 273252 550206 273254
rect 570306 273312 570366 273400
rect 590466 273400 610686 273460
rect 590466 273312 590526 273400
rect 570306 273252 590526 273312
rect 610626 273312 610686 273400
rect 674703 273312 674769 273315
rect 610626 273252 630654 273312
rect 530031 273249 530097 273252
rect 367170 273104 368766 273164
rect 630594 273164 630654 273252
rect 674703 273310 674814 273312
rect 674703 273254 674708 273310
rect 674764 273254 674814 273310
rect 674703 273249 674814 273254
rect 645135 273164 645201 273167
rect 630594 273162 645201 273164
rect 630594 273106 645140 273162
rect 645196 273106 645201 273162
rect 630594 273104 645201 273106
rect 181551 273101 181617 273104
rect 645135 273101 645201 273104
rect 674754 273060 674814 273249
rect 40378 272806 40384 272870
rect 40448 272868 40454 272870
rect 41775 272868 41841 272871
rect 40448 272866 41841 272868
rect 40448 272810 41780 272866
rect 41836 272810 41841 272866
rect 40448 272808 41841 272810
rect 40448 272806 40454 272808
rect 41775 272805 41841 272808
rect 674799 272722 674865 272723
rect 674746 272720 674752 272722
rect 674708 272660 674752 272720
rect 674816 272718 674865 272722
rect 674860 272662 674865 272718
rect 674746 272658 674752 272660
rect 674816 272658 674865 272662
rect 674799 272657 674865 272658
rect 41338 272362 41344 272426
rect 41408 272424 41414 272426
rect 41775 272424 41841 272427
rect 41408 272422 41841 272424
rect 41408 272366 41780 272422
rect 41836 272366 41841 272422
rect 41408 272364 41841 272366
rect 41408 272362 41414 272364
rect 41775 272361 41841 272364
rect 674170 272214 674176 272278
rect 674240 272276 674246 272278
rect 674240 272216 674784 272276
rect 674240 272214 674246 272216
rect 675906 270946 675966 271432
rect 675898 270882 675904 270946
rect 675968 270882 675974 270946
rect 680079 270944 680145 270947
rect 680079 270942 680190 270944
rect 680079 270886 680084 270942
rect 680140 270886 680190 270942
rect 680079 270881 680190 270886
rect 674362 270734 674368 270798
rect 674432 270796 674438 270798
rect 680130 270796 680190 270881
rect 674432 270766 680190 270796
rect 674432 270736 680160 270766
rect 674432 270734 674438 270736
rect 40954 270586 40960 270650
rect 41024 270648 41030 270650
rect 41775 270648 41841 270651
rect 41024 270646 41841 270648
rect 41024 270590 41780 270646
rect 41836 270590 41841 270646
rect 41024 270588 41841 270590
rect 41024 270586 41030 270588
rect 41775 270585 41841 270588
rect 100239 270648 100305 270651
rect 430287 270648 430353 270651
rect 100239 270646 430353 270648
rect 100239 270590 100244 270646
rect 100300 270590 430292 270646
rect 430348 270590 430353 270646
rect 100239 270588 430353 270590
rect 100239 270585 100305 270588
rect 430287 270585 430353 270588
rect 442234 270586 442240 270650
rect 442304 270648 442310 270650
rect 444015 270648 444081 270651
rect 442304 270646 444081 270648
rect 442304 270590 444020 270646
rect 444076 270590 444081 270646
rect 442304 270588 444081 270590
rect 442304 270586 442310 270588
rect 444015 270585 444081 270588
rect 449967 270648 450033 270651
rect 450682 270648 450688 270650
rect 449967 270646 450688 270648
rect 449967 270590 449972 270646
rect 450028 270590 450688 270646
rect 449967 270588 450688 270590
rect 449967 270585 450033 270588
rect 450682 270586 450688 270588
rect 450752 270586 450758 270650
rect 95535 270500 95601 270503
rect 426351 270500 426417 270503
rect 95535 270498 426417 270500
rect 95535 270442 95540 270498
rect 95596 270442 426356 270498
rect 426412 270442 426417 270498
rect 95535 270440 426417 270442
rect 95535 270437 95601 270440
rect 426351 270437 426417 270440
rect 442863 270500 442929 270503
rect 446458 270500 446464 270502
rect 442863 270498 446464 270500
rect 442863 270442 442868 270498
rect 442924 270442 446464 270498
rect 442863 270440 446464 270442
rect 442863 270437 442929 270440
rect 446458 270438 446464 270440
rect 446528 270438 446534 270502
rect 449530 270438 449536 270502
rect 449600 270500 449606 270502
rect 451119 270500 451185 270503
rect 449600 270498 451185 270500
rect 449600 270442 451124 270498
rect 451180 270442 451185 270498
rect 449600 270440 451185 270442
rect 449600 270438 449606 270440
rect 451119 270437 451185 270440
rect 93135 270352 93201 270355
rect 430095 270352 430161 270355
rect 93135 270350 430161 270352
rect 93135 270294 93140 270350
rect 93196 270294 430100 270350
rect 430156 270294 430161 270350
rect 93135 270292 430161 270294
rect 93135 270289 93201 270292
rect 430095 270289 430161 270292
rect 439311 270352 439377 270355
rect 443578 270352 443584 270354
rect 439311 270350 443584 270352
rect 439311 270294 439316 270350
rect 439372 270294 443584 270350
rect 439311 270292 443584 270294
rect 439311 270289 439377 270292
rect 443578 270290 443584 270292
rect 443648 270290 443654 270354
rect 90735 270204 90801 270207
rect 432207 270204 432273 270207
rect 443002 270204 443008 270206
rect 90735 270202 430974 270204
rect 90735 270146 90740 270202
rect 90796 270146 430974 270202
rect 90735 270144 430974 270146
rect 90735 270141 90801 270144
rect 41146 269994 41152 270058
rect 41216 270056 41222 270058
rect 41775 270056 41841 270059
rect 41216 270054 41841 270056
rect 41216 269998 41780 270054
rect 41836 269998 41841 270054
rect 41216 269996 41841 269998
rect 41216 269994 41222 269996
rect 41775 269993 41841 269996
rect 83631 270056 83697 270059
rect 428463 270056 428529 270059
rect 83631 270054 428529 270056
rect 83631 269998 83636 270054
rect 83692 269998 428468 270054
rect 428524 269998 428529 270054
rect 83631 269996 428529 269998
rect 430914 270056 430974 270144
rect 432207 270202 443008 270204
rect 432207 270146 432212 270202
rect 432268 270146 443008 270202
rect 432207 270144 443008 270146
rect 432207 270141 432273 270144
rect 443002 270142 443008 270144
rect 443072 270142 443078 270206
rect 472527 270204 472593 270207
rect 443202 270202 472593 270204
rect 443202 270146 472532 270202
rect 472588 270146 472593 270202
rect 443202 270144 472593 270146
rect 432783 270056 432849 270059
rect 430914 270054 432849 270056
rect 430914 269998 432788 270054
rect 432844 269998 432849 270054
rect 430914 269996 432849 269998
rect 83631 269993 83697 269996
rect 428463 269993 428529 269996
rect 432783 269993 432849 269996
rect 442042 269994 442048 270058
rect 442112 270056 442118 270058
rect 443202 270056 443262 270144
rect 472527 270141 472593 270144
rect 442112 269996 443262 270056
rect 442112 269994 442118 269996
rect 77679 269908 77745 269911
rect 423567 269908 423633 269911
rect 77679 269906 423633 269908
rect 77679 269850 77684 269906
rect 77740 269850 423572 269906
rect 423628 269850 423633 269906
rect 77679 269848 423633 269850
rect 77679 269845 77745 269848
rect 423567 269845 423633 269848
rect 673978 269846 673984 269910
rect 674048 269908 674054 269910
rect 674048 269848 674784 269908
rect 674048 269846 674054 269848
rect 69327 269760 69393 269763
rect 425871 269760 425937 269763
rect 69327 269758 425937 269760
rect 69327 269702 69332 269758
rect 69388 269702 425876 269758
rect 425932 269702 425937 269758
rect 69327 269700 425937 269702
rect 69327 269697 69393 269700
rect 425871 269697 425937 269700
rect 433263 269760 433329 269763
rect 449722 269760 449728 269762
rect 433263 269758 449728 269760
rect 433263 269702 433268 269758
rect 433324 269702 449728 269758
rect 433263 269700 449728 269702
rect 433263 269697 433329 269700
rect 449722 269698 449728 269700
rect 449792 269698 449798 269762
rect 81327 269612 81393 269615
rect 437199 269612 437265 269615
rect 81327 269610 437265 269612
rect 81327 269554 81332 269610
rect 81388 269554 437204 269610
rect 437260 269554 437265 269610
rect 81327 269552 437265 269554
rect 81327 269549 81393 269552
rect 437199 269549 437265 269552
rect 71727 269464 71793 269467
rect 433455 269464 433521 269467
rect 71727 269462 433521 269464
rect 71727 269406 71732 269462
rect 71788 269406 433460 269462
rect 433516 269406 433521 269462
rect 71727 269404 433521 269406
rect 71727 269401 71793 269404
rect 433455 269401 433521 269404
rect 445690 269402 445696 269466
rect 445760 269464 445766 269466
rect 465519 269464 465585 269467
rect 445760 269462 465585 269464
rect 445760 269406 465524 269462
rect 465580 269406 465585 269462
rect 445760 269404 465585 269406
rect 445760 269402 445766 269404
rect 465519 269401 465585 269404
rect 66927 269316 66993 269319
rect 431151 269316 431217 269319
rect 452218 269316 452224 269318
rect 66927 269314 431217 269316
rect 66927 269258 66932 269314
rect 66988 269258 431156 269314
rect 431212 269258 431217 269314
rect 66927 269256 431217 269258
rect 66927 269253 66993 269256
rect 431151 269253 431217 269256
rect 447426 269256 452224 269316
rect 40762 269106 40768 269170
rect 40832 269168 40838 269170
rect 41775 269168 41841 269171
rect 40832 269166 41841 269168
rect 40832 269110 41780 269166
rect 41836 269110 41841 269166
rect 40832 269108 41841 269110
rect 40832 269106 40838 269108
rect 41775 269105 41841 269108
rect 107439 269168 107505 269171
rect 435951 269168 436017 269171
rect 107439 269166 436017 269168
rect 107439 269110 107444 269166
rect 107500 269110 435956 269166
rect 436012 269110 436017 269166
rect 107439 269108 436017 269110
rect 107439 269105 107505 269108
rect 435951 269105 436017 269108
rect 290362 268958 290368 269022
rect 290432 269020 290438 269022
rect 423759 269020 423825 269023
rect 290432 269018 423825 269020
rect 290432 268962 423764 269018
rect 423820 268962 423825 269018
rect 290432 268960 423825 268962
rect 290432 268958 290438 268960
rect 423759 268957 423825 268960
rect 426159 269020 426225 269023
rect 447226 269020 447232 269022
rect 426159 269018 447232 269020
rect 426159 268962 426164 269018
rect 426220 268962 447232 269018
rect 426159 268960 447232 268962
rect 426159 268957 426225 268960
rect 447226 268958 447232 268960
rect 447296 268958 447302 269022
rect 290170 268810 290176 268874
rect 290240 268872 290246 268874
rect 416655 268872 416721 268875
rect 290240 268870 416721 268872
rect 290240 268814 416660 268870
rect 416716 268814 416721 268870
rect 290240 268812 416721 268814
rect 290240 268810 290246 268812
rect 416655 268809 416721 268812
rect 419343 268872 419409 268875
rect 447426 268872 447486 269256
rect 452218 269254 452224 269256
rect 452288 269254 452294 269318
rect 452410 269168 452416 269170
rect 419343 268870 447486 268872
rect 419343 268814 419348 268870
rect 419404 268814 447486 268870
rect 419343 268812 447486 268814
rect 447618 269108 452416 269168
rect 419343 268809 419409 268812
rect 290746 268662 290752 268726
rect 290816 268724 290822 268726
rect 409551 268724 409617 268727
rect 290816 268722 409617 268724
rect 290816 268666 409556 268722
rect 409612 268666 409617 268722
rect 290816 268664 409617 268666
rect 290816 268662 290822 268664
rect 409551 268661 409617 268664
rect 290554 268514 290560 268578
rect 290624 268576 290630 268578
rect 398895 268576 398961 268579
rect 290624 268574 398961 268576
rect 290624 268518 398900 268574
rect 398956 268518 398961 268574
rect 290624 268516 398961 268518
rect 290624 268514 290630 268516
rect 398895 268513 398961 268516
rect 401199 268576 401265 268579
rect 447618 268576 447678 269108
rect 452410 269106 452416 269108
rect 452480 269106 452486 269170
rect 469359 269168 469425 269171
rect 480879 269168 480945 269171
rect 469359 269166 480945 269168
rect 469359 269110 469364 269166
rect 469420 269110 480884 269166
rect 480940 269110 480945 269166
rect 469359 269108 480945 269110
rect 469359 269105 469425 269108
rect 480879 269105 480945 269108
rect 674754 268578 674814 269138
rect 401199 268574 447678 268576
rect 401199 268518 401204 268574
rect 401260 268518 447678 268574
rect 401199 268516 447678 268518
rect 401199 268513 401265 268516
rect 674746 268514 674752 268578
rect 674816 268514 674822 268578
rect 425007 268428 425073 268431
rect 437871 268428 437937 268431
rect 425007 268426 437937 268428
rect 425007 268370 425012 268426
rect 425068 268370 437876 268426
rect 437932 268370 437937 268426
rect 425007 268368 437937 268370
rect 425007 268365 425073 268368
rect 437871 268365 437937 268368
rect 440463 268428 440529 268431
rect 449338 268428 449344 268430
rect 440463 268426 449344 268428
rect 440463 268370 440468 268426
rect 440524 268370 449344 268426
rect 440463 268368 449344 268370
rect 440463 268365 440529 268368
rect 449338 268366 449344 268368
rect 449408 268366 449414 268430
rect 417807 268280 417873 268283
rect 443386 268280 443392 268282
rect 417807 268278 443392 268280
rect 417807 268222 417812 268278
rect 417868 268222 443392 268278
rect 417807 268220 443392 268222
rect 417807 268217 417873 268220
rect 443386 268218 443392 268220
rect 443456 268218 443462 268282
rect 344559 268132 344625 268135
rect 348207 268132 348273 268135
rect 344559 268130 348273 268132
rect 344559 268074 344564 268130
rect 344620 268074 348212 268130
rect 348268 268074 348273 268130
rect 344559 268072 348273 268074
rect 344559 268069 344625 268072
rect 348207 268069 348273 268072
rect 380175 268132 380241 268135
rect 398127 268132 398193 268135
rect 380175 268130 398193 268132
rect 380175 268074 380180 268130
rect 380236 268074 398132 268130
rect 398188 268074 398193 268130
rect 380175 268072 398193 268074
rect 380175 268069 380241 268072
rect 398127 268069 398193 268072
rect 437871 268132 437937 268135
rect 675714 268134 675774 268250
rect 446650 268132 446656 268134
rect 437871 268130 446656 268132
rect 437871 268074 437876 268130
rect 437932 268074 446656 268130
rect 437871 268072 446656 268074
rect 437871 268069 437937 268072
rect 446650 268070 446656 268072
rect 446720 268070 446726 268134
rect 675706 268070 675712 268134
rect 675776 268070 675782 268134
rect 322671 267984 322737 267987
rect 339759 267984 339825 267987
rect 322671 267982 339825 267984
rect 322671 267926 322676 267982
rect 322732 267926 339764 267982
rect 339820 267926 339825 267982
rect 322671 267924 339825 267926
rect 322671 267921 322737 267924
rect 339759 267921 339825 267924
rect 284794 267774 284800 267838
rect 284864 267836 284870 267838
rect 434895 267836 434961 267839
rect 284864 267834 434961 267836
rect 284864 267778 434900 267834
rect 434956 267778 434961 267834
rect 284864 267776 434961 267778
rect 284864 267774 284870 267776
rect 434895 267773 434961 267776
rect 289978 267626 289984 267690
rect 290048 267688 290054 267690
rect 448815 267688 448881 267691
rect 290048 267686 448881 267688
rect 290048 267630 448820 267686
rect 448876 267630 448881 267686
rect 290048 267628 448881 267630
rect 290048 267626 290054 267628
rect 448815 267625 448881 267628
rect 284410 267478 284416 267542
rect 284480 267540 284486 267542
rect 459087 267540 459153 267543
rect 284480 267538 459153 267540
rect 284480 267482 459092 267538
rect 459148 267482 459153 267538
rect 284480 267480 459153 267482
rect 284480 267478 284486 267480
rect 459087 267477 459153 267480
rect 292858 267330 292864 267394
rect 292928 267392 292934 267394
rect 470127 267392 470193 267395
rect 292928 267390 470193 267392
rect 292928 267334 470132 267390
rect 470188 267334 470193 267390
rect 292928 267332 470193 267334
rect 292928 267330 292934 267332
rect 470127 267329 470193 267332
rect 675330 267247 675390 267510
rect 289210 267182 289216 267246
rect 289280 267244 289286 267246
rect 480975 267244 481041 267247
rect 289280 267242 481041 267244
rect 289280 267186 480980 267242
rect 481036 267186 481041 267242
rect 289280 267184 481041 267186
rect 289280 267182 289286 267184
rect 480975 267181 481041 267184
rect 538479 267244 538545 267247
rect 561519 267244 561585 267247
rect 538479 267242 561585 267244
rect 538479 267186 538484 267242
rect 538540 267186 561524 267242
rect 561580 267186 561585 267242
rect 538479 267184 561585 267186
rect 675330 267242 675441 267247
rect 675330 267186 675380 267242
rect 675436 267186 675441 267242
rect 675330 267184 675441 267186
rect 538479 267181 538545 267184
rect 561519 267181 561585 267184
rect 675375 267181 675441 267184
rect 289551 267096 289617 267099
rect 559407 267096 559473 267099
rect 289551 267094 559473 267096
rect 289551 267038 289556 267094
rect 289612 267038 559412 267094
rect 559468 267038 559473 267094
rect 289551 267036 559473 267038
rect 289551 267033 289617 267036
rect 559407 267033 559473 267036
rect 289935 266948 290001 266951
rect 562959 266948 563025 266951
rect 289935 266946 563025 266948
rect 289935 266890 289940 266946
rect 289996 266890 562964 266946
rect 563020 266890 563025 266946
rect 289935 266888 563025 266890
rect 289935 266885 290001 266888
rect 562959 266885 563025 266888
rect 283695 266800 283761 266803
rect 555855 266800 555921 266803
rect 283695 266798 555921 266800
rect 283695 266742 283700 266798
rect 283756 266742 555860 266798
rect 555916 266742 555921 266798
rect 283695 266740 555921 266742
rect 283695 266737 283761 266740
rect 555855 266737 555921 266740
rect 590223 266800 590289 266803
rect 590511 266800 590577 266803
rect 590223 266798 590577 266800
rect 590223 266742 590228 266798
rect 590284 266742 590516 266798
rect 590572 266742 590577 266798
rect 590223 266740 590577 266742
rect 590223 266737 590289 266740
rect 590511 266737 590577 266740
rect 610383 266800 610449 266803
rect 610671 266800 610737 266803
rect 610383 266798 610737 266800
rect 610383 266742 610388 266798
rect 610444 266742 610676 266798
rect 610732 266742 610737 266798
rect 610383 266740 610737 266742
rect 610383 266737 610449 266740
rect 610671 266737 610737 266740
rect 290319 266652 290385 266655
rect 570063 266652 570129 266655
rect 290319 266650 570129 266652
rect 290319 266594 290324 266650
rect 290380 266594 570068 266650
rect 570124 266594 570129 266650
rect 290319 266592 570129 266594
rect 290319 266589 290385 266592
rect 570063 266589 570129 266592
rect 590127 266652 590193 266655
rect 590607 266652 590673 266655
rect 590127 266650 590673 266652
rect 590127 266594 590132 266650
rect 590188 266594 590612 266650
rect 590668 266594 590673 266650
rect 590127 266592 590673 266594
rect 590127 266589 590193 266592
rect 590607 266589 590673 266592
rect 676866 266507 676926 266622
rect 283791 266504 283857 266507
rect 573711 266504 573777 266507
rect 283791 266502 573777 266504
rect 283791 266446 283796 266502
rect 283852 266446 573716 266502
rect 573772 266446 573777 266502
rect 283791 266444 573777 266446
rect 283791 266441 283857 266444
rect 573711 266441 573777 266444
rect 676815 266502 676926 266507
rect 676815 266446 676820 266502
rect 676876 266446 676926 266502
rect 676815 266444 676926 266446
rect 676815 266441 676881 266444
rect 283887 266356 283953 266359
rect 587919 266356 587985 266359
rect 283887 266354 587985 266356
rect 283887 266298 283892 266354
rect 283948 266298 587924 266354
rect 587980 266298 587985 266354
rect 283887 266296 587985 266298
rect 283887 266293 283953 266296
rect 587919 266293 587985 266296
rect 284986 266146 284992 266210
rect 285056 266208 285062 266210
rect 432015 266208 432081 266211
rect 285056 266206 432081 266208
rect 285056 266150 432020 266206
rect 432076 266150 432081 266206
rect 285056 266148 432081 266150
rect 285056 266146 285062 266148
rect 432015 266145 432081 266148
rect 284026 265998 284032 266062
rect 284096 266060 284102 266062
rect 429135 266060 429201 266063
rect 284096 266058 429201 266060
rect 284096 266002 429140 266058
rect 429196 266002 429201 266058
rect 284096 266000 429201 266002
rect 284096 265998 284102 266000
rect 429135 265997 429201 266000
rect 290703 265912 290769 265915
rect 432303 265912 432369 265915
rect 290703 265910 432369 265912
rect 290703 265854 290708 265910
rect 290764 265854 432308 265910
rect 432364 265854 432369 265910
rect 290703 265852 432369 265854
rect 290703 265849 290769 265852
rect 432303 265849 432369 265852
rect 291087 265764 291153 265767
rect 432111 265764 432177 265767
rect 291087 265762 432177 265764
rect 291087 265706 291092 265762
rect 291148 265706 432116 265762
rect 432172 265706 432177 265762
rect 291087 265704 432177 265706
rect 291087 265701 291153 265704
rect 432111 265701 432177 265704
rect 383439 265616 383505 265619
rect 389775 265616 389841 265619
rect 383439 265614 389841 265616
rect 383439 265558 383444 265614
rect 383500 265558 389780 265614
rect 389836 265558 389841 265614
rect 383439 265556 389841 265558
rect 383439 265553 383505 265556
rect 389775 265553 389841 265556
rect 382191 265468 382257 265471
rect 385647 265468 385713 265471
rect 382191 265466 385713 265468
rect 382191 265410 382196 265466
rect 382252 265410 385652 265466
rect 385708 265410 385713 265466
rect 382191 265408 385713 265410
rect 382191 265405 382257 265408
rect 385647 265405 385713 265408
rect 674554 265406 674560 265470
rect 674624 265468 674630 265470
rect 674754 265468 674814 266030
rect 674624 265408 674814 265468
rect 674624 265406 674630 265408
rect 674362 265110 674368 265174
rect 674432 265172 674438 265174
rect 674432 265112 674784 265172
rect 674432 265110 674438 265112
rect 329199 265024 329265 265027
rect 338703 265024 338769 265027
rect 329199 265022 338769 265024
rect 329199 264966 329204 265022
rect 329260 264966 338708 265022
rect 338764 264966 338769 265022
rect 329199 264964 338769 264966
rect 329199 264961 329265 264964
rect 338703 264961 338769 264964
rect 42106 264814 42112 264878
rect 42176 264876 42182 264878
rect 43311 264876 43377 264879
rect 42176 264874 43377 264876
rect 42176 264818 43316 264874
rect 43372 264818 43377 264874
rect 42176 264816 43377 264818
rect 42176 264814 42182 264816
rect 43311 264813 43377 264816
rect 287674 264814 287680 264878
rect 287744 264876 287750 264878
rect 455919 264876 455985 264879
rect 287744 264874 455985 264876
rect 287744 264818 455924 264874
rect 455980 264818 455985 264874
rect 287744 264816 455985 264818
rect 287744 264814 287750 264816
rect 455919 264813 455985 264816
rect 197871 264728 197937 264731
rect 387471 264728 387537 264731
rect 197871 264726 387537 264728
rect 197871 264670 197876 264726
rect 197932 264670 387476 264726
rect 387532 264670 387537 264726
rect 197871 264668 387537 264670
rect 197871 264665 197937 264668
rect 387471 264665 387537 264668
rect 332655 264580 332721 264583
rect 607023 264580 607089 264583
rect 332655 264578 607089 264580
rect 332655 264522 332660 264578
rect 332716 264522 607028 264578
rect 607084 264522 607089 264578
rect 332655 264520 607089 264522
rect 332655 264517 332721 264520
rect 607023 264517 607089 264520
rect 312399 264432 312465 264435
rect 318639 264432 318705 264435
rect 312399 264430 318705 264432
rect 312399 264374 312404 264430
rect 312460 264374 318644 264430
rect 318700 264374 318705 264430
rect 312399 264372 318705 264374
rect 312399 264369 312465 264372
rect 318639 264369 318705 264372
rect 333039 264432 333105 264435
rect 610575 264432 610641 264435
rect 333039 264430 610641 264432
rect 333039 264374 333044 264430
rect 333100 264374 610580 264430
rect 610636 264374 610641 264430
rect 333039 264372 610641 264374
rect 333039 264369 333105 264372
rect 610575 264369 610641 264372
rect 42255 264284 42321 264287
rect 333423 264284 333489 264287
rect 614127 264284 614193 264287
rect 42255 264282 42366 264284
rect 42255 264226 42260 264282
rect 42316 264226 42366 264282
rect 42255 264221 42366 264226
rect 333423 264282 614193 264284
rect 333423 264226 333428 264282
rect 333484 264226 614132 264282
rect 614188 264226 614193 264282
rect 333423 264224 614193 264226
rect 333423 264221 333489 264224
rect 614127 264221 614193 264224
rect 42306 264106 42366 264221
rect 675330 264139 675390 264402
rect 333711 264136 333777 264139
rect 617679 264136 617745 264139
rect 333711 264134 617745 264136
rect 333711 264078 333716 264134
rect 333772 264078 617684 264134
rect 617740 264078 617745 264134
rect 333711 264076 617745 264078
rect 333711 264073 333777 264076
rect 617679 264073 617745 264076
rect 675279 264134 675390 264139
rect 675279 264078 675284 264134
rect 675340 264078 675390 264134
rect 675279 264076 675390 264078
rect 675279 264073 675345 264076
rect 120495 263988 120561 263991
rect 330735 263988 330801 263991
rect 120495 263986 330801 263988
rect 120495 263930 120500 263986
rect 120556 263930 330740 263986
rect 330796 263930 330801 263986
rect 120495 263928 330801 263930
rect 120495 263925 120561 263928
rect 330735 263925 330801 263928
rect 335631 263988 335697 263991
rect 631983 263988 632049 263991
rect 335631 263986 632049 263988
rect 335631 263930 335636 263986
rect 335692 263930 631988 263986
rect 632044 263930 632049 263986
rect 335631 263928 632049 263930
rect 335631 263925 335697 263928
rect 631983 263925 632049 263928
rect 116943 263840 117009 263843
rect 331119 263840 331185 263843
rect 116943 263838 331185 263840
rect 116943 263782 116948 263838
rect 117004 263782 331124 263838
rect 331180 263782 331185 263838
rect 116943 263780 331185 263782
rect 116943 263777 117009 263780
rect 331119 263777 331185 263780
rect 335919 263840 335985 263843
rect 635535 263840 635601 263843
rect 335919 263838 635601 263840
rect 335919 263782 335924 263838
rect 335980 263782 635540 263838
rect 635596 263782 635601 263838
rect 335919 263780 635601 263782
rect 335919 263777 335985 263780
rect 635535 263777 635601 263780
rect 113391 263692 113457 263695
rect 330927 263692 330993 263695
rect 113391 263690 330993 263692
rect 113391 263634 113396 263690
rect 113452 263634 330932 263690
rect 330988 263634 330993 263690
rect 113391 263632 330993 263634
rect 113391 263629 113457 263632
rect 330927 263629 330993 263632
rect 336303 263692 336369 263695
rect 639087 263692 639153 263695
rect 336303 263690 639153 263692
rect 336303 263634 336308 263690
rect 336364 263634 639092 263690
rect 639148 263634 639153 263690
rect 336303 263632 639153 263634
rect 336303 263629 336369 263632
rect 639087 263629 639153 263632
rect 42255 263544 42321 263547
rect 72975 263544 73041 263547
rect 333999 263544 334065 263547
rect 42255 263542 42366 263544
rect 42255 263486 42260 263542
rect 42316 263486 42366 263542
rect 42255 263481 42366 263486
rect 72975 263542 334065 263544
rect 72975 263486 72980 263542
rect 73036 263486 334004 263542
rect 334060 263486 334065 263542
rect 72975 263484 334065 263486
rect 72975 263481 73041 263484
rect 333999 263481 334065 263484
rect 336687 263544 336753 263547
rect 642639 263544 642705 263547
rect 336687 263542 642705 263544
rect 336687 263486 336692 263542
rect 336748 263486 642644 263542
rect 642700 263486 642705 263542
rect 336687 263484 642705 263486
rect 336687 263481 336753 263484
rect 642639 263481 642705 263484
rect 42306 263218 42366 263481
rect 675138 263399 675198 263514
rect 289018 263334 289024 263398
rect 289088 263396 289094 263398
rect 441615 263396 441681 263399
rect 289088 263394 441681 263396
rect 289088 263338 441620 263394
rect 441676 263338 441681 263394
rect 289088 263336 441681 263338
rect 675138 263394 675249 263399
rect 675138 263338 675188 263394
rect 675244 263338 675249 263394
rect 675138 263336 675249 263338
rect 289088 263334 289094 263336
rect 441615 263333 441681 263336
rect 675183 263333 675249 263336
rect 237039 263248 237105 263251
rect 384495 263248 384561 263251
rect 237039 263246 384561 263248
rect 237039 263190 237044 263246
rect 237100 263190 384500 263246
rect 384556 263190 384561 263246
rect 237039 263188 384561 263190
rect 237039 263185 237105 263188
rect 384495 263185 384561 263188
rect 291514 263038 291520 263102
rect 291584 263100 291590 263102
rect 438063 263100 438129 263103
rect 291584 263098 438129 263100
rect 291584 263042 438068 263098
rect 438124 263042 438129 263098
rect 291584 263040 438129 263042
rect 291584 263038 291590 263040
rect 438063 263037 438129 263040
rect 289786 262890 289792 262954
rect 289856 262952 289862 262954
rect 430959 262952 431025 262955
rect 289856 262950 431025 262952
rect 289856 262894 430964 262950
rect 431020 262894 431025 262950
rect 289856 262892 431025 262894
rect 289856 262890 289862 262892
rect 430959 262889 431025 262892
rect 330831 262804 330897 262807
rect 427215 262804 427281 262807
rect 330831 262802 427281 262804
rect 330831 262746 330836 262802
rect 330892 262746 427220 262802
rect 427276 262746 427281 262802
rect 330831 262744 427281 262746
rect 330831 262741 330897 262744
rect 427215 262741 427281 262744
rect 674415 262804 674481 262807
rect 674415 262802 674784 262804
rect 674415 262746 674420 262802
rect 674476 262746 674784 262802
rect 674415 262744 674784 262746
rect 674415 262741 674481 262744
rect 330447 262656 330513 262659
rect 427119 262656 427185 262659
rect 330447 262654 427185 262656
rect 330447 262598 330452 262654
rect 330508 262598 427124 262654
rect 427180 262598 427185 262654
rect 330447 262596 427185 262598
rect 330447 262593 330513 262596
rect 427119 262593 427185 262596
rect 42831 262508 42897 262511
rect 42336 262506 42897 262508
rect 42336 262450 42836 262506
rect 42892 262450 42897 262506
rect 42336 262448 42897 262450
rect 42831 262445 42897 262448
rect 332271 262508 332337 262511
rect 429711 262508 429777 262511
rect 332271 262506 429777 262508
rect 332271 262450 332276 262506
rect 332332 262450 429716 262506
rect 429772 262450 429777 262506
rect 332271 262448 429777 262450
rect 332271 262445 332337 262448
rect 429711 262445 429777 262448
rect 287482 262150 287488 262214
rect 287552 262212 287558 262214
rect 514959 262212 515025 262215
rect 287552 262210 515025 262212
rect 287552 262154 514964 262210
rect 515020 262154 515025 262210
rect 287552 262152 515025 262154
rect 287552 262150 287558 262152
rect 514959 262149 515025 262152
rect 674799 262212 674865 262215
rect 675322 262212 675328 262214
rect 674799 262210 675328 262212
rect 674799 262154 674804 262210
rect 674860 262154 675328 262210
rect 674799 262152 675328 262154
rect 674799 262149 674865 262152
rect 675322 262150 675328 262152
rect 675392 262150 675398 262214
rect 291471 262064 291537 262067
rect 584367 262064 584433 262067
rect 291471 262062 584433 262064
rect 291471 262006 291476 262062
rect 291532 262006 584372 262062
rect 584428 262006 584433 262062
rect 291471 262004 584433 262006
rect 291471 262001 291537 262004
rect 584367 262001 584433 262004
rect 291759 261916 291825 261919
rect 591567 261916 591633 261919
rect 291759 261914 591633 261916
rect 291759 261858 291764 261914
rect 291820 261858 591572 261914
rect 591628 261858 591633 261914
rect 291759 261856 591633 261858
rect 291759 261853 291825 261856
rect 591567 261853 591633 261856
rect 674946 261771 675006 261886
rect 292143 261768 292209 261771
rect 595119 261768 595185 261771
rect 292143 261766 595185 261768
rect 292143 261710 292148 261766
rect 292204 261710 595124 261766
rect 595180 261710 595185 261766
rect 292143 261708 595185 261710
rect 292143 261705 292209 261708
rect 595119 261705 595185 261708
rect 674895 261766 675006 261771
rect 674895 261710 674900 261766
rect 674956 261710 675006 261766
rect 674895 261708 675006 261710
rect 674895 261705 674961 261708
rect 43791 261620 43857 261623
rect 42336 261618 43857 261620
rect 42336 261562 43796 261618
rect 43852 261562 43857 261618
rect 42336 261560 43857 261562
rect 43791 261557 43857 261560
rect 292527 261620 292593 261623
rect 602223 261620 602289 261623
rect 292527 261618 602289 261620
rect 292527 261562 292532 261618
rect 292588 261562 602228 261618
rect 602284 261562 602289 261618
rect 292527 261560 602289 261562
rect 292527 261557 292593 261560
rect 602223 261557 602289 261560
rect 292911 261472 292977 261475
rect 609327 261472 609393 261475
rect 292911 261470 609393 261472
rect 292911 261414 292916 261470
rect 292972 261414 609332 261470
rect 609388 261414 609393 261470
rect 292911 261412 609393 261414
rect 292911 261409 292977 261412
rect 609327 261409 609393 261412
rect 293295 261324 293361 261327
rect 612975 261324 613041 261327
rect 293295 261322 613041 261324
rect 293295 261266 293300 261322
rect 293356 261266 612980 261322
rect 613036 261266 613041 261322
rect 293295 261264 613041 261266
rect 293295 261261 293361 261264
rect 612975 261261 613041 261264
rect 293967 261176 294033 261179
rect 623631 261176 623697 261179
rect 293967 261174 623697 261176
rect 293967 261118 293972 261174
rect 294028 261118 623636 261174
rect 623692 261118 623697 261174
rect 293967 261116 623697 261118
rect 293967 261113 294033 261116
rect 623631 261113 623697 261116
rect 674127 261176 674193 261179
rect 674754 261176 674814 261220
rect 674127 261174 674814 261176
rect 674127 261118 674132 261174
rect 674188 261118 674814 261174
rect 674127 261116 674814 261118
rect 674127 261113 674193 261116
rect 294351 261028 294417 261031
rect 627183 261028 627249 261031
rect 294351 261026 627249 261028
rect 294351 260970 294356 261026
rect 294412 260970 627188 261026
rect 627244 260970 627249 261026
rect 294351 260968 627249 260970
rect 294351 260965 294417 260968
rect 627183 260965 627249 260968
rect 43215 260880 43281 260883
rect 42336 260878 43281 260880
rect 42336 260822 43220 260878
rect 43276 260822 43281 260878
rect 42336 260820 43281 260822
rect 43215 260817 43281 260820
rect 294735 260880 294801 260883
rect 634287 260880 634353 260883
rect 294735 260878 634353 260880
rect 294735 260822 294740 260878
rect 294796 260822 634292 260878
rect 634348 260822 634353 260878
rect 294735 260820 634353 260822
rect 294735 260817 294801 260820
rect 634287 260817 634353 260820
rect 198735 260732 198801 260735
rect 295119 260732 295185 260735
rect 641487 260732 641553 260735
rect 198735 260730 204414 260732
rect 198735 260674 198740 260730
rect 198796 260674 204414 260730
rect 198735 260672 204414 260674
rect 198735 260669 198801 260672
rect 204354 260584 204414 260672
rect 295119 260730 641553 260732
rect 295119 260674 295124 260730
rect 295180 260674 641492 260730
rect 641548 260674 641553 260730
rect 295119 260672 641553 260674
rect 295119 260669 295185 260672
rect 641487 260669 641553 260672
rect 218799 260584 218865 260587
rect 204354 260582 218865 260584
rect 204354 260526 218804 260582
rect 218860 260526 218865 260582
rect 204354 260524 218865 260526
rect 218799 260521 218865 260524
rect 295503 260584 295569 260587
rect 645039 260584 645105 260587
rect 295503 260582 645105 260584
rect 295503 260526 295508 260582
rect 295564 260526 645044 260582
rect 645100 260526 645105 260582
rect 295503 260524 645105 260526
rect 295503 260521 295569 260524
rect 645039 260521 645105 260524
rect 299631 260436 299697 260439
rect 309135 260436 309201 260439
rect 299631 260434 309201 260436
rect 299631 260378 299636 260434
rect 299692 260378 309140 260434
rect 309196 260378 309201 260434
rect 299631 260376 309201 260378
rect 299631 260373 299697 260376
rect 309135 260373 309201 260376
rect 327471 260436 327537 260439
rect 560655 260436 560721 260439
rect 327471 260434 560721 260436
rect 327471 260378 327476 260434
rect 327532 260378 560660 260434
rect 560716 260378 560721 260434
rect 327471 260376 560721 260378
rect 327471 260373 327537 260376
rect 560655 260373 560721 260376
rect 327087 260288 327153 260291
rect 557007 260288 557073 260291
rect 327087 260286 557073 260288
rect 327087 260230 327092 260286
rect 327148 260230 557012 260286
rect 557068 260230 557073 260286
rect 327087 260228 557073 260230
rect 327087 260225 327153 260228
rect 557007 260225 557073 260228
rect 675138 260143 675198 260406
rect 43311 260140 43377 260143
rect 42336 260138 43377 260140
rect 42336 260082 43316 260138
rect 43372 260082 43377 260138
rect 42336 260080 43377 260082
rect 43311 260077 43377 260080
rect 314991 260140 315057 260143
rect 545199 260140 545265 260143
rect 314991 260138 545265 260140
rect 314991 260082 314996 260138
rect 315052 260082 545204 260138
rect 545260 260082 545265 260138
rect 314991 260080 545265 260082
rect 314991 260077 315057 260080
rect 545199 260077 545265 260080
rect 675087 260138 675198 260143
rect 675087 260082 675092 260138
rect 675148 260082 675198 260138
rect 675087 260080 675198 260082
rect 675087 260077 675153 260080
rect 334479 259992 334545 259995
rect 426831 259992 426897 259995
rect 334479 259990 426897 259992
rect 334479 259934 334484 259990
rect 334540 259934 426836 259990
rect 426892 259934 426897 259990
rect 334479 259932 426897 259934
rect 334479 259929 334545 259932
rect 426831 259929 426897 259932
rect 40570 259486 40576 259550
rect 40640 259486 40646 259550
rect 40578 259400 40638 259486
rect 674946 259403 675006 259592
rect 43599 259400 43665 259403
rect 40578 259398 43665 259400
rect 40578 259370 43604 259398
rect 40608 259342 43604 259370
rect 43660 259342 43665 259398
rect 40608 259340 43665 259342
rect 674946 259398 675057 259403
rect 674946 259342 674996 259398
rect 675052 259342 675057 259398
rect 674946 259340 675057 259342
rect 43599 259337 43665 259340
rect 674991 259337 675057 259340
rect 65871 259104 65937 259107
rect 391599 259104 391665 259107
rect 65871 259102 391665 259104
rect 65871 259046 65876 259102
rect 65932 259046 391604 259102
rect 391660 259046 391665 259102
rect 65871 259044 391665 259046
rect 65871 259041 65937 259044
rect 391599 259041 391665 259044
rect 420975 259104 421041 259107
rect 443194 259104 443200 259106
rect 420975 259102 443200 259104
rect 420975 259046 420980 259102
rect 421036 259046 443200 259102
rect 420975 259044 443200 259046
rect 420975 259041 421041 259044
rect 443194 259042 443200 259044
rect 443264 259042 443270 259106
rect 70575 258956 70641 258959
rect 371439 258956 371505 258959
rect 70575 258954 371505 258956
rect 70575 258898 70580 258954
rect 70636 258898 371444 258954
rect 371500 258898 371505 258954
rect 70575 258896 371505 258898
rect 70575 258893 70641 258896
rect 371439 258893 371505 258896
rect 414735 258956 414801 258959
rect 442618 258956 442624 258958
rect 414735 258954 442624 258956
rect 414735 258898 414740 258954
rect 414796 258898 442624 258954
rect 414735 258896 442624 258898
rect 414735 258893 414801 258896
rect 442618 258894 442624 258896
rect 442688 258894 442694 258958
rect 74127 258808 74193 258811
rect 367119 258808 367185 258811
rect 74127 258806 367185 258808
rect 74127 258750 74132 258806
rect 74188 258750 367124 258806
rect 367180 258750 367185 258806
rect 74127 258748 367185 258750
rect 74127 258745 74193 258748
rect 367119 258745 367185 258748
rect 411759 258808 411825 258811
rect 442810 258808 442816 258810
rect 411759 258806 442816 258808
rect 411759 258750 411764 258806
rect 411820 258750 442816 258806
rect 411759 258748 442816 258750
rect 411759 258745 411825 258748
rect 442810 258746 442816 258748
rect 442880 258746 442886 258810
rect 674319 258808 674385 258811
rect 674319 258806 674784 258808
rect 674319 258750 674324 258806
rect 674380 258750 674784 258806
rect 674319 258748 674784 258750
rect 674319 258745 674385 258748
rect 76527 258660 76593 258663
rect 367791 258660 367857 258663
rect 76527 258658 367857 258660
rect 76527 258602 76532 258658
rect 76588 258602 367796 258658
rect 367852 258602 367857 258658
rect 76527 258600 367857 258602
rect 76527 258597 76593 258600
rect 367791 258597 367857 258600
rect 415119 258660 415185 258663
rect 446842 258660 446848 258662
rect 415119 258658 446848 258660
rect 415119 258602 415124 258658
rect 415180 258602 446848 258658
rect 415119 258600 446848 258602
rect 415119 258597 415185 258600
rect 446842 258598 446848 258600
rect 446912 258598 446918 258662
rect 78927 258512 78993 258515
rect 367599 258512 367665 258515
rect 78927 258510 367665 258512
rect 40386 257922 40446 258482
rect 78927 258454 78932 258510
rect 78988 258454 367604 258510
rect 367660 258454 367665 258510
rect 78927 258452 367665 258454
rect 78927 258449 78993 258452
rect 367599 258449 367665 258452
rect 413199 258512 413265 258515
rect 451066 258512 451072 258514
rect 413199 258510 451072 258512
rect 413199 258454 413204 258510
rect 413260 258454 451072 258510
rect 413199 258452 451072 258454
rect 413199 258449 413265 258452
rect 451066 258450 451072 258452
rect 451136 258450 451142 258514
rect 86031 258364 86097 258367
rect 370287 258364 370353 258367
rect 86031 258362 370353 258364
rect 86031 258306 86036 258362
rect 86092 258306 370292 258362
rect 370348 258306 370353 258362
rect 86031 258304 370353 258306
rect 86031 258301 86097 258304
rect 370287 258301 370353 258304
rect 412527 258364 412593 258367
rect 446074 258364 446080 258366
rect 412527 258362 446080 258364
rect 412527 258306 412532 258362
rect 412588 258306 446080 258362
rect 412527 258304 446080 258306
rect 412527 258301 412593 258304
rect 446074 258302 446080 258304
rect 446144 258302 446150 258366
rect 91983 258216 92049 258219
rect 435663 258216 435729 258219
rect 91983 258214 435729 258216
rect 91983 258158 91988 258214
rect 92044 258158 435668 258214
rect 435724 258158 435729 258214
rect 91983 258156 435729 258158
rect 91983 258153 92049 258156
rect 435663 258153 435729 258156
rect 87183 258068 87249 258071
rect 435279 258068 435345 258071
rect 87183 258066 435345 258068
rect 87183 258010 87188 258066
rect 87244 258010 435284 258066
rect 435340 258010 435345 258066
rect 87183 258008 435345 258010
rect 87183 258005 87249 258008
rect 435279 258005 435345 258008
rect 40378 257858 40384 257922
rect 40448 257858 40454 257922
rect 96783 257920 96849 257923
rect 448143 257920 448209 257923
rect 96783 257918 448209 257920
rect 96783 257862 96788 257918
rect 96844 257862 448148 257918
rect 448204 257862 448209 257918
rect 96783 257860 448209 257862
rect 96783 257857 96849 257860
rect 448143 257857 448209 257860
rect 88431 257772 88497 257775
rect 447471 257772 447537 257775
rect 88431 257770 447537 257772
rect 42306 257183 42366 257742
rect 88431 257714 88436 257770
rect 88492 257714 447476 257770
rect 447532 257714 447537 257770
rect 88431 257712 447537 257714
rect 88431 257709 88497 257712
rect 447471 257709 447537 257712
rect 282543 257624 282609 257627
rect 434223 257624 434289 257627
rect 282543 257622 434289 257624
rect 282543 257566 282548 257622
rect 282604 257566 434228 257622
rect 434284 257566 434289 257622
rect 282543 257564 434289 257566
rect 282543 257561 282609 257564
rect 434223 257561 434289 257564
rect 679746 257479 679806 257964
rect 289594 257414 289600 257478
rect 289664 257476 289670 257478
rect 290746 257476 290752 257478
rect 289664 257416 290752 257476
rect 289664 257414 289670 257416
rect 290746 257414 290752 257416
rect 290816 257414 290822 257478
rect 333999 257476 334065 257479
rect 426063 257476 426129 257479
rect 333999 257474 426129 257476
rect 333999 257418 334004 257474
rect 334060 257418 426068 257474
rect 426124 257418 426129 257474
rect 333999 257416 426129 257418
rect 333999 257413 334065 257416
rect 426063 257413 426129 257416
rect 679695 257474 679806 257479
rect 679695 257418 679700 257474
rect 679756 257418 679806 257474
rect 679695 257416 679806 257418
rect 679695 257413 679761 257416
rect 378447 257328 378513 257331
rect 388431 257328 388497 257331
rect 378447 257326 388497 257328
rect 378447 257270 378452 257326
rect 378508 257270 388436 257326
rect 388492 257270 388497 257326
rect 378447 257268 388497 257270
rect 378447 257265 378513 257268
rect 388431 257265 388497 257268
rect 409551 257328 409617 257331
rect 441466 257328 441472 257330
rect 409551 257326 441472 257328
rect 409551 257270 409556 257326
rect 409612 257270 441472 257326
rect 409551 257268 441472 257270
rect 409551 257265 409617 257268
rect 441466 257266 441472 257268
rect 441536 257266 441542 257330
rect 674938 257266 674944 257330
rect 675008 257328 675014 257330
rect 675514 257328 675520 257330
rect 675008 257268 675520 257328
rect 675008 257266 675014 257268
rect 675514 257266 675520 257268
rect 675584 257266 675590 257330
rect 42255 257178 42366 257183
rect 351471 257182 351537 257183
rect 351418 257180 351424 257182
rect 42255 257122 42260 257178
rect 42316 257122 42366 257178
rect 42255 257120 42366 257122
rect 351380 257120 351424 257180
rect 351488 257178 351537 257182
rect 351532 257122 351537 257178
rect 42255 257117 42321 257120
rect 351418 257118 351424 257120
rect 351488 257118 351537 257122
rect 351471 257117 351537 257118
rect 383151 257180 383217 257183
rect 397071 257180 397137 257183
rect 383151 257178 397137 257180
rect 383151 257122 383156 257178
rect 383212 257122 397076 257178
rect 397132 257122 397137 257178
rect 383151 257120 397137 257122
rect 383151 257117 383217 257120
rect 397071 257117 397137 257120
rect 412911 257180 412977 257183
rect 448378 257180 448384 257182
rect 412911 257178 448384 257180
rect 412911 257122 412916 257178
rect 412972 257122 448384 257178
rect 412911 257120 448384 257122
rect 412911 257117 412977 257120
rect 448378 257118 448384 257120
rect 448448 257118 448454 257182
rect 321999 257032 322065 257035
rect 445114 257032 445120 257034
rect 321999 257030 445120 257032
rect 321999 256974 322004 257030
rect 322060 256974 445120 257030
rect 321999 256972 445120 256974
rect 321999 256969 322065 256972
rect 445114 256970 445120 256972
rect 445184 256970 445190 257034
rect 40578 256442 40638 256854
rect 287098 256822 287104 256886
rect 287168 256884 287174 256886
rect 319023 256884 319089 256887
rect 287168 256847 287934 256884
rect 288018 256882 319089 256884
rect 288018 256847 319028 256882
rect 287168 256826 319028 256847
rect 319084 256826 319089 256882
rect 287168 256824 319089 256826
rect 287168 256822 287174 256824
rect 287874 256787 288078 256824
rect 319023 256821 319089 256824
rect 320175 256884 320241 256887
rect 445306 256884 445312 256886
rect 320175 256882 445312 256884
rect 320175 256826 320180 256882
rect 320236 256826 445312 256882
rect 320175 256824 445312 256826
rect 320175 256821 320241 256824
rect 445306 256822 445312 256824
rect 445376 256822 445382 256886
rect 679695 256884 679761 256887
rect 679695 256882 679806 256884
rect 679695 256826 679700 256882
rect 679756 256826 679806 256882
rect 679695 256821 679806 256826
rect 300783 256736 300849 256739
rect 310863 256736 310929 256739
rect 300783 256734 310929 256736
rect 300783 256678 300788 256734
rect 300844 256678 310868 256734
rect 310924 256678 310929 256734
rect 300783 256676 310929 256678
rect 300783 256673 300849 256676
rect 310863 256673 310929 256676
rect 317967 256736 318033 256739
rect 443770 256736 443776 256738
rect 317967 256734 443776 256736
rect 317967 256678 317972 256734
rect 318028 256678 443776 256734
rect 317967 256676 443776 256678
rect 317967 256673 318033 256676
rect 443770 256674 443776 256676
rect 443840 256674 443846 256738
rect 292090 256526 292096 256590
rect 292160 256588 292166 256590
rect 310959 256588 311025 256591
rect 292160 256586 311025 256588
rect 292160 256530 310964 256586
rect 311020 256530 311025 256586
rect 292160 256528 311025 256530
rect 292160 256526 292166 256528
rect 310959 256525 311025 256528
rect 317199 256588 317265 256591
rect 447802 256588 447808 256590
rect 317199 256586 447808 256588
rect 317199 256530 317204 256586
rect 317260 256530 447808 256586
rect 317199 256528 447808 256530
rect 317199 256525 317265 256528
rect 447802 256526 447808 256528
rect 447872 256526 447878 256590
rect 40570 256378 40576 256442
rect 40640 256378 40646 256442
rect 286906 256378 286912 256442
rect 286976 256440 286982 256442
rect 424623 256440 424689 256443
rect 286976 256438 424689 256440
rect 286976 256382 424628 256438
rect 424684 256382 424689 256438
rect 679746 256410 679806 256821
rect 286976 256380 424689 256382
rect 286976 256378 286982 256380
rect 424623 256377 424689 256380
rect 286714 256230 286720 256294
rect 286784 256292 286790 256294
rect 424239 256292 424305 256295
rect 286784 256290 424305 256292
rect 286784 256234 424244 256290
rect 424300 256234 424305 256290
rect 286784 256232 424305 256234
rect 286784 256230 286790 256232
rect 424239 256229 424305 256232
rect 424431 256292 424497 256295
rect 448762 256292 448768 256294
rect 424431 256290 448768 256292
rect 424431 256234 424436 256290
rect 424492 256234 448768 256290
rect 424431 256232 448768 256234
rect 424431 256229 424497 256232
rect 448762 256230 448768 256232
rect 448832 256230 448838 256294
rect 676666 256230 676672 256294
rect 676736 256292 676742 256294
rect 680079 256292 680145 256295
rect 676736 256290 680145 256292
rect 676736 256234 680084 256290
rect 680140 256234 680145 256290
rect 676736 256232 680145 256234
rect 676736 256230 676742 256232
rect 680079 256229 680145 256232
rect 40962 255702 41022 256114
rect 290746 256082 290752 256146
rect 290816 256144 290822 256146
rect 319695 256144 319761 256147
rect 290816 256142 319761 256144
rect 290816 256086 319700 256142
rect 319756 256086 319761 256142
rect 290816 256084 319761 256086
rect 290816 256082 290822 256084
rect 319695 256081 319761 256084
rect 320463 256144 320529 256147
rect 408975 256144 409041 256147
rect 320463 256142 409041 256144
rect 320463 256086 320468 256142
rect 320524 256086 408980 256142
rect 409036 256086 409041 256142
rect 320463 256084 409041 256086
rect 320463 256081 320529 256084
rect 408975 256081 409041 256084
rect 443002 256082 443008 256146
rect 443072 256144 443078 256146
rect 448954 256144 448960 256146
rect 443072 256084 448960 256144
rect 443072 256082 443078 256084
rect 448954 256082 448960 256084
rect 449024 256082 449030 256146
rect 290938 255934 290944 255998
rect 291008 255996 291014 255998
rect 337210 255996 337216 255998
rect 291008 255936 337216 255996
rect 291008 255934 291014 255936
rect 337210 255934 337216 255936
rect 337280 255934 337286 255998
rect 337455 255996 337521 255999
rect 446650 255996 446656 255998
rect 337455 255994 446656 255996
rect 337455 255938 337460 255994
rect 337516 255938 446656 255994
rect 337455 255936 446656 255938
rect 337455 255933 337521 255936
rect 446650 255934 446656 255936
rect 446720 255934 446726 255998
rect 138159 255848 138225 255851
rect 118146 255846 138225 255848
rect 118146 255790 138164 255846
rect 138220 255790 138225 255846
rect 118146 255788 138225 255790
rect 118146 255703 118206 255788
rect 138159 255785 138225 255788
rect 291322 255786 291328 255850
rect 291392 255848 291398 255850
rect 351418 255848 351424 255850
rect 291392 255788 351424 255848
rect 291392 255786 291398 255788
rect 351418 255786 351424 255788
rect 351488 255786 351494 255850
rect 408975 255848 409041 255851
rect 421551 255848 421617 255851
rect 408975 255846 421617 255848
rect 408975 255790 408980 255846
rect 409036 255790 421556 255846
rect 421612 255790 421617 255846
rect 408975 255788 421617 255790
rect 408975 255785 409041 255788
rect 421551 255785 421617 255788
rect 421743 255848 421809 255851
rect 448570 255848 448576 255850
rect 421743 255846 448576 255848
rect 421743 255790 421748 255846
rect 421804 255790 448576 255846
rect 421743 255788 448576 255790
rect 421743 255785 421809 255788
rect 448570 255786 448576 255788
rect 448640 255786 448646 255850
rect 621999 255848 622065 255851
rect 601986 255846 622065 255848
rect 601986 255790 622004 255846
rect 622060 255790 622065 255846
rect 601986 255788 622065 255790
rect 601986 255703 602046 255788
rect 621999 255785 622065 255788
rect 40954 255638 40960 255702
rect 41024 255638 41030 255702
rect 80655 255700 80721 255703
rect 86703 255700 86769 255703
rect 80655 255698 86769 255700
rect 80655 255642 80660 255698
rect 80716 255642 86708 255698
rect 86764 255642 86769 255698
rect 80655 255640 86769 255642
rect 80655 255637 80721 255640
rect 86703 255637 86769 255640
rect 118095 255698 118206 255703
rect 118095 255642 118100 255698
rect 118156 255642 118206 255698
rect 118095 255640 118206 255642
rect 118095 255637 118161 255640
rect 291706 255638 291712 255702
rect 291776 255700 291782 255702
rect 359343 255700 359409 255703
rect 291776 255698 359409 255700
rect 291776 255642 359348 255698
rect 359404 255642 359409 255698
rect 291776 255640 359409 255642
rect 291776 255638 291782 255640
rect 359343 255637 359409 255640
rect 410703 255700 410769 255703
rect 452986 255700 452992 255702
rect 410703 255698 452992 255700
rect 410703 255642 410708 255698
rect 410764 255642 452992 255698
rect 410703 255640 452992 255642
rect 410703 255637 410769 255640
rect 452986 255638 452992 255640
rect 453056 255638 453062 255702
rect 501135 255700 501201 255703
rect 501135 255698 538494 255700
rect 501135 255642 501140 255698
rect 501196 255666 538494 255698
rect 601935 255698 602046 255703
rect 501196 255661 538545 255666
rect 501196 255642 538484 255661
rect 501135 255640 538484 255642
rect 501135 255637 501201 255640
rect 538434 255605 538484 255640
rect 538540 255605 538545 255661
rect 601935 255642 601940 255698
rect 601996 255642 602046 255698
rect 601935 255640 602046 255642
rect 642255 255700 642321 255703
rect 671055 255700 671121 255703
rect 673978 255700 673984 255702
rect 642255 255698 642366 255700
rect 642255 255642 642260 255698
rect 642316 255642 642366 255698
rect 601935 255637 602001 255640
rect 642255 255637 642366 255642
rect 671055 255698 673984 255700
rect 671055 255642 671060 255698
rect 671116 255642 673984 255698
rect 671055 255640 673984 255642
rect 671055 255637 671121 255640
rect 673978 255638 673984 255640
rect 674048 255638 674054 255702
rect 538434 255603 538545 255605
rect 538479 255600 538545 255603
rect 291898 255490 291904 255554
rect 291968 255552 291974 255554
rect 364431 255552 364497 255555
rect 291968 255550 364497 255552
rect 291968 255494 364436 255550
rect 364492 255494 364497 255550
rect 291968 255492 364497 255494
rect 291968 255490 291974 255492
rect 364431 255489 364497 255492
rect 419151 255552 419217 255555
rect 448186 255552 448192 255554
rect 419151 255550 448192 255552
rect 419151 255494 419156 255550
rect 419212 255494 448192 255550
rect 419151 255492 448192 255494
rect 419151 255489 419217 255492
rect 448186 255490 448192 255492
rect 448256 255490 448262 255554
rect 642306 255552 642366 255637
rect 662319 255552 662385 255555
rect 642306 255550 662385 255552
rect 642306 255494 662324 255550
rect 662380 255494 662385 255550
rect 642306 255492 662385 255494
rect 662319 255489 662385 255492
rect 41346 254814 41406 255374
rect 292282 255342 292288 255406
rect 292352 255404 292358 255406
rect 364335 255404 364401 255407
rect 292352 255402 364401 255404
rect 292352 255346 364340 255402
rect 364396 255346 364401 255402
rect 292352 255344 364401 255346
rect 292352 255342 292358 255344
rect 364335 255341 364401 255344
rect 419823 255404 419889 255407
rect 453754 255404 453760 255406
rect 419823 255402 453760 255404
rect 419823 255346 419828 255402
rect 419884 255346 453760 255402
rect 419823 255344 453760 255346
rect 419823 255341 419889 255344
rect 453754 255342 453760 255344
rect 453824 255342 453830 255406
rect 292666 255194 292672 255258
rect 292736 255256 292742 255258
rect 377775 255256 377841 255259
rect 292736 255254 377841 255256
rect 292736 255198 377780 255254
rect 377836 255198 377841 255254
rect 292736 255196 377841 255198
rect 292736 255194 292742 255196
rect 377775 255193 377841 255196
rect 409935 255256 410001 255259
rect 439023 255256 439089 255259
rect 453178 255256 453184 255258
rect 409935 255254 439089 255256
rect 409935 255198 409940 255254
rect 409996 255198 439028 255254
rect 439084 255198 439089 255254
rect 409935 255196 439089 255198
rect 409935 255193 410001 255196
rect 439023 255193 439089 255196
rect 439170 255196 453184 255256
rect 293050 255046 293056 255110
rect 293120 255108 293126 255110
rect 383439 255108 383505 255111
rect 293120 255106 383505 255108
rect 293120 255050 383444 255106
rect 383500 255050 383505 255106
rect 293120 255048 383505 255050
rect 293120 255046 293126 255048
rect 383439 255045 383505 255048
rect 418767 255108 418833 255111
rect 439170 255108 439230 255196
rect 453178 255194 453184 255196
rect 453248 255194 453254 255258
rect 453370 255108 453376 255110
rect 418767 255106 439230 255108
rect 418767 255050 418772 255106
rect 418828 255050 439230 255106
rect 418767 255048 439230 255050
rect 439362 255048 453376 255108
rect 418767 255045 418833 255048
rect 65007 254960 65073 254963
rect 204922 254960 204928 254962
rect 65007 254958 204928 254960
rect 65007 254902 65012 254958
rect 65068 254902 204928 254958
rect 65007 254900 204928 254902
rect 65007 254897 65073 254900
rect 204922 254898 204928 254900
rect 204992 254898 204998 254962
rect 293242 254898 293248 254962
rect 293312 254960 293318 254962
rect 389967 254960 390033 254963
rect 293312 254958 390033 254960
rect 293312 254902 389972 254958
rect 390028 254902 390033 254958
rect 293312 254900 390033 254902
rect 293312 254898 293318 254900
rect 389967 254897 390033 254900
rect 410319 254960 410385 254963
rect 439362 254960 439422 255048
rect 453370 255046 453376 255048
rect 453440 255046 453446 255110
rect 410319 254958 439422 254960
rect 410319 254902 410324 254958
rect 410380 254902 439422 254958
rect 410319 254900 439422 254902
rect 439503 254960 439569 254963
rect 454138 254960 454144 254962
rect 439503 254958 454144 254960
rect 439503 254902 439508 254958
rect 439564 254902 454144 254958
rect 439503 254900 454144 254902
rect 410319 254897 410385 254900
rect 439503 254897 439569 254900
rect 454138 254898 454144 254900
rect 454208 254898 454214 254962
rect 41338 254750 41344 254814
rect 41408 254750 41414 254814
rect 65103 254812 65169 254815
rect 204730 254812 204736 254814
rect 65103 254810 204736 254812
rect 65103 254754 65108 254810
rect 65164 254754 204736 254810
rect 65103 254752 204736 254754
rect 65103 254749 65169 254752
rect 204730 254750 204736 254752
rect 204800 254750 204806 254814
rect 289167 254812 289233 254815
rect 387279 254812 387345 254815
rect 289167 254810 387345 254812
rect 289167 254754 289172 254810
rect 289228 254754 387284 254810
rect 387340 254754 387345 254810
rect 289167 254752 387345 254754
rect 289167 254749 289233 254752
rect 387279 254749 387345 254752
rect 417615 254812 417681 254815
rect 449914 254812 449920 254814
rect 417615 254810 449920 254812
rect 417615 254754 417620 254810
rect 417676 254754 449920 254810
rect 417615 254752 449920 254754
rect 417615 254749 417681 254752
rect 449914 254750 449920 254752
rect 449984 254750 449990 254814
rect 284218 254602 284224 254666
rect 284288 254664 284294 254666
rect 322575 254664 322641 254667
rect 284288 254662 322641 254664
rect 284288 254606 322580 254662
rect 322636 254606 322641 254662
rect 284288 254604 322641 254606
rect 284288 254602 284294 254604
rect 322575 254601 322641 254604
rect 324879 254664 324945 254667
rect 337455 254664 337521 254667
rect 324879 254662 337521 254664
rect 324879 254606 324884 254662
rect 324940 254606 337460 254662
rect 337516 254606 337521 254662
rect 324879 254604 337521 254606
rect 324879 254601 324945 254604
rect 337455 254601 337521 254604
rect 337594 254602 337600 254666
rect 337664 254664 337670 254666
rect 345039 254664 345105 254667
rect 453946 254664 453952 254666
rect 337664 254662 345105 254664
rect 337664 254606 345044 254662
rect 345100 254606 345105 254662
rect 337664 254604 345105 254606
rect 337664 254602 337670 254604
rect 345039 254601 345105 254604
rect 439170 254604 453952 254664
rect 37314 254075 37374 254560
rect 287290 254454 287296 254518
rect 287360 254516 287366 254518
rect 425391 254516 425457 254519
rect 287360 254514 425457 254516
rect 287360 254458 425396 254514
rect 425452 254458 425457 254514
rect 287360 254456 425457 254458
rect 287360 254454 287366 254456
rect 425391 254453 425457 254456
rect 425679 254516 425745 254519
rect 439170 254516 439230 254604
rect 453946 254602 453952 254604
rect 454016 254602 454022 254666
rect 425679 254514 439230 254516
rect 425679 254458 425684 254514
rect 425740 254458 439230 254514
rect 425679 254456 439230 254458
rect 440655 254516 440721 254519
rect 441850 254516 441856 254518
rect 440655 254514 441856 254516
rect 440655 254458 440660 254514
rect 440716 254458 441856 254514
rect 440655 254456 441856 254458
rect 425679 254453 425745 254456
rect 440655 254453 440721 254456
rect 441850 254454 441856 254456
rect 441920 254454 441926 254518
rect 443535 254516 443601 254519
rect 444154 254516 444160 254518
rect 443535 254514 444160 254516
rect 443535 254458 443540 254514
rect 443596 254458 444160 254514
rect 443535 254456 444160 254458
rect 443535 254453 443601 254456
rect 444154 254454 444160 254456
rect 444224 254454 444230 254518
rect 324495 254368 324561 254371
rect 316290 254366 324561 254368
rect 316290 254310 324500 254366
rect 324556 254310 324561 254366
rect 316290 254308 324561 254310
rect 293434 254158 293440 254222
rect 293504 254220 293510 254222
rect 316290 254220 316350 254308
rect 324495 254305 324561 254308
rect 325263 254368 325329 254371
rect 437007 254368 437073 254371
rect 325263 254366 437073 254368
rect 325263 254310 325268 254366
rect 325324 254310 437012 254366
rect 437068 254310 437073 254366
rect 325263 254308 437073 254310
rect 325263 254305 325329 254308
rect 437007 254305 437073 254308
rect 440751 254368 440817 254371
rect 442426 254368 442432 254370
rect 440751 254366 442432 254368
rect 440751 254310 440756 254366
rect 440812 254310 442432 254366
rect 440751 254308 442432 254310
rect 440751 254305 440817 254308
rect 442426 254306 442432 254308
rect 442496 254306 442502 254370
rect 443631 254368 443697 254371
rect 444346 254368 444352 254370
rect 443631 254366 444352 254368
rect 443631 254310 443636 254366
rect 443692 254310 444352 254366
rect 443631 254308 444352 254310
rect 443631 254305 443697 254308
rect 444346 254306 444352 254308
rect 444416 254306 444422 254370
rect 446415 254368 446481 254371
rect 447610 254368 447616 254370
rect 446415 254366 447616 254368
rect 446415 254310 446420 254366
rect 446476 254310 447616 254366
rect 446415 254308 447616 254310
rect 446415 254305 446481 254308
rect 447610 254306 447616 254308
rect 447680 254306 447686 254370
rect 293504 254160 316350 254220
rect 319695 254220 319761 254223
rect 321231 254220 321297 254223
rect 319695 254218 321297 254220
rect 319695 254162 319700 254218
rect 319756 254162 321236 254218
rect 321292 254162 321297 254218
rect 319695 254160 321297 254162
rect 293504 254158 293510 254160
rect 319695 254157 319761 254160
rect 321231 254157 321297 254160
rect 323823 254220 323889 254223
rect 444538 254220 444544 254222
rect 323823 254218 444544 254220
rect 323823 254162 323828 254218
rect 323884 254162 444544 254218
rect 323823 254160 444544 254162
rect 323823 254157 323889 254160
rect 444538 254158 444544 254160
rect 444608 254158 444614 254222
rect 446415 254220 446481 254223
rect 447994 254220 448000 254222
rect 446415 254218 448000 254220
rect 446415 254162 446420 254218
rect 446476 254162 448000 254218
rect 446415 254160 448000 254162
rect 446415 254157 446481 254160
rect 447994 254158 448000 254160
rect 448064 254158 448070 254222
rect 37263 254070 37374 254075
rect 37263 254014 37268 254070
rect 37324 254014 37374 254070
rect 37263 254012 37374 254014
rect 37263 254009 37329 254012
rect 288058 254010 288064 254074
rect 288128 254072 288134 254074
rect 315663 254072 315729 254075
rect 288128 254070 315729 254072
rect 288128 254014 315668 254070
rect 315724 254014 315729 254070
rect 288128 254012 315729 254014
rect 288128 254010 288134 254012
rect 315663 254009 315729 254012
rect 316719 254072 316785 254075
rect 322575 254072 322641 254075
rect 316719 254070 322641 254072
rect 316719 254014 316724 254070
rect 316780 254014 322580 254070
rect 322636 254014 322641 254070
rect 316719 254012 322641 254014
rect 316719 254009 316785 254012
rect 322575 254009 322641 254012
rect 323439 254072 323505 254075
rect 443962 254072 443968 254074
rect 323439 254070 443968 254072
rect 323439 254014 323444 254070
rect 323500 254014 443968 254070
rect 323439 254012 443968 254014
rect 323439 254009 323505 254012
rect 443962 254010 443968 254012
rect 444032 254010 444038 254074
rect 444303 254072 444369 254075
rect 451258 254072 451264 254074
rect 444303 254070 451264 254072
rect 444303 254014 444308 254070
rect 444364 254014 451264 254070
rect 444303 254012 451264 254014
rect 444303 254009 444369 254012
rect 451258 254010 451264 254012
rect 451328 254010 451334 254074
rect 288207 253924 288273 253927
rect 322671 253924 322737 253927
rect 288207 253922 322737 253924
rect 288207 253866 288212 253922
rect 288268 253866 322676 253922
rect 322732 253866 322737 253922
rect 288207 253864 322737 253866
rect 288207 253861 288273 253864
rect 322671 253861 322737 253864
rect 418383 253924 418449 253927
rect 452602 253924 452608 253926
rect 418383 253922 452608 253924
rect 418383 253866 418388 253922
rect 418444 253866 452608 253922
rect 418383 253864 452608 253866
rect 418383 253861 418449 253864
rect 452602 253862 452608 253864
rect 452672 253862 452678 253926
rect 40770 253482 40830 253746
rect 288250 253714 288256 253778
rect 288320 253776 288326 253778
rect 316431 253776 316497 253779
rect 319407 253776 319473 253779
rect 288320 253774 316497 253776
rect 288320 253718 316436 253774
rect 316492 253718 316497 253774
rect 288320 253716 316497 253718
rect 288320 253714 288326 253716
rect 316431 253713 316497 253716
rect 316674 253774 319473 253776
rect 316674 253718 319412 253774
rect 319468 253718 319473 253774
rect 316674 253716 319473 253718
rect 288442 253566 288448 253630
rect 288512 253628 288518 253630
rect 316674 253628 316734 253716
rect 319407 253713 319473 253716
rect 416175 253776 416241 253779
rect 452794 253776 452800 253778
rect 416175 253774 452800 253776
rect 416175 253718 416180 253774
rect 416236 253718 452800 253774
rect 416175 253716 452800 253718
rect 416175 253713 416241 253716
rect 452794 253714 452800 253716
rect 452864 253714 452870 253778
rect 288512 253568 316734 253628
rect 419535 253628 419601 253631
rect 441658 253628 441664 253630
rect 419535 253626 441664 253628
rect 419535 253570 419540 253626
rect 419596 253570 441664 253626
rect 419535 253568 441664 253570
rect 288512 253566 288518 253568
rect 419535 253565 419601 253568
rect 441658 253566 441664 253568
rect 441728 253566 441734 253630
rect 442618 253566 442624 253630
rect 442688 253628 442694 253630
rect 445882 253628 445888 253630
rect 442688 253568 445888 253628
rect 442688 253566 442694 253568
rect 445882 253566 445888 253568
rect 445952 253566 445958 253630
rect 40762 253418 40768 253482
rect 40832 253418 40838 253482
rect 288826 253418 288832 253482
rect 288896 253480 288902 253482
rect 318639 253480 318705 253483
rect 288896 253478 318705 253480
rect 288896 253422 318644 253478
rect 318700 253422 318705 253478
rect 288896 253420 318705 253422
rect 288896 253418 288902 253420
rect 318639 253417 318705 253420
rect 410991 253480 411057 253483
rect 425679 253480 425745 253483
rect 410991 253478 425745 253480
rect 410991 253422 410996 253478
rect 411052 253422 425684 253478
rect 425740 253422 425745 253478
rect 410991 253420 425745 253422
rect 410991 253417 411057 253420
rect 425679 253417 425745 253420
rect 437007 253480 437073 253483
rect 444922 253480 444928 253482
rect 437007 253478 444928 253480
rect 437007 253422 437012 253478
rect 437068 253422 444928 253478
rect 437007 253420 444928 253422
rect 437007 253417 437073 253420
rect 444922 253418 444928 253420
rect 444992 253418 444998 253482
rect 445359 253480 445425 253483
rect 450106 253480 450112 253482
rect 445359 253478 450112 253480
rect 445359 253422 445364 253478
rect 445420 253422 450112 253478
rect 445359 253420 450112 253422
rect 445359 253417 445425 253420
rect 450106 253418 450112 253420
rect 450176 253418 450182 253482
rect 282831 253332 282897 253335
rect 283066 253332 283072 253334
rect 282831 253330 283072 253332
rect 282831 253274 282836 253330
rect 282892 253274 283072 253330
rect 282831 253272 283072 253274
rect 282831 253269 282897 253272
rect 283066 253270 283072 253272
rect 283136 253270 283142 253334
rect 292474 253270 292480 253334
rect 292544 253332 292550 253334
rect 293199 253332 293265 253335
rect 444730 253332 444736 253334
rect 292544 253330 293265 253332
rect 292544 253274 293204 253330
rect 293260 253274 293265 253330
rect 292544 253272 293265 253274
rect 292544 253270 292550 253272
rect 293199 253269 293265 253272
rect 436866 253272 444736 253332
rect 413583 253184 413649 253187
rect 436866 253184 436926 253272
rect 444730 253270 444736 253272
rect 444800 253270 444806 253334
rect 444975 253332 445041 253335
rect 450490 253332 450496 253334
rect 444975 253330 450496 253332
rect 444975 253274 444980 253330
rect 445036 253274 450496 253330
rect 444975 253272 450496 253274
rect 444975 253269 445041 253272
rect 450490 253270 450496 253272
rect 450560 253270 450566 253334
rect 450874 253184 450880 253186
rect 413583 253182 436926 253184
rect 413583 253126 413588 253182
rect 413644 253126 436926 253182
rect 413583 253124 436926 253126
rect 439170 253124 450880 253184
rect 413583 253121 413649 253124
rect 286522 252974 286528 253038
rect 286592 253036 286598 253038
rect 287823 253036 287889 253039
rect 286592 253034 287889 253036
rect 286592 252978 287828 253034
rect 287884 252978 287889 253034
rect 286592 252976 287889 252978
rect 286592 252974 286598 252976
rect 287823 252973 287889 252976
rect 288634 252974 288640 253038
rect 288704 253036 288710 253038
rect 288879 253036 288945 253039
rect 289167 253036 289233 253039
rect 289455 253038 289521 253039
rect 289402 253036 289408 253038
rect 288704 253034 288945 253036
rect 288704 252978 288884 253034
rect 288940 252978 288945 253034
rect 288704 252976 288945 252978
rect 288704 252974 288710 252976
rect 288879 252973 288945 252976
rect 289026 253034 289233 253036
rect 289026 252978 289172 253034
rect 289228 252978 289233 253034
rect 289026 252976 289233 252978
rect 289364 252976 289408 253036
rect 289472 253034 289521 253038
rect 289516 252978 289521 253034
rect 41154 252446 41214 252932
rect 289026 252888 289086 252976
rect 289167 252973 289233 252976
rect 289402 252974 289408 252976
rect 289472 252974 289521 252978
rect 291130 252974 291136 253038
rect 291200 253036 291206 253038
rect 295311 253036 295377 253039
rect 291200 253034 295377 253036
rect 291200 252978 295316 253034
rect 295372 252978 295377 253034
rect 291200 252976 295377 252978
rect 291200 252974 291206 252976
rect 289455 252973 289521 252974
rect 295311 252973 295377 252976
rect 415407 253036 415473 253039
rect 415791 253036 415857 253039
rect 439170 253036 439230 253124
rect 450874 253122 450880 253124
rect 450944 253122 450950 253186
rect 415407 253034 415614 253036
rect 415407 252978 415412 253034
rect 415468 252978 415614 253034
rect 415407 252976 415614 252978
rect 415407 252973 415473 252976
rect 288642 252828 289086 252888
rect 415554 252888 415614 252976
rect 415791 253034 439230 253036
rect 415791 252978 415796 253034
rect 415852 252978 439230 253034
rect 415791 252976 439230 252978
rect 440271 253036 440337 253039
rect 442618 253036 442624 253038
rect 440271 253034 442624 253036
rect 440271 252978 440276 253034
rect 440332 252978 442624 253034
rect 440271 252976 442624 252978
rect 415791 252973 415857 252976
rect 440271 252973 440337 252976
rect 442618 252974 442624 252976
rect 442688 252974 442694 253038
rect 443578 252974 443584 253038
rect 443648 252974 443654 253038
rect 445359 253034 445425 253039
rect 446223 253038 446289 253039
rect 446223 253036 446272 253038
rect 445359 252978 445364 253034
rect 445420 252978 445425 253034
rect 443586 252888 443646 252974
rect 445359 252973 445425 252978
rect 446180 253034 446272 253036
rect 446180 252978 446228 253034
rect 446180 252976 446272 252978
rect 446223 252974 446272 252976
rect 446336 252974 446342 253038
rect 446415 253036 446481 253039
rect 447418 253036 447424 253038
rect 446415 253034 447424 253036
rect 446415 252978 446420 253034
rect 446476 252978 447424 253034
rect 446415 252976 447424 252978
rect 446223 252973 446289 252974
rect 446415 252973 446481 252976
rect 447418 252974 447424 252976
rect 447488 252974 447494 253038
rect 453562 252974 453568 253038
rect 453632 252974 453638 253038
rect 415554 252828 443646 252888
rect 445362 252888 445422 252973
rect 453570 252888 453630 252974
rect 445362 252828 453630 252888
rect 41146 252382 41152 252446
rect 41216 252382 41222 252446
rect 45903 252148 45969 252151
rect 208378 252148 208384 252150
rect 45903 252146 208384 252148
rect 41922 251559 41982 252118
rect 45903 252090 45908 252146
rect 45964 252090 208384 252146
rect 45903 252088 208384 252090
rect 45903 252085 45969 252088
rect 208378 252086 208384 252088
rect 208448 252086 208454 252150
rect 45615 252000 45681 252003
rect 207418 252000 207424 252002
rect 45615 251998 207424 252000
rect 45615 251942 45620 251998
rect 45676 251942 207424 251998
rect 45615 251940 207424 251942
rect 45615 251937 45681 251940
rect 207418 251938 207424 251940
rect 207488 251938 207494 252002
rect 288642 251822 288702 252828
rect 41922 251554 42033 251559
rect 41922 251498 41972 251554
rect 42028 251498 42033 251554
rect 41922 251496 42033 251498
rect 41967 251493 42033 251496
rect 37314 250819 37374 251304
rect 283695 251260 283761 251263
rect 283695 251258 288288 251260
rect 283695 251202 283700 251258
rect 283756 251202 288288 251258
rect 283695 251200 288288 251202
rect 283695 251197 283761 251200
rect 288495 251112 288561 251115
rect 288450 251110 288561 251112
rect 288450 251054 288500 251110
rect 288556 251054 288561 251110
rect 288450 251049 288561 251054
rect 37167 250816 37233 250819
rect 37122 250814 37233 250816
rect 37122 250758 37172 250814
rect 37228 250758 37233 250814
rect 37122 250753 37233 250758
rect 37314 250814 37425 250819
rect 37314 250758 37364 250814
rect 37420 250758 37425 250814
rect 37314 250756 37425 250758
rect 37359 250753 37425 250756
rect 37122 250638 37182 250753
rect 145402 250668 145408 250670
rect 140802 250608 145408 250668
rect 140802 250566 140862 250608
rect 145402 250606 145408 250608
rect 145472 250606 145478 250670
rect 288450 250638 288510 251049
rect 283791 250224 283857 250227
rect 283791 250222 288288 250224
rect 283791 250166 283796 250222
rect 283852 250166 288288 250222
rect 283791 250164 288288 250166
rect 283791 250161 283857 250164
rect 43119 249780 43185 249783
rect 42336 249778 43185 249780
rect 42336 249722 43124 249778
rect 43180 249722 43185 249778
rect 42336 249720 43185 249722
rect 43119 249717 43185 249720
rect 282735 249632 282801 249635
rect 282735 249630 288288 249632
rect 282735 249574 282740 249630
rect 282796 249574 288288 249630
rect 282735 249572 288288 249574
rect 282735 249569 282801 249572
rect 674746 249570 674752 249634
rect 674816 249632 674822 249634
rect 675375 249632 675441 249635
rect 674816 249630 675441 249632
rect 674816 249574 675380 249630
rect 675436 249574 675441 249630
rect 674816 249572 675441 249574
rect 674816 249570 674822 249572
rect 675375 249569 675441 249572
rect 145455 249336 145521 249339
rect 140832 249334 145521 249336
rect 140832 249278 145460 249334
rect 145516 249278 145521 249334
rect 140832 249276 145521 249278
rect 145455 249273 145521 249276
rect 288015 249336 288081 249339
rect 288399 249336 288465 249339
rect 288015 249334 288465 249336
rect 288015 249278 288020 249334
rect 288076 249278 288404 249334
rect 288460 249278 288465 249334
rect 288015 249276 288465 249278
rect 288015 249273 288081 249276
rect 288399 249273 288465 249276
rect 283887 249040 283953 249043
rect 283887 249038 288288 249040
rect 42114 248451 42174 249010
rect 283887 248982 283892 249038
rect 283948 248982 288288 249038
rect 283887 248980 288288 248982
rect 283887 248977 283953 248980
rect 283119 248894 283185 248895
rect 283066 248830 283072 248894
rect 283136 248892 283185 248894
rect 288495 248892 288561 248895
rect 288634 248892 288640 248894
rect 283136 248890 283228 248892
rect 283180 248834 283228 248890
rect 283136 248832 283228 248834
rect 288495 248890 288640 248892
rect 288495 248834 288500 248890
rect 288556 248834 288640 248890
rect 288495 248832 288640 248834
rect 283136 248830 283185 248832
rect 283119 248829 283185 248830
rect 288495 248829 288561 248832
rect 288634 248830 288640 248832
rect 288704 248830 288710 248894
rect 288207 248744 288273 248747
rect 288634 248744 288640 248746
rect 288207 248742 288640 248744
rect 288207 248686 288212 248742
rect 288268 248686 288640 248742
rect 288207 248684 288640 248686
rect 288207 248681 288273 248684
rect 288634 248682 288640 248684
rect 288704 248682 288710 248746
rect 284794 248534 284800 248598
rect 284864 248596 284870 248598
rect 284864 248536 288288 248596
rect 284864 248534 284870 248536
rect 42063 248446 42174 248451
rect 42063 248390 42068 248446
rect 42124 248390 42174 248446
rect 42063 248388 42174 248390
rect 42063 248385 42129 248388
rect 284026 248386 284032 248450
rect 284096 248448 284102 248450
rect 284794 248448 284800 248450
rect 284096 248388 284800 248448
rect 284096 248386 284102 248388
rect 284794 248386 284800 248388
rect 284864 248386 284870 248450
rect 288207 248300 288273 248303
rect 288495 248300 288561 248303
rect 288207 248298 288561 248300
rect 288207 248242 288212 248298
rect 288268 248242 288500 248298
rect 288556 248242 288561 248298
rect 288207 248240 288561 248242
rect 288207 248237 288273 248240
rect 288495 248237 288561 248240
rect 43023 248152 43089 248155
rect 144015 248152 144081 248155
rect 42336 248150 43089 248152
rect 42336 248094 43028 248150
rect 43084 248094 43089 248150
rect 42336 248092 43089 248094
rect 140832 248150 144081 248152
rect 140832 248094 144020 248150
rect 144076 248094 144081 248150
rect 140832 248092 144081 248094
rect 43023 248089 43089 248092
rect 144015 248089 144081 248092
rect 285754 248090 285760 248154
rect 285824 248152 285830 248154
rect 285903 248152 285969 248155
rect 285824 248150 285969 248152
rect 285824 248094 285908 248150
rect 285964 248094 285969 248150
rect 285824 248092 285969 248094
rect 285824 248090 285830 248092
rect 285903 248089 285969 248092
rect 284986 247942 284992 248006
rect 285056 248004 285062 248006
rect 285056 247944 288288 248004
rect 285056 247942 285062 247944
rect 40570 247794 40576 247858
rect 40640 247794 40646 247858
rect 40578 247708 40638 247794
rect 41530 247708 41536 247710
rect 40578 247648 41536 247708
rect 41530 247646 41536 247648
rect 41600 247646 41606 247710
rect 34626 247119 34686 247382
rect 284794 247350 284800 247414
rect 284864 247412 284870 247414
rect 284864 247352 288288 247412
rect 284864 247350 284870 247352
rect 285807 247266 285873 247267
rect 285754 247264 285760 247266
rect 285716 247204 285760 247264
rect 285824 247262 285873 247266
rect 285868 247206 285873 247262
rect 285754 247202 285760 247204
rect 285824 247202 285873 247206
rect 285807 247201 285873 247202
rect 34575 247114 34686 247119
rect 34575 247058 34580 247114
rect 34636 247058 34686 247114
rect 34575 247056 34686 247058
rect 34575 247053 34641 247056
rect 284410 246906 284416 246970
rect 284480 246968 284486 246970
rect 284480 246908 288288 246968
rect 284480 246906 284486 246908
rect 140802 246376 140862 246864
rect 288634 246610 288640 246674
rect 288704 246610 288710 246674
rect 144111 246376 144177 246379
rect 140802 246374 144177 246376
rect 140802 246318 144116 246374
rect 144172 246318 144177 246374
rect 288642 246346 288702 246610
rect 140802 246316 144177 246318
rect 144111 246313 144177 246316
rect 34575 246080 34641 246083
rect 34575 246078 34686 246080
rect 34575 246022 34580 246078
rect 34636 246022 34686 246078
rect 34575 246017 34686 246022
rect 34626 245902 34686 246017
rect 284218 245722 284224 245786
rect 284288 245784 284294 245786
rect 284288 245724 288288 245784
rect 284288 245722 284294 245724
rect 140802 245340 140862 245670
rect 144015 245340 144081 245343
rect 140802 245338 144081 245340
rect 140802 245282 144020 245338
rect 144076 245282 144081 245338
rect 140802 245280 144081 245282
rect 144015 245277 144081 245280
rect 282351 245340 282417 245343
rect 282351 245338 288288 245340
rect 282351 245282 282356 245338
rect 282412 245282 288288 245338
rect 282351 245280 288288 245282
rect 282351 245277 282417 245280
rect 675279 245046 675345 245047
rect 674938 244982 674944 245046
rect 675008 245044 675014 245046
rect 675279 245044 675328 245046
rect 675008 245042 675328 245044
rect 675008 244986 675284 245042
rect 675008 244984 675328 244986
rect 675008 244982 675014 244984
rect 675279 244982 675328 244984
rect 675392 244982 675398 245046
rect 675279 244981 675345 244982
rect 282255 244748 282321 244751
rect 675471 244750 675537 244751
rect 675471 244748 675520 244750
rect 282255 244746 288288 244748
rect 282255 244690 282260 244746
rect 282316 244690 288288 244746
rect 282255 244688 288288 244690
rect 675428 244746 675520 244748
rect 675428 244690 675476 244746
rect 675428 244688 675520 244690
rect 282255 244685 282321 244688
rect 675471 244686 675520 244688
rect 675584 244686 675590 244750
rect 675471 244685 675537 244686
rect 145594 244452 145600 244454
rect 140832 244392 145600 244452
rect 145594 244390 145600 244392
rect 145664 244390 145670 244454
rect 284271 244156 284337 244159
rect 284271 244154 288288 244156
rect 284271 244098 284276 244154
rect 284332 244098 288288 244154
rect 284271 244096 288288 244098
rect 284271 244093 284337 244096
rect 282255 243712 282321 243715
rect 282255 243710 288288 243712
rect 282255 243654 282260 243710
rect 282316 243654 288288 243710
rect 282255 243652 288288 243654
rect 282255 243649 282321 243652
rect 674554 243502 674560 243566
rect 674624 243564 674630 243566
rect 675471 243564 675537 243567
rect 674624 243562 675537 243564
rect 674624 243506 675476 243562
rect 675532 243506 675537 243562
rect 674624 243504 675537 243506
rect 674624 243502 674630 243504
rect 675471 243501 675537 243504
rect 140802 242824 140862 243312
rect 283023 243120 283089 243123
rect 283023 243118 288288 243120
rect 283023 243062 283028 243118
rect 283084 243062 288288 243118
rect 283023 243060 288288 243062
rect 283023 243057 283089 243060
rect 144015 242824 144081 242827
rect 140802 242822 144081 242824
rect 140802 242766 144020 242822
rect 144076 242766 144081 242822
rect 140802 242764 144081 242766
rect 144015 242761 144081 242764
rect 282447 242528 282513 242531
rect 282447 242526 288288 242528
rect 282447 242470 282452 242526
rect 282508 242470 288288 242526
rect 282447 242468 288288 242470
rect 282447 242465 282513 242468
rect 282351 242380 282417 242383
rect 282351 242378 288318 242380
rect 282351 242322 282356 242378
rect 282412 242322 288318 242378
rect 282351 242320 288318 242322
rect 282351 242317 282417 242320
rect 286522 242170 286528 242234
rect 286592 242232 286598 242234
rect 288015 242232 288081 242235
rect 286592 242230 288081 242232
rect 286592 242174 288020 242230
rect 288076 242174 288081 242230
rect 286592 242172 288081 242174
rect 286592 242170 286598 242172
rect 288015 242169 288081 242172
rect 140802 242084 140862 242128
rect 145743 242084 145809 242087
rect 140802 242082 145809 242084
rect 140802 242026 145748 242082
rect 145804 242026 145809 242082
rect 140802 242024 145809 242026
rect 145743 242021 145809 242024
rect 288258 241980 288318 242320
rect 288399 242232 288465 242235
rect 288634 242232 288640 242234
rect 288399 242230 288640 242232
rect 288399 242174 288404 242230
rect 288460 242174 288640 242230
rect 288399 242172 288640 242174
rect 288399 242169 288465 242172
rect 288634 242170 288640 242172
rect 288704 242170 288710 242234
rect 284943 241492 285009 241495
rect 284943 241490 288288 241492
rect 284943 241434 284948 241490
rect 285004 241434 288288 241490
rect 284943 241432 288288 241434
rect 284943 241429 285009 241432
rect 145786 240900 145792 240902
rect 140832 240840 145792 240900
rect 145786 240838 145792 240840
rect 145856 240838 145862 240902
rect 42298 240690 42304 240754
rect 42368 240752 42374 240754
rect 42639 240752 42705 240755
rect 42368 240750 42705 240752
rect 42368 240694 42644 240750
rect 42700 240694 42705 240750
rect 42368 240692 42705 240694
rect 42368 240690 42374 240692
rect 42639 240689 42705 240692
rect 288450 240311 288510 240870
rect 288399 240306 288510 240311
rect 288399 240250 288404 240306
rect 288460 240250 288510 240306
rect 288399 240248 288510 240250
rect 288399 240245 288465 240248
rect 140802 239124 140862 239658
rect 290178 239656 294078 239716
rect 287482 239506 287488 239570
rect 287552 239568 287558 239570
rect 288975 239568 289041 239571
rect 287552 239566 289041 239568
rect 287552 239510 288980 239566
rect 289036 239510 289041 239566
rect 287552 239508 289041 239510
rect 287552 239506 287558 239508
rect 288975 239505 289041 239508
rect 289402 239506 289408 239570
rect 289472 239568 289478 239570
rect 289743 239568 289809 239571
rect 290178 239570 290238 239656
rect 290895 239570 290961 239571
rect 291183 239570 291249 239571
rect 291375 239570 291441 239571
rect 289472 239566 289809 239568
rect 289472 239510 289748 239566
rect 289804 239510 289809 239566
rect 289472 239508 289809 239510
rect 289472 239506 289478 239508
rect 289743 239505 289809 239508
rect 290170 239506 290176 239570
rect 290240 239506 290246 239570
rect 290895 239568 290944 239570
rect 290852 239566 290944 239568
rect 290852 239510 290900 239566
rect 290852 239508 290944 239510
rect 290895 239506 290944 239508
rect 291008 239506 291014 239570
rect 291130 239568 291136 239570
rect 291092 239508 291136 239568
rect 291200 239566 291249 239570
rect 291244 239510 291249 239566
rect 291130 239506 291136 239508
rect 291200 239506 291249 239510
rect 291322 239506 291328 239570
rect 291392 239568 291441 239570
rect 291567 239568 291633 239571
rect 291951 239570 292017 239571
rect 292335 239570 292401 239571
rect 292719 239570 292785 239571
rect 293103 239570 293169 239571
rect 291706 239568 291712 239570
rect 291392 239566 291484 239568
rect 291436 239510 291484 239566
rect 291392 239508 291484 239510
rect 291567 239566 291712 239568
rect 291567 239510 291572 239566
rect 291628 239510 291712 239566
rect 291567 239508 291712 239510
rect 291392 239506 291441 239508
rect 290895 239505 290961 239506
rect 291183 239505 291249 239506
rect 291375 239505 291441 239506
rect 291567 239505 291633 239508
rect 291706 239506 291712 239508
rect 291776 239506 291782 239570
rect 291898 239506 291904 239570
rect 291968 239568 292017 239570
rect 291968 239566 292060 239568
rect 292012 239510 292060 239566
rect 291968 239508 292060 239510
rect 291968 239506 292017 239508
rect 292282 239506 292288 239570
rect 292352 239568 292401 239570
rect 292352 239566 292444 239568
rect 292396 239510 292444 239566
rect 292352 239508 292444 239510
rect 292352 239506 292401 239508
rect 292666 239506 292672 239570
rect 292736 239568 292785 239570
rect 292736 239566 292828 239568
rect 292780 239510 292828 239566
rect 292736 239508 292828 239510
rect 292736 239506 292785 239508
rect 293050 239506 293056 239570
rect 293120 239568 293169 239570
rect 294018 239568 294078 239656
rect 385554 239656 398718 239716
rect 385554 239571 385614 239656
rect 294927 239568 294993 239571
rect 293120 239566 293212 239568
rect 293164 239510 293212 239566
rect 293120 239508 293212 239510
rect 294018 239566 294993 239568
rect 294018 239510 294932 239566
rect 294988 239510 294993 239566
rect 294018 239508 294993 239510
rect 293120 239506 293169 239508
rect 291951 239505 292017 239506
rect 292335 239505 292401 239506
rect 292719 239505 292785 239506
rect 293103 239505 293169 239506
rect 294927 239505 294993 239508
rect 385551 239566 385617 239571
rect 385551 239510 385556 239566
rect 385612 239510 385617 239566
rect 385551 239505 385617 239510
rect 288634 239358 288640 239422
rect 288704 239420 288710 239422
rect 289551 239420 289617 239423
rect 288704 239418 289617 239420
rect 288704 239362 289556 239418
rect 289612 239362 289617 239418
rect 288704 239360 289617 239362
rect 288704 239358 288710 239360
rect 289551 239357 289617 239360
rect 290746 239358 290752 239422
rect 290816 239420 290822 239422
rect 293103 239420 293169 239423
rect 290816 239418 293169 239420
rect 290816 239362 293108 239418
rect 293164 239362 293169 239418
rect 290816 239360 293169 239362
rect 290816 239358 290822 239360
rect 293103 239357 293169 239360
rect 293242 239358 293248 239422
rect 293312 239420 293318 239422
rect 293391 239420 293457 239423
rect 293312 239418 293457 239420
rect 293312 239362 293396 239418
rect 293452 239362 293457 239418
rect 293312 239360 293457 239362
rect 398658 239420 398718 239656
rect 408258 239656 411822 239716
rect 408258 239420 408318 239656
rect 411762 239571 411822 239656
rect 437775 239605 437841 239608
rect 437634 239603 437841 239605
rect 408879 239568 408945 239571
rect 410703 239568 410769 239571
rect 408879 239566 410769 239568
rect 408879 239510 408884 239566
rect 408940 239510 410708 239566
rect 410764 239510 410769 239566
rect 408879 239508 410769 239510
rect 408879 239505 408945 239508
rect 410703 239505 410769 239508
rect 411759 239566 411825 239571
rect 411759 239510 411764 239566
rect 411820 239510 411825 239566
rect 411759 239505 411825 239510
rect 437634 239547 437780 239603
rect 437836 239547 437841 239603
rect 437634 239545 437841 239547
rect 398658 239360 408318 239420
rect 408879 239420 408945 239423
rect 415503 239420 415569 239423
rect 408879 239418 415569 239420
rect 408879 239362 408884 239418
rect 408940 239362 415508 239418
rect 415564 239362 415569 239418
rect 408879 239360 415569 239362
rect 293312 239358 293318 239360
rect 293391 239357 293457 239360
rect 408879 239357 408945 239360
rect 415503 239357 415569 239360
rect 421935 239420 422001 239423
rect 437634 239420 437694 239545
rect 437775 239542 437841 239545
rect 442618 239506 442624 239570
rect 442688 239506 442694 239570
rect 443727 239568 443793 239571
rect 446266 239568 446272 239570
rect 443727 239566 446272 239568
rect 443727 239510 443732 239566
rect 443788 239510 446272 239566
rect 443727 239508 446272 239510
rect 442626 239423 442686 239506
rect 443727 239505 443793 239508
rect 446266 239506 446272 239508
rect 446336 239506 446342 239570
rect 421935 239418 437694 239420
rect 421935 239362 421940 239418
rect 421996 239362 437694 239418
rect 421935 239360 437694 239362
rect 421935 239357 422001 239360
rect 441082 239358 441088 239422
rect 441152 239420 441158 239422
rect 442426 239420 442432 239422
rect 441152 239360 442432 239420
rect 441152 239358 441158 239360
rect 442426 239358 442432 239360
rect 442496 239358 442502 239422
rect 442626 239418 442737 239423
rect 442626 239362 442676 239418
rect 442732 239362 442737 239418
rect 442626 239360 442737 239362
rect 442671 239357 442737 239360
rect 443535 239420 443601 239423
rect 444303 239422 444369 239423
rect 445263 239422 445329 239423
rect 443962 239420 443968 239422
rect 443535 239418 443968 239420
rect 443535 239362 443540 239418
rect 443596 239362 443968 239418
rect 443535 239360 443968 239362
rect 443535 239357 443601 239360
rect 443962 239358 443968 239360
rect 444032 239358 444038 239422
rect 444303 239420 444352 239422
rect 444260 239418 444352 239420
rect 444260 239362 444308 239418
rect 444260 239360 444352 239362
rect 444303 239358 444352 239360
rect 444416 239358 444422 239422
rect 445263 239420 445312 239422
rect 445220 239418 445312 239420
rect 445220 239362 445268 239418
rect 445220 239360 445312 239362
rect 445263 239358 445312 239360
rect 445376 239358 445382 239422
rect 446607 239420 446673 239423
rect 447802 239420 447808 239422
rect 446607 239418 447808 239420
rect 446607 239362 446612 239418
rect 446668 239362 447808 239418
rect 446607 239360 447808 239362
rect 444303 239357 444369 239358
rect 445263 239357 445329 239358
rect 446607 239357 446673 239360
rect 447802 239358 447808 239360
rect 447872 239358 447878 239422
rect 447951 239420 448017 239423
rect 450106 239420 450112 239422
rect 447951 239418 450112 239420
rect 447951 239362 447956 239418
rect 448012 239362 450112 239418
rect 447951 239360 450112 239362
rect 447951 239357 448017 239360
rect 450106 239358 450112 239360
rect 450176 239358 450182 239422
rect 292858 239210 292864 239274
rect 292928 239272 292934 239274
rect 297807 239272 297873 239275
rect 292928 239270 297873 239272
rect 292928 239214 297812 239270
rect 297868 239214 297873 239270
rect 292928 239212 297873 239214
rect 292928 239210 292934 239212
rect 297807 239209 297873 239212
rect 398511 239272 398577 239275
rect 444111 239274 444177 239275
rect 443578 239272 443584 239274
rect 398511 239270 443584 239272
rect 398511 239214 398516 239270
rect 398572 239214 443584 239270
rect 398511 239212 443584 239214
rect 398511 239209 398577 239212
rect 443578 239210 443584 239212
rect 443648 239210 443654 239274
rect 444111 239272 444160 239274
rect 444068 239270 444160 239272
rect 444068 239214 444116 239270
rect 444068 239212 444160 239214
rect 444111 239210 444160 239212
rect 444224 239210 444230 239274
rect 444399 239272 444465 239275
rect 445114 239272 445120 239274
rect 444399 239270 445120 239272
rect 444399 239214 444404 239270
rect 444460 239214 445120 239270
rect 444399 239212 445120 239214
rect 444111 239209 444177 239210
rect 444399 239209 444465 239212
rect 445114 239210 445120 239212
rect 445184 239210 445190 239274
rect 446703 239272 446769 239275
rect 447610 239272 447616 239274
rect 446703 239270 447616 239272
rect 446703 239214 446708 239270
rect 446764 239214 447616 239270
rect 446703 239212 447616 239214
rect 446703 239209 446769 239212
rect 447610 239210 447616 239212
rect 447680 239210 447686 239274
rect 448143 239272 448209 239275
rect 448762 239272 448768 239274
rect 448143 239270 448768 239272
rect 448143 239214 448148 239270
rect 448204 239214 448768 239270
rect 448143 239212 448768 239214
rect 448143 239209 448209 239212
rect 448762 239210 448768 239212
rect 448832 239210 448838 239274
rect 144015 239124 144081 239127
rect 140802 239122 144081 239124
rect 140802 239066 144020 239122
rect 144076 239066 144081 239122
rect 140802 239064 144081 239066
rect 144015 239061 144081 239064
rect 290554 239062 290560 239126
rect 290624 239124 290630 239126
rect 293775 239124 293841 239127
rect 290624 239122 293841 239124
rect 290624 239066 293780 239122
rect 293836 239066 293841 239122
rect 290624 239064 293841 239066
rect 290624 239062 290630 239064
rect 293775 239061 293841 239064
rect 389871 239124 389937 239127
rect 450298 239124 450304 239126
rect 389871 239122 450304 239124
rect 389871 239066 389876 239122
rect 389932 239066 450304 239122
rect 389871 239064 450304 239066
rect 389871 239061 389937 239064
rect 450298 239062 450304 239064
rect 450368 239062 450374 239126
rect 291514 238914 291520 238978
rect 291584 238976 291590 238978
rect 295983 238976 296049 238979
rect 291584 238974 296049 238976
rect 291584 238918 295988 238974
rect 296044 238918 296049 238974
rect 291584 238916 296049 238918
rect 291584 238914 291590 238916
rect 295983 238913 296049 238916
rect 297999 238976 298065 238979
rect 341679 238976 341745 238979
rect 297999 238974 341745 238976
rect 297999 238918 298004 238974
rect 298060 238918 341684 238974
rect 341740 238918 341745 238974
rect 297999 238916 341745 238918
rect 297999 238913 298065 238916
rect 341679 238913 341745 238916
rect 390639 238976 390705 238979
rect 442234 238976 442240 238978
rect 390639 238974 442240 238976
rect 390639 238918 390644 238974
rect 390700 238918 442240 238974
rect 390639 238916 442240 238918
rect 390639 238913 390705 238916
rect 442234 238914 442240 238916
rect 442304 238914 442310 238978
rect 442426 238914 442432 238978
rect 442496 238976 442502 238978
rect 445882 238976 445888 238978
rect 442496 238916 445888 238976
rect 442496 238914 442502 238916
rect 445882 238914 445888 238916
rect 445952 238914 445958 238978
rect 674746 238914 674752 238978
rect 674816 238976 674822 238978
rect 675087 238976 675153 238979
rect 674816 238974 675153 238976
rect 674816 238918 675092 238974
rect 675148 238918 675153 238974
rect 674816 238916 675153 238918
rect 674816 238914 674822 238916
rect 675087 238913 675153 238916
rect 212943 238828 213009 238831
rect 388335 238828 388401 238831
rect 212943 238826 388401 238828
rect 212943 238770 212948 238826
rect 213004 238770 388340 238826
rect 388396 238770 388401 238826
rect 212943 238768 388401 238770
rect 212943 238765 213009 238768
rect 388335 238765 388401 238768
rect 392079 238828 392145 238831
rect 442042 238828 442048 238830
rect 392079 238826 442048 238828
rect 392079 238770 392084 238826
rect 392140 238770 442048 238826
rect 392079 238768 442048 238770
rect 392079 238765 392145 238768
rect 442042 238766 442048 238768
rect 442112 238766 442118 238830
rect 442618 238766 442624 238830
rect 442688 238828 442694 238830
rect 448954 238828 448960 238830
rect 442688 238768 448960 238828
rect 442688 238766 442694 238768
rect 448954 238766 448960 238768
rect 449024 238766 449030 238830
rect 287866 238618 287872 238682
rect 287936 238680 287942 238682
rect 297999 238680 298065 238683
rect 287936 238678 298065 238680
rect 287936 238622 298004 238678
rect 298060 238622 298065 238678
rect 287936 238620 298065 238622
rect 287936 238618 287942 238620
rect 297999 238617 298065 238620
rect 342447 238680 342513 238683
rect 675663 238682 675729 238683
rect 447034 238680 447040 238682
rect 342447 238678 447040 238680
rect 342447 238622 342452 238678
rect 342508 238622 447040 238678
rect 342447 238620 447040 238622
rect 342447 238617 342513 238620
rect 447034 238618 447040 238620
rect 447104 238618 447110 238682
rect 675663 238678 675712 238682
rect 675776 238680 675782 238682
rect 675663 238622 675668 238678
rect 675663 238618 675712 238622
rect 675776 238620 675820 238680
rect 675776 238618 675782 238620
rect 675663 238617 675729 238618
rect 221487 238532 221553 238535
rect 392463 238532 392529 238535
rect 221487 238530 392529 238532
rect 221487 238474 221492 238530
rect 221548 238474 392468 238530
rect 392524 238474 392529 238530
rect 221487 238472 392529 238474
rect 221487 238469 221553 238472
rect 392463 238469 392529 238472
rect 392655 238532 392721 238535
rect 392655 238530 400446 238532
rect 392655 238474 392660 238530
rect 392716 238474 400446 238530
rect 392655 238472 400446 238474
rect 392655 238469 392721 238472
rect 140802 237940 140862 238428
rect 227439 238384 227505 238387
rect 396495 238384 396561 238387
rect 227439 238382 396561 238384
rect 227439 238326 227444 238382
rect 227500 238326 396500 238382
rect 396556 238326 396561 238382
rect 227439 238324 396561 238326
rect 400386 238384 400446 238472
rect 400570 238470 400576 238534
rect 400640 238532 400646 238534
rect 447226 238532 447232 238534
rect 400640 238472 447232 238532
rect 400640 238470 400646 238472
rect 447226 238470 447232 238472
rect 447296 238470 447302 238534
rect 445690 238384 445696 238386
rect 400386 238324 445696 238384
rect 227439 238321 227505 238324
rect 396495 238321 396561 238324
rect 445690 238322 445696 238324
rect 445760 238322 445766 238386
rect 292090 238174 292096 238238
rect 292160 238236 292166 238238
rect 305103 238236 305169 238239
rect 292160 238234 305169 238236
rect 292160 238178 305108 238234
rect 305164 238178 305169 238234
rect 292160 238176 305169 238178
rect 292160 238174 292166 238176
rect 305103 238173 305169 238176
rect 345615 238236 345681 238239
rect 345903 238236 345969 238239
rect 345615 238234 345969 238236
rect 345615 238178 345620 238234
rect 345676 238178 345908 238234
rect 345964 238178 345969 238234
rect 345615 238176 345969 238178
rect 345615 238173 345681 238176
rect 345903 238173 345969 238176
rect 347535 238236 347601 238239
rect 512847 238236 512913 238239
rect 347535 238234 512913 238236
rect 347535 238178 347540 238234
rect 347596 238178 512852 238234
rect 512908 238178 512913 238234
rect 347535 238176 512913 238178
rect 347535 238173 347601 238176
rect 512847 238173 512913 238176
rect 347151 238088 347217 238091
rect 509871 238088 509937 238091
rect 347151 238086 509937 238088
rect 347151 238030 347156 238086
rect 347212 238030 509876 238086
rect 509932 238030 509937 238086
rect 347151 238028 509937 238030
rect 347151 238025 347217 238028
rect 509871 238025 509937 238028
rect 144015 237940 144081 237943
rect 140802 237938 144081 237940
rect 140802 237882 144020 237938
rect 144076 237882 144081 237938
rect 140802 237880 144081 237882
rect 144015 237877 144081 237880
rect 301551 237940 301617 237943
rect 406095 237940 406161 237943
rect 301551 237938 406161 237940
rect 301551 237882 301556 237938
rect 301612 237882 406100 237938
rect 406156 237882 406161 237938
rect 301551 237880 406161 237882
rect 301551 237877 301617 237880
rect 406095 237877 406161 237880
rect 411759 237940 411825 237943
rect 421935 237940 422001 237943
rect 411759 237938 422001 237940
rect 411759 237882 411764 237938
rect 411820 237882 421940 237938
rect 421996 237882 422001 237938
rect 411759 237880 422001 237882
rect 411759 237877 411825 237880
rect 421935 237877 422001 237880
rect 435279 237940 435345 237943
rect 445498 237940 445504 237942
rect 435279 237938 445504 237940
rect 435279 237882 435284 237938
rect 435340 237882 445504 237938
rect 435279 237880 445504 237882
rect 435279 237877 435345 237880
rect 445498 237878 445504 237880
rect 445568 237878 445574 237942
rect 325551 237792 325617 237795
rect 325935 237792 326001 237795
rect 325551 237790 326001 237792
rect 325551 237734 325556 237790
rect 325612 237734 325940 237790
rect 325996 237734 326001 237790
rect 325551 237732 326001 237734
rect 325551 237729 325617 237732
rect 325935 237729 326001 237732
rect 343887 237792 343953 237795
rect 450682 237792 450688 237794
rect 343887 237790 450688 237792
rect 343887 237734 343892 237790
rect 343948 237734 450688 237790
rect 343887 237732 450688 237734
rect 343887 237729 343953 237732
rect 450682 237730 450688 237732
rect 450752 237730 450758 237794
rect 293434 237582 293440 237646
rect 293504 237644 293510 237646
rect 396303 237644 396369 237647
rect 293504 237642 396369 237644
rect 293504 237586 396308 237642
rect 396364 237586 396369 237642
rect 293504 237584 396369 237586
rect 293504 237582 293510 237584
rect 396303 237581 396369 237584
rect 396495 237644 396561 237647
rect 411279 237644 411345 237647
rect 396495 237642 411345 237644
rect 396495 237586 396500 237642
rect 396556 237586 411284 237642
rect 411340 237586 411345 237642
rect 396495 237584 411345 237586
rect 396495 237581 396561 237584
rect 411279 237581 411345 237584
rect 413967 237644 414033 237647
rect 446650 237644 446656 237646
rect 413967 237642 446656 237644
rect 413967 237586 413972 237642
rect 414028 237586 446656 237642
rect 413967 237584 446656 237586
rect 413967 237581 414033 237584
rect 446650 237582 446656 237584
rect 446720 237582 446726 237646
rect 447226 237582 447232 237646
rect 447296 237644 447302 237646
rect 448186 237644 448192 237646
rect 447296 237584 448192 237644
rect 447296 237582 447302 237584
rect 448186 237582 448192 237584
rect 448256 237582 448262 237646
rect 301167 237496 301233 237499
rect 403215 237496 403281 237499
rect 301167 237494 403281 237496
rect 301167 237438 301172 237494
rect 301228 237438 403220 237494
rect 403276 237438 403281 237494
rect 301167 237436 403281 237438
rect 301167 237433 301233 237436
rect 403215 237433 403281 237436
rect 408207 237496 408273 237499
rect 444538 237496 444544 237498
rect 408207 237494 444544 237496
rect 408207 237438 408212 237494
rect 408268 237438 444544 237494
rect 408207 237436 444544 237438
rect 408207 237433 408273 237436
rect 444538 237434 444544 237436
rect 444608 237434 444614 237498
rect 286906 237286 286912 237350
rect 286976 237348 286982 237350
rect 353679 237348 353745 237351
rect 286976 237346 353745 237348
rect 286976 237290 353684 237346
rect 353740 237290 353745 237346
rect 286976 237288 353745 237290
rect 286976 237286 286982 237288
rect 353679 237285 353745 237288
rect 385167 237348 385233 237351
rect 398799 237348 398865 237351
rect 441658 237348 441664 237350
rect 385167 237346 390078 237348
rect 385167 237290 385172 237346
rect 385228 237290 390078 237346
rect 385167 237288 390078 237290
rect 385167 237285 385233 237288
rect 140802 236756 140862 237238
rect 300495 237200 300561 237203
rect 354543 237200 354609 237203
rect 300495 237198 354609 237200
rect 300495 237142 300500 237198
rect 300556 237142 354548 237198
rect 354604 237142 354609 237198
rect 300495 237140 354609 237142
rect 390018 237200 390078 237288
rect 398799 237346 441664 237348
rect 398799 237290 398804 237346
rect 398860 237290 441664 237346
rect 398799 237288 441664 237290
rect 398799 237285 398865 237288
rect 441658 237286 441664 237288
rect 441728 237286 441734 237350
rect 442671 237348 442737 237351
rect 442810 237348 442816 237350
rect 442671 237346 442816 237348
rect 442671 237290 442676 237346
rect 442732 237290 442816 237346
rect 442671 237288 442816 237290
rect 442671 237285 442737 237288
rect 442810 237286 442816 237288
rect 442880 237286 442886 237350
rect 449914 237200 449920 237202
rect 390018 237140 449920 237200
rect 300495 237137 300561 237140
rect 354543 237137 354609 237140
rect 449914 237138 449920 237140
rect 449984 237138 449990 237202
rect 301935 237052 302001 237055
rect 357039 237052 357105 237055
rect 301935 237050 357105 237052
rect 301935 236994 301940 237050
rect 301996 236994 357044 237050
rect 357100 236994 357105 237050
rect 301935 236992 357105 236994
rect 301935 236989 302001 236992
rect 357039 236989 357105 236992
rect 383343 237052 383409 237055
rect 398799 237052 398865 237055
rect 399183 237054 399249 237055
rect 399183 237052 399232 237054
rect 383343 237050 398865 237052
rect 383343 236994 383348 237050
rect 383404 236994 398804 237050
rect 398860 236994 398865 237050
rect 383343 236992 398865 236994
rect 399140 237050 399232 237052
rect 399140 236994 399188 237050
rect 399140 236992 399232 236994
rect 383343 236989 383409 236992
rect 398799 236989 398865 236992
rect 399183 236990 399232 236992
rect 399296 236990 399302 237054
rect 399375 237052 399441 237055
rect 446074 237052 446080 237054
rect 399375 237050 446080 237052
rect 399375 236994 399380 237050
rect 399436 236994 446080 237050
rect 399375 236992 446080 236994
rect 399183 236989 399249 236990
rect 399375 236989 399441 236992
rect 446074 236990 446080 236992
rect 446144 236990 446150 237054
rect 300783 236904 300849 236907
rect 354831 236904 354897 236907
rect 300783 236902 354897 236904
rect 300783 236846 300788 236902
rect 300844 236846 354836 236902
rect 354892 236846 354897 236902
rect 300783 236844 354897 236846
rect 300783 236841 300849 236844
rect 354831 236841 354897 236844
rect 389487 236904 389553 236907
rect 400570 236904 400576 236906
rect 389487 236902 400576 236904
rect 389487 236846 389492 236902
rect 389548 236846 400576 236902
rect 389487 236844 400576 236846
rect 389487 236841 389553 236844
rect 400570 236842 400576 236844
rect 400640 236842 400646 236906
rect 404463 236904 404529 236907
rect 408783 236904 408849 236907
rect 404463 236902 408849 236904
rect 404463 236846 404468 236902
rect 404524 236846 408788 236902
rect 408844 236846 408849 236902
rect 404463 236844 408849 236846
rect 404463 236841 404529 236844
rect 408783 236841 408849 236844
rect 411322 236842 411328 236906
rect 411392 236904 411398 236906
rect 444730 236904 444736 236906
rect 411392 236844 444736 236904
rect 411392 236842 411398 236844
rect 444730 236842 444736 236844
rect 444800 236842 444806 236906
rect 674362 236842 674368 236906
rect 674432 236904 674438 236906
rect 675375 236904 675441 236907
rect 674432 236902 675441 236904
rect 674432 236846 675380 236902
rect 675436 236846 675441 236902
rect 674432 236844 675441 236846
rect 674432 236842 674438 236844
rect 675375 236841 675441 236844
rect 145978 236756 145984 236758
rect 140802 236696 145984 236756
rect 145978 236694 145984 236696
rect 146048 236694 146054 236758
rect 300111 236756 300177 236759
rect 359151 236756 359217 236759
rect 300111 236754 359217 236756
rect 300111 236698 300116 236754
rect 300172 236698 359156 236754
rect 359212 236698 359217 236754
rect 300111 236696 359217 236698
rect 300111 236693 300177 236696
rect 359151 236693 359217 236696
rect 387951 236756 388017 236759
rect 442426 236756 442432 236758
rect 387951 236754 442432 236756
rect 387951 236698 387956 236754
rect 388012 236698 442432 236754
rect 387951 236696 442432 236698
rect 387951 236693 388017 236696
rect 442426 236694 442432 236696
rect 442496 236694 442502 236758
rect 299727 236608 299793 236611
rect 360495 236608 360561 236611
rect 299727 236606 360561 236608
rect 299727 236550 299732 236606
rect 299788 236550 360500 236606
rect 360556 236550 360561 236606
rect 299727 236548 360561 236550
rect 299727 236545 299793 236548
rect 360495 236545 360561 236548
rect 396303 236608 396369 236611
rect 406671 236608 406737 236611
rect 396303 236606 406737 236608
rect 396303 236550 396308 236606
rect 396364 236550 406676 236606
rect 406732 236550 406737 236606
rect 396303 236548 406737 236550
rect 396303 236545 396369 236548
rect 406671 236545 406737 236548
rect 406863 236608 406929 236611
rect 444922 236608 444928 236610
rect 406863 236606 444928 236608
rect 406863 236550 406868 236606
rect 406924 236550 444928 236606
rect 406863 236548 444928 236550
rect 406863 236545 406929 236548
rect 444922 236546 444928 236548
rect 444992 236546 444998 236610
rect 292474 236398 292480 236462
rect 292544 236460 292550 236462
rect 296559 236460 296625 236463
rect 292544 236458 296625 236460
rect 292544 236402 296564 236458
rect 296620 236402 296625 236458
rect 292544 236400 296625 236402
rect 292544 236398 292550 236400
rect 296559 236397 296625 236400
rect 298959 236460 299025 236463
rect 487023 236460 487089 236463
rect 298959 236458 487089 236460
rect 298959 236402 298964 236458
rect 299020 236402 487028 236458
rect 487084 236402 487089 236458
rect 298959 236400 487089 236402
rect 298959 236397 299025 236400
rect 487023 236397 487089 236400
rect 299343 236312 299409 236315
rect 492687 236312 492753 236315
rect 299343 236310 492753 236312
rect 299343 236254 299348 236310
rect 299404 236254 492692 236310
rect 492748 236254 492753 236310
rect 299343 236252 492753 236254
rect 299343 236249 299409 236252
rect 492687 236249 492753 236252
rect 145359 236164 145425 236167
rect 140832 236162 145425 236164
rect 140832 236106 145364 236162
rect 145420 236106 145425 236162
rect 140832 236104 145425 236106
rect 145359 236101 145425 236104
rect 290362 236102 290368 236166
rect 290432 236164 290438 236166
rect 295311 236164 295377 236167
rect 290432 236162 295377 236164
rect 290432 236106 295316 236162
rect 295372 236106 295377 236162
rect 290432 236104 295377 236106
rect 290432 236102 290438 236104
rect 295311 236101 295377 236104
rect 358191 236164 358257 236167
rect 405231 236164 405297 236167
rect 358191 236162 405297 236164
rect 358191 236106 358196 236162
rect 358252 236106 405236 236162
rect 405292 236106 405297 236162
rect 358191 236104 405297 236106
rect 358191 236101 358257 236104
rect 405231 236101 405297 236104
rect 405423 236164 405489 236167
rect 411759 236164 411825 236167
rect 405423 236162 411825 236164
rect 405423 236106 405428 236162
rect 405484 236106 411764 236162
rect 411820 236106 411825 236162
rect 405423 236104 411825 236106
rect 405423 236101 405489 236104
rect 411759 236101 411825 236104
rect 420111 236164 420177 236167
rect 420879 236164 420945 236167
rect 420111 236162 420945 236164
rect 420111 236106 420116 236162
rect 420172 236106 420884 236162
rect 420940 236106 420945 236162
rect 420111 236104 420945 236106
rect 420111 236101 420177 236104
rect 420879 236101 420945 236104
rect 424239 236164 424305 236167
rect 441423 236164 441489 236167
rect 443631 236166 443697 236167
rect 443578 236164 443584 236166
rect 424239 236162 441489 236164
rect 424239 236106 424244 236162
rect 424300 236106 441428 236162
rect 441484 236106 441489 236162
rect 424239 236104 441489 236106
rect 443540 236104 443584 236164
rect 443648 236162 443697 236166
rect 443692 236106 443697 236162
rect 424239 236101 424305 236104
rect 441423 236101 441489 236104
rect 443578 236102 443584 236104
rect 443648 236102 443697 236106
rect 443631 236101 443697 236102
rect 289594 235954 289600 236018
rect 289664 236016 289670 236018
rect 294543 236016 294609 236019
rect 289664 236014 294609 236016
rect 289664 235958 294548 236014
rect 294604 235958 294609 236014
rect 289664 235956 294609 235958
rect 289664 235954 289670 235956
rect 294543 235953 294609 235956
rect 338511 236016 338577 236019
rect 357039 236016 357105 236019
rect 338511 236014 357105 236016
rect 338511 235958 338516 236014
rect 338572 235958 357044 236014
rect 357100 235958 357105 236014
rect 338511 235956 357105 235958
rect 338511 235953 338577 235956
rect 357039 235953 357105 235956
rect 368559 236016 368625 236019
rect 486639 236016 486705 236019
rect 368559 236014 486705 236016
rect 368559 235958 368564 236014
rect 368620 235958 486644 236014
rect 486700 235958 486705 236014
rect 368559 235956 486705 235958
rect 368559 235953 368625 235956
rect 486639 235953 486705 235956
rect 289786 235806 289792 235870
rect 289856 235868 289862 235870
rect 295599 235868 295665 235871
rect 289856 235866 295665 235868
rect 289856 235810 295604 235866
rect 295660 235810 295665 235866
rect 289856 235808 295665 235810
rect 289856 235806 289862 235808
rect 295599 235805 295665 235808
rect 297519 235868 297585 235871
rect 342735 235868 342801 235871
rect 297519 235866 342801 235868
rect 297519 235810 297524 235866
rect 297580 235810 342740 235866
rect 342796 235810 342801 235866
rect 297519 235808 342801 235810
rect 297519 235805 297585 235808
rect 342735 235805 342801 235808
rect 360303 235868 360369 235871
rect 360687 235868 360753 235871
rect 360303 235866 360753 235868
rect 360303 235810 360308 235866
rect 360364 235810 360692 235866
rect 360748 235810 360753 235866
rect 360303 235808 360753 235810
rect 360303 235805 360369 235808
rect 360687 235805 360753 235808
rect 371343 235868 371409 235871
rect 488079 235868 488145 235871
rect 371343 235866 488145 235868
rect 371343 235810 371348 235866
rect 371404 235810 488084 235866
rect 488140 235810 488145 235866
rect 371343 235808 488145 235810
rect 371343 235805 371409 235808
rect 488079 235805 488145 235808
rect 289978 235658 289984 235722
rect 290048 235720 290054 235722
rect 296751 235720 296817 235723
rect 290048 235718 296817 235720
rect 290048 235662 296756 235718
rect 296812 235662 296817 235718
rect 290048 235660 296817 235662
rect 290048 235658 290054 235660
rect 296751 235657 296817 235660
rect 314799 235720 314865 235723
rect 358287 235720 358353 235723
rect 314799 235718 358353 235720
rect 314799 235662 314804 235718
rect 314860 235662 358292 235718
rect 358348 235662 358353 235718
rect 314799 235660 358353 235662
rect 314799 235657 314865 235660
rect 358287 235657 358353 235660
rect 360111 235720 360177 235723
rect 360495 235720 360561 235723
rect 360111 235718 360561 235720
rect 360111 235662 360116 235718
rect 360172 235662 360500 235718
rect 360556 235662 360561 235718
rect 360111 235660 360561 235662
rect 360111 235657 360177 235660
rect 360495 235657 360561 235660
rect 369999 235720 370065 235723
rect 487311 235720 487377 235723
rect 369999 235718 487377 235720
rect 369999 235662 370004 235718
rect 370060 235662 487316 235718
rect 487372 235662 487377 235718
rect 369999 235660 487377 235662
rect 369999 235657 370065 235660
rect 487311 235657 487377 235660
rect 289018 235510 289024 235574
rect 289088 235572 289094 235574
rect 296367 235572 296433 235575
rect 289088 235570 296433 235572
rect 289088 235514 296372 235570
rect 296428 235514 296433 235570
rect 289088 235512 296433 235514
rect 289088 235510 289094 235512
rect 296367 235509 296433 235512
rect 316239 235572 316305 235575
rect 362223 235572 362289 235575
rect 316239 235570 362289 235572
rect 316239 235514 316244 235570
rect 316300 235514 362228 235570
rect 362284 235514 362289 235570
rect 316239 235512 362289 235514
rect 316239 235509 316305 235512
rect 362223 235509 362289 235512
rect 367023 235572 367089 235575
rect 485871 235572 485937 235575
rect 367023 235570 485937 235572
rect 367023 235514 367028 235570
rect 367084 235514 485876 235570
rect 485932 235514 485937 235570
rect 367023 235512 485937 235514
rect 367023 235509 367089 235512
rect 485871 235509 485937 235512
rect 289210 235362 289216 235426
rect 289280 235424 289286 235426
rect 298575 235424 298641 235427
rect 289280 235422 298641 235424
rect 289280 235366 298580 235422
rect 298636 235366 298641 235422
rect 289280 235364 298641 235366
rect 289280 235362 289286 235364
rect 298575 235361 298641 235364
rect 315567 235424 315633 235427
rect 362415 235424 362481 235427
rect 315567 235422 362481 235424
rect 315567 235366 315572 235422
rect 315628 235366 362420 235422
rect 362476 235366 362481 235422
rect 315567 235364 362481 235366
rect 315567 235361 315633 235364
rect 362415 235361 362481 235364
rect 365391 235424 365457 235427
rect 485103 235424 485169 235427
rect 365391 235422 485169 235424
rect 365391 235366 365396 235422
rect 365452 235366 485108 235422
rect 485164 235366 485169 235422
rect 365391 235364 485169 235366
rect 365391 235361 365457 235364
rect 485103 235361 485169 235364
rect 313359 235276 313425 235279
rect 359439 235276 359505 235279
rect 313359 235274 359505 235276
rect 313359 235218 313364 235274
rect 313420 235218 359444 235274
rect 359500 235218 359505 235274
rect 313359 235216 359505 235218
rect 313359 235213 313425 235216
rect 359439 235213 359505 235216
rect 362607 235276 362673 235279
rect 483663 235276 483729 235279
rect 362607 235274 483729 235276
rect 362607 235218 362612 235274
rect 362668 235218 483668 235274
rect 483724 235218 483729 235274
rect 362607 235216 483729 235218
rect 362607 235213 362673 235216
rect 483663 235213 483729 235216
rect 287674 235066 287680 235130
rect 287744 235128 287750 235130
rect 297135 235128 297201 235131
rect 287744 235126 297201 235128
rect 287744 235070 297140 235126
rect 297196 235070 297201 235126
rect 287744 235068 297201 235070
rect 287744 235066 287750 235068
rect 297135 235065 297201 235068
rect 312591 235128 312657 235131
rect 358863 235128 358929 235131
rect 312591 235126 358929 235128
rect 312591 235070 312596 235126
rect 312652 235070 358868 235126
rect 358924 235070 358929 235126
rect 312591 235068 358929 235070
rect 312591 235065 312657 235068
rect 358863 235065 358929 235068
rect 364143 235128 364209 235131
rect 484431 235128 484497 235131
rect 364143 235126 484497 235128
rect 364143 235070 364148 235126
rect 364204 235070 484436 235126
rect 484492 235070 484497 235126
rect 364143 235068 484497 235070
rect 364143 235065 364209 235068
rect 484431 235065 484497 235068
rect 213039 234980 213105 234983
rect 341295 234980 341361 234983
rect 213039 234978 341361 234980
rect 213039 234922 213044 234978
rect 213100 234922 341300 234978
rect 341356 234922 341361 234978
rect 213039 234920 341361 234922
rect 213039 234917 213105 234920
rect 341295 234917 341361 234920
rect 356751 234980 356817 234983
rect 480687 234980 480753 234983
rect 356751 234978 480753 234980
rect 356751 234922 356756 234978
rect 356812 234922 480692 234978
rect 480748 234922 480753 234978
rect 356751 234920 480753 234922
rect 356751 234917 356817 234920
rect 480687 234917 480753 234920
rect 42159 234832 42225 234835
rect 42298 234832 42304 234834
rect 42159 234830 42304 234832
rect 42159 234774 42164 234830
rect 42220 234774 42304 234830
rect 42159 234772 42304 234774
rect 42159 234769 42225 234772
rect 42298 234770 42304 234772
rect 42368 234770 42374 234834
rect 140802 234388 140862 234876
rect 310383 234832 310449 234835
rect 348783 234832 348849 234835
rect 310383 234830 348849 234832
rect 310383 234774 310388 234830
rect 310444 234774 348788 234830
rect 348844 234774 348849 234830
rect 310383 234772 348849 234774
rect 310383 234769 310449 234772
rect 348783 234769 348849 234772
rect 355119 234832 355185 234835
rect 480015 234832 480081 234835
rect 355119 234830 480081 234832
rect 355119 234774 355124 234830
rect 355180 234774 480020 234830
rect 480076 234774 480081 234830
rect 355119 234772 480081 234774
rect 355119 234769 355185 234772
rect 480015 234769 480081 234772
rect 309615 234684 309681 234687
rect 351759 234684 351825 234687
rect 309615 234682 351825 234684
rect 309615 234626 309620 234682
rect 309676 234626 351764 234682
rect 351820 234626 351825 234682
rect 309615 234624 351825 234626
rect 309615 234621 309681 234624
rect 351759 234621 351825 234624
rect 357519 234684 357585 234687
rect 481071 234684 481137 234687
rect 357519 234682 481137 234684
rect 357519 234626 357524 234682
rect 357580 234626 481076 234682
rect 481132 234626 481137 234682
rect 357519 234624 481137 234626
rect 357519 234621 357585 234624
rect 481071 234621 481137 234624
rect 385071 234536 385137 234539
rect 499887 234536 499953 234539
rect 385071 234534 499953 234536
rect 385071 234478 385076 234534
rect 385132 234478 499892 234534
rect 499948 234478 499953 234534
rect 385071 234476 499953 234478
rect 385071 234473 385137 234476
rect 499887 234473 499953 234476
rect 144111 234388 144177 234391
rect 140802 234386 144177 234388
rect 140802 234330 144116 234386
rect 144172 234330 144177 234386
rect 140802 234328 144177 234330
rect 144111 234325 144177 234328
rect 385839 234388 385905 234391
rect 500655 234388 500721 234391
rect 385839 234386 500721 234388
rect 385839 234330 385844 234386
rect 385900 234330 500660 234386
rect 500716 234330 500721 234386
rect 385839 234328 500721 234330
rect 385839 234325 385905 234328
rect 500655 234325 500721 234328
rect 302703 234240 302769 234243
rect 399663 234240 399729 234243
rect 302703 234238 399729 234240
rect 302703 234182 302708 234238
rect 302764 234182 399668 234238
rect 399724 234182 399729 234238
rect 302703 234180 399729 234182
rect 302703 234177 302769 234180
rect 399663 234177 399729 234180
rect 400239 234240 400305 234243
rect 406095 234240 406161 234243
rect 400239 234238 406161 234240
rect 400239 234182 400244 234238
rect 400300 234182 406100 234238
rect 406156 234182 406161 234238
rect 400239 234180 406161 234182
rect 400239 234177 400305 234180
rect 406095 234177 406161 234180
rect 406287 234240 406353 234243
rect 411759 234240 411825 234243
rect 406287 234238 411825 234240
rect 406287 234182 406292 234238
rect 406348 234182 411764 234238
rect 411820 234182 411825 234238
rect 406287 234180 411825 234182
rect 406287 234177 406353 234180
rect 411759 234177 411825 234180
rect 412335 234240 412401 234243
rect 441082 234240 441088 234242
rect 412335 234238 441088 234240
rect 412335 234182 412340 234238
rect 412396 234182 441088 234238
rect 412335 234180 441088 234182
rect 412335 234177 412401 234180
rect 441082 234178 441088 234180
rect 441152 234178 441158 234242
rect 441519 234240 441585 234243
rect 535695 234240 535761 234243
rect 441519 234238 535761 234240
rect 441519 234182 441524 234238
rect 441580 234182 535700 234238
rect 535756 234182 535761 234238
rect 441519 234180 535761 234182
rect 441519 234177 441585 234180
rect 535695 234177 535761 234180
rect 363375 234092 363441 234095
rect 435375 234092 435441 234095
rect 363375 234090 435441 234092
rect 363375 234034 363380 234090
rect 363436 234034 435380 234090
rect 435436 234034 435441 234090
rect 363375 234032 435441 234034
rect 363375 234029 363441 234032
rect 435375 234029 435441 234032
rect 435567 234092 435633 234095
rect 495375 234092 495441 234095
rect 435567 234090 495441 234092
rect 435567 234034 435572 234090
rect 435628 234034 495380 234090
rect 495436 234034 495441 234090
rect 435567 234032 495441 234034
rect 435567 234029 435633 234032
rect 495375 234029 495441 234032
rect 359727 233944 359793 233947
rect 404463 233944 404529 233947
rect 359727 233942 404529 233944
rect 359727 233886 359732 233942
rect 359788 233886 404468 233942
rect 404524 233886 404529 233942
rect 359727 233884 404529 233886
rect 359727 233881 359793 233884
rect 404463 233881 404529 233884
rect 408399 233944 408465 233947
rect 409455 233944 409521 233947
rect 408399 233942 409521 233944
rect 408399 233886 408404 233942
rect 408460 233886 409460 233942
rect 409516 233886 409521 233942
rect 408399 233884 409521 233886
rect 408399 233881 408465 233884
rect 409455 233881 409521 233884
rect 414351 233944 414417 233947
rect 451258 233944 451264 233946
rect 414351 233942 451264 233944
rect 414351 233886 414356 233942
rect 414412 233886 451264 233942
rect 414351 233884 451264 233886
rect 414351 233881 414417 233884
rect 451258 233882 451264 233884
rect 451328 233882 451334 233946
rect 401871 233796 401937 233799
rect 407247 233796 407313 233799
rect 401871 233794 407313 233796
rect 401871 233738 401876 233794
rect 401932 233738 407252 233794
rect 407308 233738 407313 233794
rect 401871 233736 407313 233738
rect 401871 233733 401937 233736
rect 407247 233733 407313 233736
rect 416751 233796 416817 233799
rect 447994 233796 448000 233798
rect 416751 233794 448000 233796
rect 416751 233738 416756 233794
rect 416812 233738 448000 233794
rect 416751 233736 448000 233738
rect 416751 233733 416817 233736
rect 447994 233734 448000 233736
rect 448064 233734 448070 233798
rect 140802 233500 140862 233692
rect 358959 233648 359025 233651
rect 403311 233648 403377 233651
rect 410895 233648 410961 233651
rect 358959 233646 403377 233648
rect 358959 233590 358964 233646
rect 359020 233590 403316 233646
rect 403372 233590 403377 233646
rect 358959 233588 403377 233590
rect 358959 233585 359025 233588
rect 403311 233585 403377 233588
rect 403458 233646 410961 233648
rect 403458 233590 410900 233646
rect 410956 233590 410961 233646
rect 403458 233588 410961 233590
rect 144015 233500 144081 233503
rect 140802 233498 144081 233500
rect 140802 233442 144020 233498
rect 144076 233442 144081 233498
rect 140802 233440 144081 233442
rect 144015 233437 144081 233440
rect 302991 233500 303057 233503
rect 398991 233500 399057 233503
rect 302991 233498 399057 233500
rect 302991 233442 302996 233498
rect 303052 233442 398996 233498
rect 399052 233442 399057 233498
rect 302991 233440 399057 233442
rect 302991 233437 303057 233440
rect 398991 233437 399057 233440
rect 401199 233500 401265 233503
rect 403458 233500 403518 233588
rect 410895 233585 410961 233588
rect 414447 233648 414513 233651
rect 442810 233648 442816 233650
rect 414447 233646 442816 233648
rect 414447 233590 414452 233646
rect 414508 233590 442816 233646
rect 414447 233588 442816 233590
rect 414447 233585 414513 233588
rect 442810 233586 442816 233588
rect 442880 233586 442886 233650
rect 443631 233648 443697 233651
rect 444111 233648 444177 233651
rect 443631 233646 444177 233648
rect 443631 233590 443636 233646
rect 443692 233590 444116 233646
rect 444172 233590 444177 233646
rect 443631 233588 444177 233590
rect 443631 233585 443697 233588
rect 444111 233585 444177 233588
rect 401199 233498 403518 233500
rect 401199 233442 401204 233498
rect 401260 233442 403518 233498
rect 401199 233440 403518 233442
rect 408687 233500 408753 233503
rect 408975 233500 409041 233503
rect 408687 233498 409041 233500
rect 408687 233442 408692 233498
rect 408748 233442 408980 233498
rect 409036 233442 409041 233498
rect 408687 233440 409041 233442
rect 401199 233437 401265 233440
rect 408687 233437 408753 233440
rect 408975 233437 409041 233440
rect 413487 233500 413553 233503
rect 418287 233500 418353 233503
rect 413487 233498 418353 233500
rect 413487 233442 413492 233498
rect 413548 233442 418292 233498
rect 418348 233442 418353 233498
rect 413487 233440 418353 233442
rect 413487 233437 413553 233440
rect 418287 233437 418353 233440
rect 423375 233500 423441 233503
rect 443002 233500 443008 233502
rect 423375 233498 443008 233500
rect 423375 233442 423380 233498
rect 423436 233442 443008 233498
rect 423375 233440 443008 233442
rect 423375 233437 423441 233440
rect 443002 233438 443008 233440
rect 443072 233438 443078 233502
rect 443919 233500 443985 233503
rect 460815 233500 460881 233503
rect 443919 233498 460881 233500
rect 443919 233442 443924 233498
rect 443980 233442 460820 233498
rect 460876 233442 460881 233498
rect 443919 233440 460881 233442
rect 443919 233437 443985 233440
rect 460815 233437 460881 233440
rect 41338 233290 41344 233354
rect 41408 233352 41414 233354
rect 41775 233352 41841 233355
rect 41408 233350 41841 233352
rect 41408 233294 41780 233350
rect 41836 233294 41841 233350
rect 41408 233292 41841 233294
rect 41408 233290 41414 233292
rect 41775 233289 41841 233292
rect 384399 233352 384465 233355
rect 499119 233352 499185 233355
rect 384399 233350 499185 233352
rect 384399 233294 384404 233350
rect 384460 233294 499124 233350
rect 499180 233294 499185 233350
rect 384399 233292 499185 233294
rect 384399 233289 384465 233292
rect 499119 233289 499185 233292
rect 380271 233204 380337 233207
rect 495087 233204 495153 233207
rect 380271 233202 495153 233204
rect 380271 233146 380276 233202
rect 380332 233146 495092 233202
rect 495148 233146 495153 233202
rect 380271 233144 495153 233146
rect 380271 233141 380337 233144
rect 495087 233141 495153 233144
rect 383631 233056 383697 233059
rect 498351 233056 498417 233059
rect 383631 233054 498417 233056
rect 383631 232998 383636 233054
rect 383692 232998 498356 233054
rect 498412 232998 498417 233054
rect 383631 232996 498417 232998
rect 383631 232993 383697 232996
rect 498351 232993 498417 232996
rect 332847 232908 332913 232911
rect 447567 232908 447633 232911
rect 332847 232906 447633 232908
rect 332847 232850 332852 232906
rect 332908 232850 447572 232906
rect 447628 232850 447633 232906
rect 332847 232848 447633 232850
rect 332847 232845 332913 232848
rect 447567 232845 447633 232848
rect 331023 232760 331089 232763
rect 445743 232760 445809 232763
rect 331023 232758 445809 232760
rect 331023 232702 331028 232758
rect 331084 232702 445748 232758
rect 445804 232702 445809 232758
rect 331023 232700 445809 232702
rect 331023 232697 331089 232700
rect 445743 232697 445809 232700
rect 446074 232698 446080 232762
rect 446144 232760 446150 232762
rect 450874 232760 450880 232762
rect 446144 232700 450880 232760
rect 446144 232698 446150 232700
rect 450874 232698 450880 232700
rect 450944 232698 450950 232762
rect 343119 232612 343185 232615
rect 435279 232612 435345 232615
rect 343119 232610 435345 232612
rect 343119 232554 343124 232610
rect 343180 232554 435284 232610
rect 435340 232554 435345 232610
rect 343119 232552 435345 232554
rect 343119 232549 343185 232552
rect 435279 232549 435345 232552
rect 435471 232612 435537 232615
rect 503919 232612 503985 232615
rect 435471 232610 503985 232612
rect 435471 232554 435476 232610
rect 435532 232554 503924 232610
rect 503980 232554 503985 232610
rect 435471 232552 503985 232554
rect 435471 232549 435537 232552
rect 503919 232549 503985 232552
rect 145455 232464 145521 232467
rect 140832 232462 145521 232464
rect 140832 232406 145460 232462
rect 145516 232406 145521 232462
rect 140832 232404 145521 232406
rect 145455 232401 145521 232404
rect 330639 232464 330705 232467
rect 445359 232464 445425 232467
rect 330639 232462 445425 232464
rect 330639 232406 330644 232462
rect 330700 232406 445364 232462
rect 445420 232406 445425 232462
rect 330639 232404 445425 232406
rect 330639 232401 330705 232404
rect 445359 232401 445425 232404
rect 453327 232464 453393 232467
rect 453711 232464 453777 232467
rect 453327 232462 453777 232464
rect 453327 232406 453332 232462
rect 453388 232406 453716 232462
rect 453772 232406 453777 232462
rect 453327 232404 453777 232406
rect 453327 232401 453393 232404
rect 453711 232401 453777 232404
rect 331695 232316 331761 232319
rect 446511 232316 446577 232319
rect 331695 232314 446577 232316
rect 331695 232258 331700 232314
rect 331756 232258 446516 232314
rect 446572 232258 446577 232314
rect 331695 232256 446577 232258
rect 331695 232253 331761 232256
rect 446511 232253 446577 232256
rect 287098 232106 287104 232170
rect 287168 232168 287174 232170
rect 389679 232168 389745 232171
rect 412623 232168 412689 232171
rect 287168 232166 389745 232168
rect 287168 232110 389684 232166
rect 389740 232110 389745 232166
rect 287168 232108 389745 232110
rect 287168 232106 287174 232108
rect 389679 232105 389745 232108
rect 389826 232166 412689 232168
rect 389826 232110 412628 232166
rect 412684 232110 412689 232166
rect 389826 232108 412689 232110
rect 288442 231958 288448 232022
rect 288512 232020 288518 232022
rect 389826 232020 389886 232108
rect 412623 232105 412689 232108
rect 414543 232168 414609 232171
rect 429039 232168 429105 232171
rect 443386 232168 443392 232170
rect 414543 232166 428478 232168
rect 414543 232110 414548 232166
rect 414604 232110 428478 232166
rect 414543 232108 428478 232110
rect 414543 232105 414609 232108
rect 413391 232020 413457 232023
rect 288512 231960 389886 232020
rect 390018 232018 413457 232020
rect 390018 231962 413396 232018
rect 413452 231962 413457 232018
rect 390018 231960 413457 231962
rect 288512 231958 288518 231960
rect 288826 231810 288832 231874
rect 288896 231872 288902 231874
rect 390018 231872 390078 231960
rect 413391 231957 413457 231960
rect 414639 232020 414705 232023
rect 428418 232020 428478 232108
rect 429039 232166 443392 232168
rect 429039 232110 429044 232166
rect 429100 232110 443392 232166
rect 429039 232108 443392 232110
rect 429039 232105 429105 232108
rect 443386 232106 443392 232108
rect 443456 232106 443462 232170
rect 443535 232168 443601 232171
rect 453423 232168 453489 232171
rect 443535 232166 453489 232168
rect 443535 232110 443540 232166
rect 443596 232110 453428 232166
rect 453484 232110 453489 232166
rect 443535 232108 453489 232110
rect 443535 232105 443601 232108
rect 453423 232105 453489 232108
rect 453999 232168 454065 232171
rect 509871 232168 509937 232171
rect 453999 232166 509937 232168
rect 453999 232110 454004 232166
rect 454060 232110 509876 232166
rect 509932 232110 509937 232166
rect 453999 232108 509937 232110
rect 453999 232105 454065 232108
rect 509871 232105 509937 232108
rect 436815 232020 436881 232023
rect 414639 232018 428286 232020
rect 414639 231962 414644 232018
rect 414700 231962 428286 232018
rect 414639 231960 428286 231962
rect 428418 232018 436881 232020
rect 428418 231962 436820 232018
rect 436876 231962 436881 232018
rect 428418 231960 436881 231962
rect 414639 231957 414705 231960
rect 288896 231812 390078 231872
rect 397359 231872 397425 231875
rect 406575 231872 406641 231875
rect 397359 231870 406641 231872
rect 397359 231814 397364 231870
rect 397420 231814 406580 231870
rect 406636 231814 406641 231870
rect 397359 231812 406641 231814
rect 288896 231810 288902 231812
rect 397359 231809 397425 231812
rect 406575 231809 406641 231812
rect 406959 231872 407025 231875
rect 427983 231872 428049 231875
rect 406959 231870 428049 231872
rect 406959 231814 406964 231870
rect 407020 231814 427988 231870
rect 428044 231814 428049 231870
rect 406959 231812 428049 231814
rect 428226 231872 428286 231960
rect 436815 231957 436881 231960
rect 438447 232020 438513 232023
rect 506991 232020 507057 232023
rect 438447 232018 507057 232020
rect 438447 231962 438452 232018
rect 438508 231962 506996 232018
rect 507052 231962 507057 232018
rect 438447 231960 507057 231962
rect 438447 231957 438513 231960
rect 506991 231957 507057 231960
rect 435087 231872 435153 231875
rect 428226 231870 435153 231872
rect 428226 231814 435092 231870
rect 435148 231814 435153 231870
rect 428226 231812 435153 231814
rect 406959 231809 407025 231812
rect 427983 231809 428049 231812
rect 435087 231809 435153 231812
rect 435855 231872 435921 231875
rect 504303 231872 504369 231875
rect 435855 231870 504369 231872
rect 435855 231814 435860 231870
rect 435916 231814 504308 231870
rect 504364 231814 504369 231870
rect 435855 231812 504369 231814
rect 435855 231809 435921 231812
rect 504303 231809 504369 231812
rect 41775 231726 41841 231727
rect 41722 231662 41728 231726
rect 41792 231724 41841 231726
rect 383247 231724 383313 231727
rect 498159 231724 498225 231727
rect 41792 231722 41884 231724
rect 41836 231666 41884 231722
rect 41792 231664 41884 231666
rect 383247 231722 498225 231724
rect 383247 231666 383252 231722
rect 383308 231666 498164 231722
rect 498220 231666 498225 231722
rect 383247 231664 498225 231666
rect 41792 231662 41841 231664
rect 41775 231661 41841 231662
rect 383247 231661 383313 231664
rect 498159 231661 498225 231664
rect 41871 231578 41937 231579
rect 41871 231576 41920 231578
rect 41828 231574 41920 231576
rect 41828 231518 41876 231574
rect 41828 231516 41920 231518
rect 41871 231514 41920 231516
rect 41984 231514 41990 231578
rect 377391 231576 377457 231579
rect 492111 231576 492177 231579
rect 377391 231574 492177 231576
rect 377391 231518 377396 231574
rect 377452 231518 492116 231574
rect 492172 231518 492177 231574
rect 377391 231516 492177 231518
rect 41871 231513 41937 231514
rect 377391 231513 377457 231516
rect 492111 231513 492177 231516
rect 337935 231428 338001 231431
rect 440079 231428 440145 231431
rect 337935 231426 440145 231428
rect 337935 231370 337940 231426
rect 337996 231370 440084 231426
rect 440140 231370 440145 231426
rect 337935 231368 440145 231370
rect 337935 231365 338001 231368
rect 440079 231365 440145 231368
rect 440559 231428 440625 231431
rect 506511 231428 506577 231431
rect 440559 231426 506577 231428
rect 440559 231370 440564 231426
rect 440620 231370 506516 231426
rect 506572 231370 506577 231426
rect 440559 231368 506577 231370
rect 440559 231365 440625 231368
rect 506511 231365 506577 231368
rect 144015 231280 144081 231283
rect 140832 231278 144081 231280
rect 140832 231222 144020 231278
rect 144076 231222 144081 231278
rect 140832 231220 144081 231222
rect 144015 231217 144081 231220
rect 389679 231280 389745 231283
rect 406383 231280 406449 231283
rect 389679 231278 406449 231280
rect 389679 231222 389684 231278
rect 389740 231222 406388 231278
rect 406444 231222 406449 231278
rect 389679 231220 406449 231222
rect 389679 231217 389745 231220
rect 406383 231217 406449 231220
rect 406575 231280 406641 231283
rect 489615 231280 489681 231283
rect 406575 231278 489681 231280
rect 406575 231222 406580 231278
rect 406636 231222 489620 231278
rect 489676 231222 489681 231278
rect 406575 231220 489681 231222
rect 406575 231217 406641 231220
rect 489615 231217 489681 231220
rect 356175 231132 356241 231135
rect 452079 231132 452145 231135
rect 356175 231130 452145 231132
rect 356175 231074 356180 231130
rect 356236 231074 452084 231130
rect 452140 231074 452145 231130
rect 356175 231072 452145 231074
rect 356175 231069 356241 231072
rect 452079 231069 452145 231072
rect 342831 230984 342897 230987
rect 436911 230984 436977 230987
rect 439983 230984 440049 230987
rect 342831 230982 430590 230984
rect 342831 230926 342836 230982
rect 342892 230926 430590 230982
rect 342831 230924 430590 230926
rect 342831 230921 342897 230924
rect 342063 230836 342129 230839
rect 428847 230836 428913 230839
rect 342063 230834 428913 230836
rect 342063 230778 342068 230834
rect 342124 230778 428852 230834
rect 428908 230778 428913 230834
rect 342063 230776 428913 230778
rect 430530 230836 430590 230924
rect 436911 230982 440049 230984
rect 436911 230926 436916 230982
rect 436972 230926 439988 230982
rect 440044 230926 440049 230982
rect 436911 230924 440049 230926
rect 436911 230921 436977 230924
rect 439983 230921 440049 230924
rect 441039 230984 441105 230987
rect 508335 230984 508401 230987
rect 441039 230982 508401 230984
rect 441039 230926 441044 230982
rect 441100 230926 508340 230982
rect 508396 230926 508401 230982
rect 441039 230924 508401 230926
rect 441039 230921 441105 230924
rect 508335 230921 508401 230924
rect 442618 230836 442624 230838
rect 430530 230776 442624 230836
rect 342063 230773 342129 230776
rect 428847 230773 428913 230776
rect 442618 230774 442624 230776
rect 442688 230774 442694 230838
rect 442767 230836 442833 230839
rect 450927 230836 450993 230839
rect 442767 230834 450993 230836
rect 442767 230778 442772 230834
rect 442828 230778 450932 230834
rect 450988 230778 450993 230834
rect 442767 230776 450993 230778
rect 442767 230773 442833 230776
rect 450927 230773 450993 230776
rect 398127 230688 398193 230691
rect 451695 230688 451761 230691
rect 398127 230686 451761 230688
rect 398127 230630 398132 230686
rect 398188 230630 451700 230686
rect 451756 230630 451761 230686
rect 398127 230628 451761 230630
rect 398127 230625 398193 230628
rect 451695 230625 451761 230628
rect 372207 230540 372273 230543
rect 488463 230540 488529 230543
rect 372207 230538 488529 230540
rect 372207 230482 372212 230538
rect 372268 230482 488468 230538
rect 488524 230482 488529 230538
rect 372207 230480 488529 230482
rect 372207 230477 372273 230480
rect 488463 230477 488529 230480
rect 204879 230394 204945 230395
rect 204879 230392 204928 230394
rect 204836 230390 204928 230392
rect 204836 230334 204884 230390
rect 204836 230332 204928 230334
rect 204879 230330 204928 230332
rect 204992 230330 204998 230394
rect 207418 230330 207424 230394
rect 207488 230392 207494 230394
rect 208047 230392 208113 230395
rect 208431 230394 208497 230395
rect 208378 230392 208384 230394
rect 207488 230390 208113 230392
rect 207488 230334 208052 230390
rect 208108 230334 208113 230390
rect 207488 230332 208113 230334
rect 208340 230332 208384 230392
rect 208448 230390 208497 230394
rect 208492 230334 208497 230390
rect 207488 230330 207494 230332
rect 204879 230329 204945 230330
rect 208047 230329 208113 230332
rect 208378 230330 208384 230332
rect 208448 230330 208497 230334
rect 288250 230330 288256 230394
rect 288320 230392 288326 230394
rect 360015 230392 360081 230395
rect 288320 230390 360081 230392
rect 288320 230334 360020 230390
rect 360076 230334 360081 230390
rect 288320 230332 360081 230334
rect 288320 230330 288326 230332
rect 208431 230329 208497 230330
rect 360015 230329 360081 230332
rect 402255 230392 402321 230395
rect 404367 230392 404433 230395
rect 402255 230390 404433 230392
rect 402255 230334 402260 230390
rect 402316 230334 404372 230390
rect 404428 230334 404433 230390
rect 402255 230332 404433 230334
rect 402255 230329 402321 230332
rect 404367 230329 404433 230332
rect 409071 230392 409137 230395
rect 413103 230392 413169 230395
rect 409071 230390 413169 230392
rect 409071 230334 409076 230390
rect 409132 230334 413108 230390
rect 413164 230334 413169 230390
rect 409071 230332 413169 230334
rect 409071 230329 409137 230332
rect 413103 230329 413169 230332
rect 415215 230392 415281 230395
rect 443631 230394 443697 230395
rect 441850 230392 441856 230394
rect 415215 230390 441856 230392
rect 415215 230334 415220 230390
rect 415276 230334 441856 230390
rect 415215 230332 441856 230334
rect 415215 230329 415281 230332
rect 441850 230330 441856 230332
rect 441920 230330 441926 230394
rect 443578 230330 443584 230394
rect 443648 230392 443697 230394
rect 443648 230390 443740 230392
rect 443692 230334 443740 230390
rect 443648 230332 443740 230334
rect 443648 230330 443697 230332
rect 443631 230329 443697 230330
rect 204730 230182 204736 230246
rect 204800 230244 204806 230246
rect 205455 230244 205521 230247
rect 204800 230242 205521 230244
rect 204800 230186 205460 230242
rect 205516 230186 205521 230242
rect 204800 230184 205521 230186
rect 204800 230182 204806 230184
rect 205455 230181 205521 230184
rect 383919 230244 383985 230247
rect 498735 230244 498801 230247
rect 383919 230242 498801 230244
rect 383919 230186 383924 230242
rect 383980 230186 498740 230242
rect 498796 230186 498801 230242
rect 383919 230184 498801 230186
rect 383919 230181 383985 230184
rect 498735 230181 498801 230184
rect 204495 230096 204561 230099
rect 204975 230096 205041 230099
rect 204495 230094 205041 230096
rect 204495 230038 204500 230094
rect 204556 230038 204980 230094
rect 205036 230038 205041 230094
rect 204495 230036 205041 230038
rect 204495 230033 204561 230036
rect 204975 230033 205041 230036
rect 379599 230096 379665 230099
rect 494319 230096 494385 230099
rect 379599 230094 494385 230096
rect 379599 230038 379604 230094
rect 379660 230038 494324 230094
rect 494380 230038 494385 230094
rect 379599 230036 494385 230038
rect 379599 230033 379665 230036
rect 494319 230033 494385 230036
rect 41146 229738 41152 229802
rect 41216 229800 41222 229802
rect 41775 229800 41841 229803
rect 41216 229798 41841 229800
rect 41216 229742 41780 229798
rect 41836 229742 41841 229798
rect 41216 229740 41841 229742
rect 41216 229738 41222 229740
rect 41775 229737 41841 229740
rect 140802 229504 140862 229992
rect 378159 229948 378225 229951
rect 492879 229948 492945 229951
rect 378159 229946 492945 229948
rect 378159 229890 378164 229946
rect 378220 229890 492884 229946
rect 492940 229890 492945 229946
rect 378159 229888 492945 229890
rect 378159 229885 378225 229888
rect 492879 229885 492945 229888
rect 381807 229800 381873 229803
rect 496527 229800 496593 229803
rect 381807 229798 496593 229800
rect 381807 229742 381812 229798
rect 381868 229742 496532 229798
rect 496588 229742 496593 229798
rect 381807 229740 496593 229742
rect 381807 229737 381873 229740
rect 496527 229737 496593 229740
rect 368079 229652 368145 229655
rect 373359 229652 373425 229655
rect 368079 229650 373425 229652
rect 368079 229594 368084 229650
rect 368140 229594 373364 229650
rect 373420 229594 373425 229650
rect 368079 229592 373425 229594
rect 368079 229589 368145 229592
rect 373359 229589 373425 229592
rect 385455 229652 385521 229655
rect 500271 229652 500337 229655
rect 385455 229650 500337 229652
rect 385455 229594 385460 229650
rect 385516 229594 500276 229650
rect 500332 229594 500337 229650
rect 385455 229592 500337 229594
rect 385455 229589 385521 229592
rect 500271 229589 500337 229592
rect 144111 229504 144177 229507
rect 140802 229502 144177 229504
rect 140802 229446 144116 229502
rect 144172 229446 144177 229502
rect 140802 229444 144177 229446
rect 144111 229441 144177 229444
rect 354063 229504 354129 229507
rect 358767 229504 358833 229507
rect 354063 229502 358833 229504
rect 354063 229446 354068 229502
rect 354124 229446 358772 229502
rect 358828 229446 358833 229502
rect 354063 229444 358833 229446
rect 354063 229441 354129 229444
rect 358767 229441 358833 229444
rect 384687 229504 384753 229507
rect 499503 229504 499569 229507
rect 384687 229502 499569 229504
rect 384687 229446 384692 229502
rect 384748 229446 499508 229502
rect 499564 229446 499569 229502
rect 384687 229444 499569 229446
rect 384687 229441 384753 229444
rect 499503 229441 499569 229444
rect 674415 229504 674481 229507
rect 674415 229502 674784 229504
rect 674415 229446 674420 229502
rect 674476 229446 674784 229502
rect 674415 229444 674784 229446
rect 674415 229441 674481 229444
rect 369231 229356 369297 229359
rect 487023 229356 487089 229359
rect 369231 229354 487089 229356
rect 369231 229298 369236 229354
rect 369292 229298 487028 229354
rect 487084 229298 487089 229354
rect 369231 229296 487089 229298
rect 369231 229293 369297 229296
rect 487023 229293 487089 229296
rect 286714 229146 286720 229210
rect 286784 229208 286790 229210
rect 354159 229208 354225 229211
rect 286784 229206 354225 229208
rect 286784 229150 354164 229206
rect 354220 229150 354225 229206
rect 286784 229148 354225 229150
rect 286784 229146 286790 229148
rect 354159 229145 354225 229148
rect 367791 229208 367857 229211
rect 486255 229208 486321 229211
rect 367791 229206 486321 229208
rect 367791 229150 367796 229206
rect 367852 229150 486260 229206
rect 486316 229150 486321 229206
rect 367791 229148 486321 229150
rect 367791 229145 367857 229148
rect 486255 229145 486321 229148
rect 40954 228998 40960 229062
rect 41024 229060 41030 229062
rect 41775 229060 41841 229063
rect 41024 229058 41841 229060
rect 41024 229002 41780 229058
rect 41836 229002 41841 229058
rect 41024 229000 41841 229002
rect 41024 228998 41030 229000
rect 41775 228997 41841 229000
rect 287290 228998 287296 229062
rect 287360 229060 287366 229062
rect 353007 229060 353073 229063
rect 287360 229058 353073 229060
rect 287360 229002 353012 229058
rect 353068 229002 353073 229058
rect 287360 229000 353073 229002
rect 287360 228998 287366 229000
rect 353007 228997 353073 229000
rect 370671 229060 370737 229063
rect 487695 229060 487761 229063
rect 370671 229058 487761 229060
rect 370671 229002 370676 229058
rect 370732 229002 487700 229058
rect 487756 229002 487761 229058
rect 370671 229000 487761 229002
rect 370671 228997 370737 229000
rect 487695 228997 487761 229000
rect 144015 228912 144081 228915
rect 140832 228910 144081 228912
rect 140832 228854 144020 228910
rect 144076 228854 144081 228910
rect 140832 228852 144081 228854
rect 144015 228849 144081 228852
rect 288058 228850 288064 228914
rect 288128 228912 288134 228914
rect 416367 228912 416433 228915
rect 288128 228910 416433 228912
rect 288128 228854 416372 228910
rect 416428 228854 416433 228910
rect 288128 228852 416433 228854
rect 288128 228850 288134 228852
rect 416367 228849 416433 228852
rect 416559 228912 416625 228915
rect 422319 228912 422385 228915
rect 416559 228910 422385 228912
rect 416559 228854 416564 228910
rect 416620 228854 422324 228910
rect 422380 228854 422385 228910
rect 416559 228852 422385 228854
rect 416559 228849 416625 228852
rect 422319 228849 422385 228852
rect 425871 228912 425937 228915
rect 437583 228912 437649 228915
rect 425871 228910 437649 228912
rect 425871 228854 425876 228910
rect 425932 228854 437588 228910
rect 437644 228854 437649 228910
rect 425871 228852 437649 228854
rect 425871 228849 425937 228852
rect 437583 228849 437649 228852
rect 440559 228912 440625 228915
rect 448719 228912 448785 228915
rect 440559 228910 448785 228912
rect 440559 228854 440564 228910
rect 440620 228854 448724 228910
rect 448780 228854 448785 228910
rect 440559 228852 448785 228854
rect 440559 228849 440625 228852
rect 448719 228849 448785 228852
rect 674703 228912 674769 228915
rect 674703 228910 674814 228912
rect 674703 228854 674708 228910
rect 674764 228854 674814 228910
rect 674703 228849 674814 228854
rect 202575 228764 202641 228767
rect 167106 228762 202641 228764
rect 167106 228706 202580 228762
rect 202636 228706 202641 228762
rect 167106 228704 202641 228706
rect 156879 228616 156945 228619
rect 167106 228616 167166 228704
rect 202575 228701 202641 228704
rect 378927 228764 378993 228767
rect 493647 228764 493713 228767
rect 378927 228762 493713 228764
rect 378927 228706 378932 228762
rect 378988 228706 493652 228762
rect 493708 228706 493713 228762
rect 378927 228704 493713 228706
rect 378927 228701 378993 228704
rect 493647 228701 493713 228704
rect 674754 228660 674814 228849
rect 156879 228614 167166 228616
rect 156879 228558 156884 228614
rect 156940 228558 167166 228614
rect 156879 228556 167166 228558
rect 382575 228616 382641 228619
rect 497295 228616 497361 228619
rect 382575 228614 497361 228616
rect 382575 228558 382580 228614
rect 382636 228558 497300 228614
rect 497356 228558 497361 228614
rect 382575 228556 497361 228558
rect 156879 228553 156945 228556
rect 382575 228553 382641 228556
rect 497295 228553 497361 228556
rect 358479 228468 358545 228471
rect 361071 228468 361137 228471
rect 358479 228466 361137 228468
rect 358479 228410 358484 228466
rect 358540 228410 361076 228466
rect 361132 228410 361137 228466
rect 358479 228408 361137 228410
rect 358479 228405 358545 228408
rect 361071 228405 361137 228408
rect 374319 228468 374385 228471
rect 484815 228468 484881 228471
rect 374319 228466 484881 228468
rect 374319 228410 374324 228466
rect 374380 228410 484820 228466
rect 484876 228410 484881 228466
rect 374319 228408 484881 228410
rect 374319 228405 374385 228408
rect 484815 228405 484881 228408
rect 344943 228320 345009 228323
rect 453039 228320 453105 228323
rect 344943 228318 453105 228320
rect 344943 228262 344948 228318
rect 345004 228262 453044 228318
rect 453100 228262 453105 228318
rect 344943 228260 453105 228262
rect 344943 228257 345009 228260
rect 453039 228257 453105 228260
rect 345327 228172 345393 228175
rect 393039 228172 393105 228175
rect 345327 228170 393105 228172
rect 345327 228114 345332 228170
rect 345388 228114 393044 228170
rect 393100 228114 393105 228170
rect 345327 228112 393105 228114
rect 345327 228109 345393 228112
rect 393039 228109 393105 228112
rect 395439 228172 395505 228175
rect 403311 228172 403377 228175
rect 395439 228170 403377 228172
rect 395439 228114 395444 228170
rect 395500 228114 403316 228170
rect 403372 228114 403377 228170
rect 395439 228112 403377 228114
rect 395439 228109 395505 228112
rect 403311 228109 403377 228112
rect 408879 228172 408945 228175
rect 409359 228172 409425 228175
rect 408879 228170 409425 228172
rect 408879 228114 408884 228170
rect 408940 228114 409364 228170
rect 409420 228114 409425 228170
rect 408879 228112 409425 228114
rect 408879 228109 408945 228112
rect 409359 228109 409425 228112
rect 409647 228172 409713 228175
rect 413242 228172 413248 228174
rect 409647 228170 413248 228172
rect 409647 228114 409652 228170
rect 409708 228114 413248 228170
rect 409647 228112 413248 228114
rect 409647 228109 409713 228112
rect 413242 228110 413248 228112
rect 413312 228110 413318 228174
rect 413967 228172 414033 228175
rect 483279 228172 483345 228175
rect 413967 228170 483345 228172
rect 413967 228114 413972 228170
rect 414028 228114 483284 228170
rect 483340 228114 483345 228170
rect 413967 228112 483345 228114
rect 413967 228109 414033 228112
rect 483279 228109 483345 228112
rect 393135 228024 393201 228027
rect 441274 228024 441280 228026
rect 393135 228022 441280 228024
rect 393135 227966 393140 228022
rect 393196 227966 441280 228022
rect 393135 227964 441280 227966
rect 393135 227961 393201 227964
rect 441274 227962 441280 227964
rect 441344 227962 441350 228026
rect 358383 227876 358449 227879
rect 359151 227876 359217 227879
rect 358383 227874 359217 227876
rect 358383 227818 358388 227874
rect 358444 227818 359156 227874
rect 359212 227818 359217 227874
rect 358383 227816 359217 227818
rect 358383 227813 358449 227816
rect 359151 227813 359217 227816
rect 398895 227876 398961 227879
rect 413967 227876 414033 227879
rect 398895 227874 414033 227876
rect 398895 227818 398900 227874
rect 398956 227818 413972 227874
rect 414028 227818 414033 227874
rect 398895 227816 414033 227818
rect 398895 227813 398961 227816
rect 413967 227813 414033 227816
rect 414159 227876 414225 227879
rect 443770 227876 443776 227878
rect 414159 227874 443776 227876
rect 414159 227818 414164 227874
rect 414220 227818 443776 227874
rect 414159 227816 443776 227818
rect 414159 227813 414225 227816
rect 443770 227814 443776 227816
rect 443840 227814 443846 227878
rect 674415 227876 674481 227879
rect 674415 227874 674784 227876
rect 674415 227818 674420 227874
rect 674476 227818 674784 227874
rect 674415 227816 674784 227818
rect 674415 227813 674481 227816
rect 145551 227728 145617 227731
rect 140832 227726 145617 227728
rect 140832 227670 145556 227726
rect 145612 227670 145617 227726
rect 140832 227668 145617 227670
rect 145551 227665 145617 227668
rect 202575 227728 202641 227731
rect 207610 227728 207616 227730
rect 202575 227726 207616 227728
rect 202575 227670 202580 227726
rect 202636 227670 207616 227726
rect 202575 227668 207616 227670
rect 202575 227665 202641 227668
rect 207610 227666 207616 227668
rect 207680 227728 207686 227730
rect 343791 227728 343857 227731
rect 207680 227726 343857 227728
rect 207680 227670 343796 227726
rect 343852 227670 343857 227726
rect 207680 227668 343857 227670
rect 207680 227666 207686 227668
rect 343791 227665 343857 227668
rect 381135 227728 381201 227731
rect 495855 227728 495921 227731
rect 381135 227726 495921 227728
rect 381135 227670 381140 227726
rect 381196 227670 495860 227726
rect 495916 227670 495921 227726
rect 381135 227668 495921 227670
rect 381135 227665 381201 227668
rect 495855 227665 495921 227668
rect 40570 227518 40576 227582
rect 40640 227580 40646 227582
rect 41530 227580 41536 227582
rect 40640 227520 41536 227580
rect 40640 227518 40646 227520
rect 41530 227518 41536 227520
rect 41600 227518 41606 227582
rect 345711 227580 345777 227583
rect 432591 227580 432657 227583
rect 345711 227578 432657 227580
rect 345711 227522 345716 227578
rect 345772 227522 432596 227578
rect 432652 227522 432657 227578
rect 345711 227520 432657 227522
rect 345711 227517 345777 227520
rect 432591 227517 432657 227520
rect 303759 227432 303825 227435
rect 423375 227432 423441 227435
rect 303759 227430 423441 227432
rect 303759 227374 303764 227430
rect 303820 227374 423380 227430
rect 423436 227374 423441 227430
rect 303759 227372 423441 227374
rect 303759 227369 303825 227372
rect 423375 227369 423441 227372
rect 435183 227432 435249 227435
rect 443194 227432 443200 227434
rect 435183 227430 443200 227432
rect 435183 227374 435188 227430
rect 435244 227374 443200 227430
rect 435183 227372 443200 227374
rect 435183 227369 435249 227372
rect 443194 227370 443200 227372
rect 443264 227370 443270 227434
rect 40378 227222 40384 227286
rect 40448 227284 40454 227286
rect 41775 227284 41841 227287
rect 40448 227282 41841 227284
rect 40448 227226 41780 227282
rect 41836 227226 41841 227282
rect 40448 227224 41841 227226
rect 40448 227222 40454 227224
rect 41775 227221 41841 227224
rect 305199 227284 305265 227287
rect 423471 227284 423537 227287
rect 432879 227284 432945 227287
rect 305199 227282 423537 227284
rect 305199 227226 305204 227282
rect 305260 227226 423476 227282
rect 423532 227226 423537 227282
rect 305199 227224 423537 227226
rect 305199 227221 305265 227224
rect 423471 227221 423537 227224
rect 423618 227282 432945 227284
rect 423618 227226 432884 227282
rect 432940 227226 432945 227282
rect 423618 227224 432945 227226
rect 303375 227136 303441 227139
rect 423375 227136 423441 227139
rect 303375 227134 423441 227136
rect 303375 227078 303380 227134
rect 303436 227078 423380 227134
rect 423436 227078 423441 227134
rect 303375 227076 423441 227078
rect 303375 227073 303441 227076
rect 423375 227073 423441 227076
rect 304527 226988 304593 226991
rect 419194 226988 419200 226990
rect 304527 226986 419200 226988
rect 304527 226930 304532 226986
rect 304588 226930 419200 226986
rect 304527 226928 419200 226930
rect 304527 226925 304593 226928
rect 419194 226926 419200 226928
rect 419264 226926 419270 226990
rect 419343 226988 419409 226991
rect 423618 226988 423678 227224
rect 432879 227221 432945 227224
rect 433071 227284 433137 227287
rect 452218 227284 452224 227286
rect 433071 227282 452224 227284
rect 433071 227226 433076 227282
rect 433132 227226 452224 227282
rect 433071 227224 452224 227226
rect 433071 227221 433137 227224
rect 452218 227222 452224 227224
rect 452288 227222 452294 227286
rect 675898 227222 675904 227286
rect 675968 227222 675974 227286
rect 426063 227136 426129 227139
rect 432303 227136 432369 227139
rect 426063 227134 432369 227136
rect 426063 227078 426068 227134
rect 426124 227078 432308 227134
rect 432364 227078 432369 227134
rect 426063 227076 432369 227078
rect 426063 227073 426129 227076
rect 432303 227073 432369 227076
rect 432495 227136 432561 227139
rect 453178 227136 453184 227138
rect 432495 227134 453184 227136
rect 432495 227078 432500 227134
rect 432556 227078 453184 227134
rect 432495 227076 453184 227078
rect 432495 227073 432561 227076
rect 453178 227074 453184 227076
rect 453248 227074 453254 227138
rect 675906 227032 675966 227222
rect 419343 226986 423678 226988
rect 419343 226930 419348 226986
rect 419404 226930 423678 226986
rect 419343 226928 423678 226930
rect 427599 226988 427665 226991
rect 453946 226988 453952 226990
rect 427599 226986 453952 226988
rect 427599 226930 427604 226986
rect 427660 226930 453952 226986
rect 427599 226928 453952 226930
rect 419343 226925 419409 226928
rect 427599 226925 427665 226928
rect 453946 226926 453952 226928
rect 454016 226926 454022 226990
rect 40762 226778 40768 226842
rect 40832 226840 40838 226842
rect 41775 226840 41841 226843
rect 40832 226838 41841 226840
rect 40832 226782 41780 226838
rect 41836 226782 41841 226838
rect 40832 226780 41841 226782
rect 40832 226778 40838 226780
rect 41775 226777 41841 226780
rect 207855 226840 207921 226843
rect 207994 226840 208000 226842
rect 207855 226838 208000 226840
rect 207855 226782 207860 226838
rect 207916 226782 208000 226838
rect 207855 226780 208000 226782
rect 207855 226777 207921 226780
rect 207994 226778 208000 226780
rect 208064 226778 208070 226842
rect 307407 226840 307473 226843
rect 427503 226840 427569 226843
rect 307407 226838 427569 226840
rect 307407 226782 307412 226838
rect 307468 226782 427508 226838
rect 427564 226782 427569 226838
rect 307407 226780 427569 226782
rect 307407 226777 307473 226780
rect 427503 226777 427569 226780
rect 427791 226840 427857 226843
rect 452986 226840 452992 226842
rect 427791 226838 452992 226840
rect 427791 226782 427796 226838
rect 427852 226782 452992 226838
rect 427791 226780 452992 226782
rect 427791 226777 427857 226780
rect 452986 226778 452992 226780
rect 453056 226778 453062 226842
rect 207759 226694 207825 226695
rect 207759 226690 207808 226694
rect 207872 226692 207878 226694
rect 306735 226692 306801 226695
rect 419002 226692 419008 226694
rect 207759 226634 207764 226690
rect 207759 226630 207808 226634
rect 207872 226632 207916 226692
rect 306735 226690 419008 226692
rect 306735 226634 306740 226690
rect 306796 226634 419008 226690
rect 306735 226632 419008 226634
rect 207872 226630 207878 226632
rect 207759 226629 207825 226630
rect 306735 226629 306801 226632
rect 419002 226630 419008 226632
rect 419072 226630 419078 226694
rect 419194 226630 419200 226694
rect 419264 226692 419270 226694
rect 423567 226692 423633 226695
rect 419264 226690 423633 226692
rect 419264 226634 423572 226690
rect 423628 226634 423633 226690
rect 419264 226632 423633 226634
rect 419264 226630 419270 226632
rect 423567 226629 423633 226632
rect 426159 226692 426225 226695
rect 432111 226692 432177 226695
rect 426159 226690 432177 226692
rect 426159 226634 426164 226690
rect 426220 226634 432116 226690
rect 432172 226634 432177 226690
rect 426159 226632 432177 226634
rect 426159 226629 426225 226632
rect 432111 226629 432177 226632
rect 432303 226692 432369 226695
rect 448378 226692 448384 226694
rect 432303 226690 448384 226692
rect 432303 226634 432308 226690
rect 432364 226634 448384 226690
rect 432303 226632 448384 226634
rect 432303 226629 432369 226632
rect 448378 226630 448384 226632
rect 448448 226630 448454 226694
rect 208143 226546 208209 226547
rect 208143 226542 208192 226546
rect 208256 226544 208262 226546
rect 348399 226544 348465 226547
rect 426255 226544 426321 226547
rect 208143 226486 208148 226542
rect 208143 226482 208192 226486
rect 208256 226484 208300 226544
rect 348399 226542 426321 226544
rect 348399 226486 348404 226542
rect 348460 226486 426260 226542
rect 426316 226486 426321 226542
rect 348399 226484 426321 226486
rect 208256 226482 208262 226484
rect 208143 226481 208209 226482
rect 348399 226481 348465 226484
rect 426255 226481 426321 226484
rect 428079 226544 428145 226547
rect 452410 226544 452416 226546
rect 428079 226542 452416 226544
rect 428079 226486 428084 226542
rect 428140 226486 452416 226542
rect 428079 226484 452416 226486
rect 428079 226481 428145 226484
rect 452410 226482 452416 226484
rect 452480 226482 452486 226546
rect 40570 225890 40576 225954
rect 40640 225952 40646 225954
rect 41775 225952 41841 225955
rect 40640 225950 41841 225952
rect 40640 225894 41780 225950
rect 41836 225894 41841 225950
rect 40640 225892 41841 225894
rect 140802 225952 140862 226440
rect 326895 226396 326961 226399
rect 430767 226396 430833 226399
rect 431919 226396 431985 226399
rect 326895 226394 430833 226396
rect 326895 226338 326900 226394
rect 326956 226338 430772 226394
rect 430828 226338 430833 226394
rect 326895 226336 430833 226338
rect 326895 226333 326961 226336
rect 430767 226333 430833 226336
rect 430914 226394 431985 226396
rect 430914 226338 431924 226394
rect 431980 226338 431985 226394
rect 430914 226336 431985 226338
rect 308175 226248 308241 226251
rect 430914 226248 430974 226336
rect 431919 226333 431985 226336
rect 432111 226396 432177 226399
rect 446842 226396 446848 226398
rect 432111 226394 446848 226396
rect 432111 226338 432116 226394
rect 432172 226338 446848 226394
rect 432111 226336 446848 226338
rect 432111 226333 432177 226336
rect 446842 226334 446848 226336
rect 446912 226334 446918 226398
rect 446991 226396 447057 226399
rect 452794 226396 452800 226398
rect 446991 226394 452800 226396
rect 446991 226338 446996 226394
rect 447052 226338 452800 226394
rect 446991 226336 452800 226338
rect 446991 226333 447057 226336
rect 452794 226334 452800 226336
rect 452864 226334 452870 226398
rect 308175 226246 430974 226248
rect 308175 226190 308180 226246
rect 308236 226190 430974 226246
rect 308175 226188 430974 226190
rect 431151 226248 431217 226251
rect 438255 226248 438321 226251
rect 453370 226248 453376 226250
rect 431151 226246 438321 226248
rect 431151 226190 431156 226246
rect 431212 226190 438260 226246
rect 438316 226190 438321 226246
rect 431151 226188 438321 226190
rect 308175 226185 308241 226188
rect 431151 226185 431217 226188
rect 438255 226185 438321 226188
rect 438402 226188 453376 226248
rect 305967 226100 306033 226103
rect 419247 226100 419313 226103
rect 420591 226100 420657 226103
rect 305967 226098 419313 226100
rect 305967 226042 305972 226098
rect 306028 226042 419252 226098
rect 419308 226042 419313 226098
rect 305967 226040 419313 226042
rect 305967 226037 306033 226040
rect 419247 226037 419313 226040
rect 419394 226098 420657 226100
rect 419394 226042 420596 226098
rect 420652 226042 420657 226098
rect 419394 226040 420657 226042
rect 145647 225952 145713 225955
rect 140802 225950 145713 225952
rect 140802 225894 145652 225950
rect 145708 225894 145713 225950
rect 140802 225892 145713 225894
rect 40640 225890 40646 225892
rect 41775 225889 41841 225892
rect 145647 225889 145713 225892
rect 348783 225952 348849 225955
rect 419394 225952 419454 226040
rect 420591 226037 420657 226040
rect 420783 226100 420849 226103
rect 423663 226100 423729 226103
rect 420783 226098 423729 226100
rect 420783 226042 420788 226098
rect 420844 226042 423668 226098
rect 423724 226042 423729 226098
rect 420783 226040 423729 226042
rect 420783 226037 420849 226040
rect 423663 226037 423729 226040
rect 428271 226100 428337 226103
rect 438402 226100 438462 226188
rect 453370 226186 453376 226188
rect 453440 226186 453446 226250
rect 674170 226186 674176 226250
rect 674240 226248 674246 226250
rect 674240 226188 674784 226248
rect 674240 226186 674246 226188
rect 428271 226098 438462 226100
rect 428271 226042 428276 226098
rect 428332 226042 438462 226098
rect 428271 226040 438462 226042
rect 438543 226100 438609 226103
rect 453562 226100 453568 226102
rect 438543 226098 453568 226100
rect 438543 226042 438548 226098
rect 438604 226042 453568 226098
rect 438543 226040 453568 226042
rect 428271 226037 428337 226040
rect 438543 226037 438609 226040
rect 453562 226038 453568 226040
rect 453632 226038 453638 226102
rect 348783 225950 419454 225952
rect 348783 225894 348788 225950
rect 348844 225894 419454 225950
rect 348783 225892 419454 225894
rect 419535 225952 419601 225955
rect 431823 225952 431889 225955
rect 446991 225952 447057 225955
rect 419535 225950 431889 225952
rect 419535 225894 419540 225950
rect 419596 225894 431828 225950
rect 431884 225894 431889 225950
rect 419535 225892 431889 225894
rect 348783 225889 348849 225892
rect 419535 225889 419601 225892
rect 431823 225889 431889 225892
rect 432066 225950 447057 225952
rect 432066 225894 446996 225950
rect 447052 225894 447057 225950
rect 432066 225892 447057 225894
rect 351759 225804 351825 225807
rect 418959 225804 419025 225807
rect 351759 225802 419025 225804
rect 351759 225746 351764 225802
rect 351820 225746 418964 225802
rect 419020 225746 419025 225802
rect 351759 225744 419025 225746
rect 351759 225741 351825 225744
rect 418959 225741 419025 225744
rect 419194 225742 419200 225806
rect 419264 225804 419270 225806
rect 423183 225804 423249 225807
rect 429231 225804 429297 225807
rect 419264 225744 423102 225804
rect 419264 225742 419270 225744
rect 359439 225656 359505 225659
rect 420495 225656 420561 225659
rect 359439 225654 420561 225656
rect 359439 225598 359444 225654
rect 359500 225598 420500 225654
rect 420556 225598 420561 225654
rect 359439 225596 420561 225598
rect 359439 225593 359505 225596
rect 420495 225593 420561 225596
rect 420687 225656 420753 225659
rect 420975 225656 421041 225659
rect 420687 225654 421041 225656
rect 420687 225598 420692 225654
rect 420748 225598 420980 225654
rect 421036 225598 421041 225654
rect 420687 225596 421041 225598
rect 423042 225656 423102 225744
rect 423183 225802 429297 225804
rect 423183 225746 423188 225802
rect 423244 225746 429236 225802
rect 429292 225746 429297 225802
rect 423183 225744 429297 225746
rect 423183 225741 423249 225744
rect 429231 225741 429297 225744
rect 429423 225804 429489 225807
rect 432066 225804 432126 225892
rect 446991 225889 447057 225892
rect 429423 225802 432126 225804
rect 429423 225746 429428 225802
rect 429484 225746 432126 225802
rect 429423 225744 432126 225746
rect 432879 225804 432945 225807
rect 454138 225804 454144 225806
rect 432879 225802 454144 225804
rect 432879 225746 432884 225802
rect 432940 225746 454144 225802
rect 432879 225744 454144 225746
rect 429423 225741 429489 225744
rect 432879 225741 432945 225744
rect 454138 225742 454144 225744
rect 454208 225742 454214 225806
rect 676666 225742 676672 225806
rect 676736 225742 676742 225806
rect 426159 225656 426225 225659
rect 423042 225654 426225 225656
rect 423042 225598 426164 225654
rect 426220 225598 426225 225654
rect 423042 225596 426225 225598
rect 420687 225593 420753 225596
rect 420975 225593 421041 225596
rect 426159 225593 426225 225596
rect 427311 225656 427377 225659
rect 431727 225656 431793 225659
rect 427311 225654 431793 225656
rect 427311 225598 427316 225654
rect 427372 225598 431732 225654
rect 431788 225598 431793 225654
rect 427311 225596 431793 225598
rect 427311 225593 427377 225596
rect 431727 225593 431793 225596
rect 432015 225656 432081 225659
rect 432879 225656 432945 225659
rect 432015 225654 432945 225656
rect 432015 225598 432020 225654
rect 432076 225598 432884 225654
rect 432940 225598 432945 225654
rect 432015 225596 432945 225598
rect 432015 225593 432081 225596
rect 432879 225593 432945 225596
rect 433071 225656 433137 225659
rect 447418 225656 447424 225658
rect 433071 225654 447424 225656
rect 433071 225598 433076 225654
rect 433132 225598 447424 225654
rect 433071 225596 447424 225598
rect 433071 225593 433137 225596
rect 447418 225594 447424 225596
rect 447488 225594 447494 225658
rect 676674 225582 676734 225742
rect 676674 225552 679776 225582
rect 676704 225522 679806 225552
rect 358863 225508 358929 225511
rect 421935 225508 422001 225511
rect 358863 225506 422001 225508
rect 358863 225450 358868 225506
rect 358924 225450 421940 225506
rect 421996 225450 422001 225506
rect 358863 225448 422001 225450
rect 358863 225445 358929 225448
rect 421935 225445 422001 225448
rect 423951 225508 424017 225511
rect 451066 225508 451072 225510
rect 423951 225506 451072 225508
rect 423951 225450 423956 225506
rect 424012 225450 451072 225506
rect 423951 225448 451072 225450
rect 423951 225445 424017 225448
rect 451066 225446 451072 225448
rect 451136 225446 451142 225510
rect 393231 225360 393297 225363
rect 426255 225360 426321 225363
rect 393231 225358 426321 225360
rect 393231 225302 393236 225358
rect 393292 225302 426260 225358
rect 426316 225302 426321 225358
rect 393231 225300 426321 225302
rect 393231 225297 393297 225300
rect 426255 225297 426321 225300
rect 428175 225360 428241 225363
rect 452602 225360 452608 225362
rect 428175 225358 452608 225360
rect 428175 225302 428180 225358
rect 428236 225302 452608 225358
rect 428175 225300 452608 225302
rect 428175 225297 428241 225300
rect 452602 225298 452608 225300
rect 452672 225298 452678 225362
rect 140802 225064 140862 225256
rect 391023 225212 391089 225215
rect 449722 225212 449728 225214
rect 391023 225210 449728 225212
rect 391023 225154 391028 225210
rect 391084 225154 449728 225210
rect 391023 225152 449728 225154
rect 391023 225149 391089 225152
rect 449722 225150 449728 225152
rect 449792 225150 449798 225214
rect 679746 225067 679806 225522
rect 144015 225064 144081 225067
rect 140802 225062 144081 225064
rect 140802 225006 144020 225062
rect 144076 225006 144081 225062
rect 140802 225004 144081 225006
rect 144015 225001 144081 225004
rect 386223 225064 386289 225067
rect 400239 225064 400305 225067
rect 386223 225062 400305 225064
rect 386223 225006 386228 225062
rect 386284 225006 400244 225062
rect 400300 225006 400305 225062
rect 386223 225004 400305 225006
rect 386223 225001 386289 225004
rect 400239 225001 400305 225004
rect 403023 225064 403089 225067
rect 453754 225064 453760 225066
rect 403023 225062 453760 225064
rect 403023 225006 403028 225062
rect 403084 225006 453760 225062
rect 403023 225004 453760 225006
rect 403023 225001 403089 225004
rect 453754 225002 453760 225004
rect 453824 225002 453830 225066
rect 679746 225062 679857 225067
rect 679746 225006 679796 225062
rect 679852 225006 679857 225062
rect 679746 225004 679857 225006
rect 679791 225001 679857 225004
rect 385839 224916 385905 224919
rect 430767 224916 430833 224919
rect 433263 224916 433329 224919
rect 385839 224914 430590 224916
rect 385839 224858 385844 224914
rect 385900 224858 430590 224914
rect 385839 224856 430590 224858
rect 385839 224853 385905 224856
rect 388719 224770 388785 224771
rect 388666 224768 388672 224770
rect 388628 224708 388672 224768
rect 388736 224766 388785 224770
rect 388780 224710 388785 224766
rect 388666 224706 388672 224708
rect 388736 224706 388785 224710
rect 388719 224705 388785 224706
rect 391695 224770 391761 224771
rect 391695 224766 391744 224770
rect 391808 224768 391814 224770
rect 394959 224768 395025 224771
rect 426351 224768 426417 224771
rect 391695 224710 391700 224766
rect 391695 224706 391744 224710
rect 391808 224708 391852 224768
rect 394959 224766 426417 224768
rect 394959 224710 394964 224766
rect 395020 224710 426356 224766
rect 426412 224710 426417 224766
rect 394959 224708 426417 224710
rect 391808 224706 391814 224708
rect 391695 224705 391761 224706
rect 394959 224705 395025 224708
rect 426351 224705 426417 224708
rect 426543 224768 426609 224771
rect 430383 224768 430449 224771
rect 426543 224766 430449 224768
rect 426543 224710 426548 224766
rect 426604 224710 430388 224766
rect 430444 224710 430449 224766
rect 426543 224708 430449 224710
rect 430530 224768 430590 224856
rect 430767 224914 433329 224916
rect 430767 224858 430772 224914
rect 430828 224858 433268 224914
rect 433324 224858 433329 224914
rect 430767 224856 433329 224858
rect 430767 224853 430833 224856
rect 433263 224853 433329 224856
rect 433455 224916 433521 224919
rect 447226 224916 447232 224918
rect 433455 224914 447232 224916
rect 433455 224858 433460 224914
rect 433516 224858 447232 224914
rect 433455 224856 447232 224858
rect 433455 224853 433521 224856
rect 447226 224854 447232 224856
rect 447296 224854 447302 224918
rect 431535 224768 431601 224771
rect 430530 224766 431601 224768
rect 430530 224710 431540 224766
rect 431596 224710 431601 224766
rect 430530 224708 431601 224710
rect 426543 224705 426609 224708
rect 430383 224705 430449 224708
rect 431535 224705 431601 224708
rect 431727 224768 431793 224771
rect 448570 224768 448576 224770
rect 431727 224766 448576 224768
rect 431727 224710 431732 224766
rect 431788 224710 448576 224766
rect 431727 224708 448576 224710
rect 431727 224705 431793 224708
rect 448570 224706 448576 224708
rect 448640 224706 448646 224770
rect 673978 224706 673984 224770
rect 674048 224768 674054 224770
rect 674048 224708 674784 224768
rect 674048 224706 674054 224708
rect 348015 224620 348081 224623
rect 521295 224620 521361 224623
rect 348015 224618 521361 224620
rect 348015 224562 348020 224618
rect 348076 224562 521300 224618
rect 521356 224562 521361 224618
rect 348015 224560 521361 224562
rect 348015 224557 348081 224560
rect 521295 224557 521361 224560
rect 394383 224472 394449 224475
rect 509775 224472 509841 224475
rect 394383 224470 509841 224472
rect 394383 224414 394388 224470
rect 394444 224414 509780 224470
rect 509836 224414 509841 224470
rect 394383 224412 509841 224414
rect 394383 224409 394449 224412
rect 509775 224409 509841 224412
rect 343503 224324 343569 224327
rect 429178 224324 429184 224326
rect 343503 224322 429184 224324
rect 343503 224266 343508 224322
rect 343564 224266 429184 224322
rect 343503 224264 429184 224266
rect 343503 224261 343569 224264
rect 429178 224262 429184 224264
rect 429248 224262 429254 224326
rect 429370 224262 429376 224326
rect 429440 224324 429446 224326
rect 442863 224324 442929 224327
rect 429440 224322 442929 224324
rect 429440 224266 442868 224322
rect 442924 224266 442929 224322
rect 429440 224264 442929 224266
rect 429440 224262 429446 224264
rect 442863 224261 442929 224264
rect 367119 224176 367185 224179
rect 391887 224176 391953 224179
rect 367119 224174 391953 224176
rect 367119 224118 367124 224174
rect 367180 224118 391892 224174
rect 391948 224118 391953 224174
rect 367119 224116 391953 224118
rect 367119 224113 367185 224116
rect 391887 224113 391953 224116
rect 392751 224176 392817 224179
rect 480975 224176 481041 224179
rect 501039 224176 501105 224179
rect 392751 224174 481041 224176
rect 392751 224118 392756 224174
rect 392812 224118 480980 224174
rect 481036 224118 481041 224174
rect 392751 224116 481041 224118
rect 392751 224113 392817 224116
rect 480975 224113 481041 224116
rect 495234 224174 501105 224176
rect 495234 224118 501044 224174
rect 501100 224118 501105 224174
rect 495234 224116 501105 224118
rect 144015 224028 144081 224031
rect 140832 224026 144081 224028
rect 140832 223970 144020 224026
rect 144076 223970 144081 224026
rect 140832 223968 144081 223970
rect 144015 223965 144081 223968
rect 205455 224028 205521 224031
rect 207034 224028 207040 224030
rect 205455 224026 207040 224028
rect 205455 223970 205460 224026
rect 205516 223970 207040 224026
rect 205455 223968 207040 223970
rect 205455 223965 205521 223968
rect 207034 223966 207040 223968
rect 207104 223966 207110 224030
rect 360495 224028 360561 224031
rect 395919 224028 395985 224031
rect 360495 224026 395985 224028
rect 360495 223970 360500 224026
rect 360556 223970 395924 224026
rect 395980 223970 395985 224026
rect 360495 223968 395985 223970
rect 360495 223965 360561 223968
rect 395919 223965 395985 223968
rect 398895 224028 398961 224031
rect 398895 224026 399870 224028
rect 398895 223970 398900 224026
rect 398956 223970 399870 224026
rect 398895 223968 399870 223970
rect 398895 223965 398961 223968
rect 205839 223880 205905 223883
rect 206650 223880 206656 223882
rect 205839 223878 206656 223880
rect 205839 223822 205844 223878
rect 205900 223822 206656 223878
rect 205839 223820 206656 223822
rect 205839 223817 205905 223820
rect 206650 223818 206656 223820
rect 206720 223818 206726 223882
rect 207418 223818 207424 223882
rect 207488 223880 207494 223882
rect 208047 223880 208113 223883
rect 208431 223880 208497 223883
rect 207488 223878 208113 223880
rect 207488 223822 208052 223878
rect 208108 223822 208113 223878
rect 207488 223820 208113 223822
rect 207488 223818 207494 223820
rect 208047 223817 208113 223820
rect 208194 223878 208497 223880
rect 208194 223822 208436 223878
rect 208492 223822 208497 223878
rect 208194 223820 208497 223822
rect 206266 223670 206272 223734
rect 206336 223732 206342 223734
rect 208194 223732 208254 223820
rect 208431 223817 208497 223820
rect 349167 223880 349233 223883
rect 349306 223880 349312 223882
rect 349167 223878 349312 223880
rect 349167 223822 349172 223878
rect 349228 223822 349312 223878
rect 349167 223820 349312 223822
rect 349167 223817 349233 223820
rect 349306 223818 349312 223820
rect 349376 223818 349382 223882
rect 359535 223880 359601 223883
rect 362703 223882 362769 223883
rect 359674 223880 359680 223882
rect 359535 223878 359680 223880
rect 359535 223822 359540 223878
rect 359596 223822 359680 223878
rect 359535 223820 359680 223822
rect 359535 223817 359601 223820
rect 359674 223818 359680 223820
rect 359744 223818 359750 223882
rect 362703 223880 362752 223882
rect 362660 223878 362752 223880
rect 362660 223822 362708 223878
rect 362660 223820 362752 223822
rect 362703 223818 362752 223820
rect 362816 223818 362822 223882
rect 364239 223880 364305 223883
rect 379407 223880 379473 223883
rect 388719 223882 388785 223883
rect 388666 223880 388672 223882
rect 364239 223878 379473 223880
rect 364239 223822 364244 223878
rect 364300 223822 379412 223878
rect 379468 223822 379473 223878
rect 364239 223820 379473 223822
rect 388628 223820 388672 223880
rect 388736 223878 388785 223882
rect 388780 223822 388785 223878
rect 362703 223817 362769 223818
rect 364239 223817 364305 223820
rect 379407 223817 379473 223820
rect 388666 223818 388672 223820
rect 388736 223818 388785 223822
rect 388719 223817 388785 223818
rect 390351 223880 390417 223883
rect 391695 223882 391761 223883
rect 390351 223878 390462 223880
rect 390351 223822 390356 223878
rect 390412 223822 390462 223878
rect 390351 223817 390462 223822
rect 391695 223878 391744 223882
rect 391808 223880 391814 223882
rect 391695 223822 391700 223878
rect 391695 223818 391744 223822
rect 391808 223820 391852 223880
rect 399663 223878 399729 223883
rect 399663 223822 399668 223878
rect 399724 223822 399729 223878
rect 391808 223818 391814 223820
rect 391695 223817 391761 223818
rect 399663 223817 399729 223822
rect 206336 223672 208254 223732
rect 206336 223670 206342 223672
rect 302458 223584 302464 223586
rect 293826 223524 302464 223584
rect 293826 223288 293886 223524
rect 302458 223522 302464 223524
rect 302528 223522 302534 223586
rect 380026 223584 380032 223586
rect 360018 223524 380032 223584
rect 360018 223288 360078 223524
rect 380026 223522 380032 223524
rect 380096 223522 380102 223586
rect 390402 223436 390462 223817
rect 399666 223584 399726 223817
rect 399810 223732 399870 223968
rect 400186 223966 400192 224030
rect 400256 224028 400262 224030
rect 400256 223968 430590 224028
rect 400256 223966 400262 223968
rect 400239 223880 400305 223883
rect 429615 223882 429681 223883
rect 405562 223880 405568 223882
rect 400239 223878 405568 223880
rect 400239 223822 400244 223878
rect 400300 223822 405568 223878
rect 400239 223820 405568 223822
rect 400239 223817 400305 223820
rect 405562 223818 405568 223820
rect 405632 223818 405638 223882
rect 405946 223818 405952 223882
rect 406016 223880 406022 223882
rect 429562 223880 429568 223882
rect 406016 223820 429438 223880
rect 429524 223820 429568 223880
rect 429632 223878 429681 223882
rect 429676 223822 429681 223878
rect 406016 223818 406022 223820
rect 413050 223732 413056 223734
rect 399810 223672 413056 223732
rect 413050 223670 413056 223672
rect 413120 223670 413126 223734
rect 413242 223670 413248 223734
rect 413312 223732 413318 223734
rect 428986 223732 428992 223734
rect 413312 223672 428992 223732
rect 413312 223670 413318 223672
rect 428986 223670 428992 223672
rect 429056 223670 429062 223734
rect 429378 223732 429438 223820
rect 429562 223818 429568 223820
rect 429632 223818 429681 223822
rect 430530 223880 430590 223968
rect 439546 223966 439552 224030
rect 439616 224028 439622 224030
rect 439887 224028 439953 224031
rect 439616 224026 439953 224028
rect 439616 223970 439892 224026
rect 439948 223970 439953 224026
rect 439616 223968 439953 223970
rect 439616 223966 439622 223968
rect 439887 223965 439953 223968
rect 440122 223966 440128 224030
rect 440192 224028 440198 224030
rect 440655 224028 440721 224031
rect 440943 224030 441009 224031
rect 440890 224028 440896 224030
rect 440192 224026 440721 224028
rect 440192 223970 440660 224026
rect 440716 223970 440721 224026
rect 440192 223968 440721 223970
rect 440852 223968 440896 224028
rect 440960 224026 441009 224030
rect 441004 223970 441009 224026
rect 440192 223966 440198 223968
rect 440655 223965 440721 223968
rect 440890 223966 440896 223968
rect 440960 223966 441009 223970
rect 440943 223965 441009 223966
rect 449530 223880 449536 223882
rect 430530 223820 449536 223880
rect 449530 223818 449536 223820
rect 449600 223818 449606 223882
rect 429615 223817 429681 223818
rect 429378 223672 429822 223732
rect 429562 223584 429568 223586
rect 399666 223524 429568 223584
rect 429562 223522 429568 223524
rect 429632 223522 429638 223586
rect 429762 223584 429822 223672
rect 450490 223584 450496 223586
rect 429762 223524 450496 223584
rect 450490 223522 450496 223524
rect 450560 223522 450566 223586
rect 400186 223436 400192 223438
rect 390402 223376 400192 223436
rect 400186 223374 400192 223376
rect 400256 223374 400262 223438
rect 427642 223436 427648 223438
rect 403266 223376 427648 223436
rect 253506 223228 293886 223288
rect 319746 223228 360078 223288
rect 253506 223140 253566 223228
rect 249474 223080 253566 223140
rect 206842 222930 206848 222994
rect 206912 222992 206918 222994
rect 249474 222992 249534 223080
rect 302458 223078 302464 223142
rect 302528 223140 302534 223142
rect 319746 223140 319806 223228
rect 302528 223080 319806 223140
rect 302528 223078 302534 223080
rect 380026 223078 380032 223142
rect 380096 223140 380102 223142
rect 380266 223140 380272 223142
rect 380096 223080 380272 223140
rect 380096 223078 380102 223080
rect 380266 223078 380272 223080
rect 380336 223078 380342 223142
rect 400186 223078 400192 223142
rect 400256 223140 400262 223142
rect 403266 223140 403326 223376
rect 427642 223374 427648 223376
rect 427712 223374 427718 223438
rect 429370 223374 429376 223438
rect 429440 223436 429446 223438
rect 446458 223436 446464 223438
rect 429440 223376 446464 223436
rect 429440 223374 429446 223376
rect 446458 223374 446464 223376
rect 446528 223374 446534 223438
rect 413050 223226 413056 223290
rect 413120 223288 413126 223290
rect 417466 223288 417472 223290
rect 413120 223228 417472 223288
rect 413120 223226 413126 223228
rect 417466 223226 417472 223228
rect 417536 223226 417542 223290
rect 417658 223226 417664 223290
rect 417728 223288 417734 223290
rect 446074 223288 446080 223290
rect 417728 223228 446080 223288
rect 417728 223226 417734 223228
rect 446074 223226 446080 223228
rect 446144 223226 446150 223290
rect 460866 223228 480894 223288
rect 400256 223080 403326 223140
rect 400256 223078 400262 223080
rect 206912 222932 249534 222992
rect 206912 222930 206918 222932
rect 359674 222930 359680 222994
rect 359744 222992 359750 222994
rect 439546 222992 439552 222994
rect 359744 222932 439552 222992
rect 359744 222930 359750 222932
rect 439546 222930 439552 222932
rect 439616 222930 439622 222994
rect 447802 222930 447808 222994
rect 447872 222992 447878 222994
rect 460866 222992 460926 223228
rect 480834 223140 480894 223228
rect 495234 223140 495294 224116
rect 501039 224113 501105 224116
rect 631983 224176 632049 224179
rect 633466 224176 633472 224178
rect 631983 224174 633472 224176
rect 631983 224118 631988 224174
rect 632044 224118 633472 224174
rect 631983 224116 633472 224118
rect 631983 224113 632049 224116
rect 633466 224114 633472 224116
rect 633536 224114 633542 224178
rect 631311 224028 631377 224031
rect 632506 224028 632512 224030
rect 631311 224026 632512 224028
rect 631311 223970 631316 224026
rect 631372 223970 632512 224026
rect 631311 223968 632512 223970
rect 631311 223965 631377 223968
rect 632506 223966 632512 223968
rect 632576 223966 632582 224030
rect 632698 223966 632704 224030
rect 632768 224028 632774 224030
rect 633519 224028 633585 224031
rect 632768 224026 633585 224028
rect 632768 223970 633524 224026
rect 633580 223970 633585 224026
rect 632768 223968 633585 223970
rect 632768 223966 632774 223968
rect 633519 223965 633585 223968
rect 631599 223880 631665 223883
rect 632367 223882 632433 223883
rect 632122 223880 632128 223882
rect 631599 223878 632128 223880
rect 631599 223822 631604 223878
rect 631660 223822 632128 223878
rect 631599 223820 632128 223822
rect 631599 223817 631665 223820
rect 632122 223818 632128 223820
rect 632192 223818 632198 223882
rect 632314 223818 632320 223882
rect 632384 223880 632433 223882
rect 632751 223880 632817 223883
rect 632890 223880 632896 223882
rect 632384 223878 632476 223880
rect 632428 223822 632476 223878
rect 632384 223820 632476 223822
rect 632751 223878 632896 223880
rect 632751 223822 632756 223878
rect 632812 223822 632896 223878
rect 632751 223820 632896 223822
rect 632384 223818 632433 223820
rect 632367 223817 632433 223818
rect 632751 223817 632817 223820
rect 632890 223818 632896 223820
rect 632960 223818 632966 223882
rect 633135 223880 633201 223883
rect 633274 223880 633280 223882
rect 633135 223878 633280 223880
rect 633135 223822 633140 223878
rect 633196 223822 633280 223878
rect 633135 223820 633280 223822
rect 633135 223817 633201 223820
rect 633274 223818 633280 223820
rect 633344 223818 633350 223882
rect 676866 223735 676926 223850
rect 676815 223730 676926 223735
rect 676815 223674 676820 223730
rect 676876 223674 676926 223730
rect 676815 223672 676926 223674
rect 676815 223669 676881 223672
rect 480834 223080 495294 223140
rect 447872 222932 460926 222992
rect 447872 222930 447878 222932
rect 145743 222844 145809 222847
rect 140832 222842 145809 222844
rect 140832 222786 145748 222842
rect 145804 222786 145809 222842
rect 140832 222784 145809 222786
rect 145743 222781 145809 222784
rect 362746 222782 362752 222846
rect 362816 222844 362822 222846
rect 440122 222844 440128 222846
rect 362816 222784 440128 222844
rect 362816 222782 362822 222784
rect 440122 222782 440128 222784
rect 440192 222782 440198 222846
rect 204975 222696 205041 222699
rect 207226 222696 207232 222698
rect 204975 222694 207232 222696
rect 204975 222638 204980 222694
rect 205036 222638 207232 222694
rect 204975 222636 207232 222638
rect 204975 222633 205041 222636
rect 207226 222634 207232 222636
rect 207296 222634 207302 222698
rect 349306 222634 349312 222698
rect 349376 222696 349382 222698
rect 440890 222696 440896 222698
rect 349376 222636 440896 222696
rect 349376 222634 349382 222636
rect 440890 222634 440896 222636
rect 440960 222634 440966 222698
rect 674554 222486 674560 222550
rect 674624 222548 674630 222550
rect 674754 222548 674814 223110
rect 674624 222488 674814 222548
rect 674624 222486 674630 222488
rect 639663 222400 639729 222403
rect 641007 222400 641073 222403
rect 634464 222398 641073 222400
rect 199791 222104 199857 222107
rect 200271 222104 200337 222107
rect 204546 222104 204606 222370
rect 634464 222342 639668 222398
rect 639724 222342 641012 222398
rect 641068 222342 641073 222398
rect 634464 222340 641073 222342
rect 639663 222337 639729 222340
rect 641007 222337 641073 222340
rect 199791 222102 204606 222104
rect 199791 222046 199796 222102
rect 199852 222046 200276 222102
rect 200332 222046 204606 222102
rect 199791 222044 204606 222046
rect 674511 222104 674577 222107
rect 674754 222104 674814 222222
rect 674511 222102 674814 222104
rect 674511 222046 674516 222102
rect 674572 222046 674814 222102
rect 674511 222044 674814 222046
rect 199791 222041 199857 222044
rect 200271 222041 200337 222044
rect 674511 222041 674577 222044
rect 199695 221808 199761 221811
rect 200463 221808 200529 221811
rect 204546 221808 204606 221852
rect 199695 221806 204606 221808
rect 199695 221750 199700 221806
rect 199756 221750 200468 221806
rect 200524 221750 204606 221806
rect 199695 221748 204606 221750
rect 634434 221808 634494 221852
rect 639375 221808 639441 221811
rect 640719 221808 640785 221811
rect 634434 221806 640785 221808
rect 634434 221750 639380 221806
rect 639436 221750 640724 221806
rect 640780 221750 640785 221806
rect 634434 221748 640785 221750
rect 199695 221745 199761 221748
rect 200463 221745 200529 221748
rect 639375 221745 639441 221748
rect 640719 221745 640785 221748
rect 140802 221364 140862 221556
rect 144111 221364 144177 221367
rect 140802 221362 144177 221364
rect 140802 221306 144116 221362
rect 144172 221306 144177 221362
rect 140802 221304 144177 221306
rect 144111 221301 144177 221304
rect 200175 221364 200241 221367
rect 201231 221364 201297 221367
rect 639855 221364 639921 221367
rect 641295 221364 641361 221367
rect 200175 221362 204576 221364
rect 200175 221306 200180 221362
rect 200236 221306 201236 221362
rect 201292 221306 204576 221362
rect 200175 221304 204576 221306
rect 634464 221362 641361 221364
rect 634464 221306 639860 221362
rect 639916 221306 641300 221362
rect 641356 221306 641361 221362
rect 634464 221304 641361 221306
rect 200175 221301 200241 221304
rect 201231 221301 201297 221304
rect 639855 221301 639921 221304
rect 641295 221301 641361 221304
rect 674946 221219 675006 221482
rect 674946 221214 675057 221219
rect 674946 221158 674996 221214
rect 675052 221158 675057 221214
rect 674946 221156 675057 221158
rect 674991 221153 675057 221156
rect 42351 221068 42417 221071
rect 42306 221066 42417 221068
rect 42306 221010 42356 221066
rect 42412 221010 42417 221066
rect 42306 221005 42417 221010
rect 674607 221068 674673 221071
rect 675322 221068 675328 221070
rect 674607 221066 675328 221068
rect 674607 221010 674612 221066
rect 674668 221010 675328 221066
rect 674607 221008 675328 221010
rect 674607 221005 674673 221008
rect 675322 221006 675328 221008
rect 675392 221006 675398 221070
rect 42306 220890 42366 221005
rect 200367 220772 200433 220775
rect 201327 220772 201393 220775
rect 639951 220772 640017 220775
rect 641295 220772 641361 220775
rect 200367 220770 204576 220772
rect 200367 220714 200372 220770
rect 200428 220714 201332 220770
rect 201388 220714 204576 220770
rect 200367 220712 204576 220714
rect 634464 220770 641361 220772
rect 634464 220714 639956 220770
rect 640012 220714 641300 220770
rect 641356 220714 641361 220770
rect 634464 220712 641361 220714
rect 200367 220709 200433 220712
rect 201327 220709 201393 220712
rect 639951 220709 640017 220712
rect 641295 220709 641361 220712
rect 42351 220328 42417 220331
rect 42306 220326 42417 220328
rect 42306 220270 42356 220326
rect 42412 220270 42417 220326
rect 42306 220265 42417 220270
rect 42306 220076 42366 220265
rect 140802 220032 140862 220510
rect 144015 220032 144081 220035
rect 140802 220030 144081 220032
rect 140802 219974 144020 220030
rect 144076 219974 144081 220030
rect 140802 219972 144081 219974
rect 144015 219969 144081 219972
rect 200559 219884 200625 219887
rect 201135 219884 201201 219887
rect 204546 219884 204606 220224
rect 675138 220182 675198 220742
rect 675130 220118 675136 220182
rect 675200 220118 675206 220182
rect 674362 219970 674368 220034
rect 674432 220032 674438 220034
rect 674432 219972 674784 220032
rect 674432 219970 674438 219972
rect 200559 219882 204606 219884
rect 200559 219826 200564 219882
rect 200620 219826 201140 219882
rect 201196 219826 204606 219882
rect 200559 219824 204606 219826
rect 200559 219821 200625 219824
rect 201135 219821 201201 219824
rect 200751 219736 200817 219739
rect 200751 219734 204576 219736
rect 200751 219678 200756 219734
rect 200812 219678 204576 219734
rect 200751 219676 204576 219678
rect 200751 219673 200817 219676
rect 42351 219440 42417 219443
rect 42306 219438 42417 219440
rect 42306 219382 42356 219438
rect 42412 219382 42417 219438
rect 42306 219377 42417 219382
rect 42306 219262 42366 219377
rect 145839 219292 145905 219295
rect 140832 219290 145905 219292
rect 140832 219234 145844 219290
rect 145900 219234 145905 219290
rect 140832 219232 145905 219234
rect 145839 219229 145905 219232
rect 198735 219144 198801 219147
rect 198735 219142 204576 219144
rect 198735 219086 198740 219142
rect 198796 219086 204576 219142
rect 198735 219084 204576 219086
rect 198735 219081 198801 219084
rect 675138 218999 675198 219114
rect 675138 218994 675249 218999
rect 675138 218938 675188 218994
rect 675244 218938 675249 218994
rect 675138 218936 675249 218938
rect 675183 218933 675249 218936
rect 198735 218700 198801 218703
rect 198735 218698 204606 218700
rect 198735 218642 198740 218698
rect 198796 218642 204606 218698
rect 198735 218640 204606 218642
rect 198735 218637 198801 218640
rect 204546 218596 204606 218640
rect 675138 218111 675198 218374
rect 144015 218108 144081 218111
rect 140832 218106 144081 218108
rect 140832 218050 144020 218106
rect 144076 218050 144081 218106
rect 140832 218048 144081 218050
rect 144015 218045 144081 218048
rect 199023 218108 199089 218111
rect 199023 218106 204576 218108
rect 199023 218050 199028 218106
rect 199084 218050 204576 218106
rect 199023 218048 204576 218050
rect 675087 218106 675198 218111
rect 675087 218050 675092 218106
rect 675148 218050 675198 218106
rect 675087 218048 675198 218050
rect 199023 218045 199089 218048
rect 675087 218045 675153 218048
rect 43599 217664 43665 217667
rect 42336 217662 43665 217664
rect 42336 217606 43604 217662
rect 43660 217606 43665 217662
rect 42336 217604 43665 217606
rect 43599 217601 43665 217604
rect 198831 217516 198897 217519
rect 674415 217516 674481 217519
rect 198831 217514 204576 217516
rect 198831 217458 198836 217514
rect 198892 217458 204576 217514
rect 198831 217456 204576 217458
rect 674415 217514 674784 217516
rect 674415 217458 674420 217514
rect 674476 217458 674784 217514
rect 674415 217456 674784 217458
rect 198831 217453 198897 217456
rect 674415 217453 674481 217456
rect 198927 217368 198993 217371
rect 198927 217366 204606 217368
rect 198927 217310 198932 217366
rect 198988 217310 204606 217366
rect 198927 217308 204606 217310
rect 198927 217305 198993 217308
rect 204546 216968 204606 217308
rect 43311 216924 43377 216927
rect 42336 216922 43377 216924
rect 42336 216866 43316 216922
rect 43372 216866 43377 216922
rect 42336 216864 43377 216866
rect 43311 216861 43377 216864
rect 140802 216332 140862 216820
rect 198735 216480 198801 216483
rect 198735 216478 204576 216480
rect 198735 216422 198740 216478
rect 198796 216422 204576 216478
rect 198735 216420 204576 216422
rect 198735 216417 198801 216420
rect 145935 216332 146001 216335
rect 674946 216334 675006 216746
rect 140802 216330 146001 216332
rect 140802 216274 145940 216330
rect 145996 216274 146001 216330
rect 140802 216272 146001 216274
rect 145935 216269 146001 216272
rect 674938 216270 674944 216334
rect 675008 216270 675014 216334
rect 43407 216184 43473 216187
rect 42336 216182 43473 216184
rect 42336 216126 43412 216182
rect 43468 216126 43473 216182
rect 42336 216124 43473 216126
rect 43407 216121 43473 216124
rect 674127 216036 674193 216039
rect 674127 216034 674784 216036
rect 674127 215978 674132 216034
rect 674188 215978 674784 216034
rect 674127 215976 674784 215978
rect 674127 215973 674193 215976
rect 198735 215888 198801 215891
rect 198735 215886 204576 215888
rect 198735 215830 198740 215886
rect 198796 215830 204576 215886
rect 198735 215828 204576 215830
rect 198735 215825 198801 215828
rect 198831 215740 198897 215743
rect 198831 215738 204606 215740
rect 198831 215682 198836 215738
rect 198892 215682 204606 215738
rect 198831 215680 204606 215682
rect 198831 215677 198897 215680
rect 146511 215592 146577 215595
rect 140832 215590 146577 215592
rect 140832 215534 146516 215590
rect 146572 215534 146577 215590
rect 140832 215532 146577 215534
rect 146511 215529 146577 215532
rect 204546 215340 204606 215680
rect 40578 214706 40638 215266
rect 674946 215003 675006 215192
rect 674895 214998 675006 215003
rect 674895 214942 674900 214998
rect 674956 214942 675006 214998
rect 674895 214940 675006 214942
rect 674895 214937 674961 214940
rect 198735 214852 198801 214855
rect 198735 214850 204576 214852
rect 198735 214794 198740 214850
rect 198796 214794 204576 214850
rect 198735 214792 204576 214794
rect 198735 214789 198801 214792
rect 40570 214642 40576 214706
rect 40640 214642 40646 214706
rect 41922 213967 41982 214526
rect 144015 214408 144081 214411
rect 140832 214406 144081 214408
rect 140832 214350 144020 214406
rect 144076 214350 144081 214406
rect 140832 214348 144081 214350
rect 144015 214345 144081 214348
rect 674754 214263 674814 214378
rect 198831 214260 198897 214263
rect 198831 214258 204576 214260
rect 198831 214202 198836 214258
rect 198892 214202 204576 214258
rect 198831 214200 204576 214202
rect 674754 214258 674865 214263
rect 674754 214202 674804 214258
rect 674860 214202 674865 214258
rect 674754 214200 674865 214202
rect 198831 214197 198897 214200
rect 674799 214197 674865 214200
rect 198927 214112 198993 214115
rect 198927 214110 204606 214112
rect 198927 214054 198932 214110
rect 198988 214054 204606 214110
rect 198927 214052 204606 214054
rect 198927 214049 198993 214052
rect 41871 213962 41982 213967
rect 41871 213906 41876 213962
rect 41932 213906 41982 213962
rect 41871 213904 41982 213906
rect 41871 213901 41937 213904
rect 204546 213712 204606 214052
rect 40386 213226 40446 213638
rect 674754 213375 674814 213564
rect 146031 213372 146097 213375
rect 140832 213370 146097 213372
rect 140832 213314 146036 213370
rect 146092 213314 146097 213370
rect 140832 213312 146097 213314
rect 146031 213309 146097 213312
rect 674703 213370 674814 213375
rect 674703 213314 674708 213370
rect 674764 213314 674814 213370
rect 674703 213312 674814 213314
rect 674703 213309 674769 213312
rect 40378 213162 40384 213226
rect 40448 213162 40454 213226
rect 199023 213224 199089 213227
rect 199023 213222 204576 213224
rect 199023 213166 199028 213222
rect 199084 213166 204576 213222
rect 199023 213164 204576 213166
rect 199023 213161 199089 213164
rect 40962 212486 41022 212898
rect 198735 212632 198801 212635
rect 198735 212630 204576 212632
rect 198735 212574 198740 212630
rect 198796 212574 204576 212630
rect 198735 212572 204576 212574
rect 198735 212569 198801 212572
rect 40954 212422 40960 212486
rect 41024 212422 41030 212486
rect 679746 212191 679806 212750
rect 679695 212186 679806 212191
rect 41154 211598 41214 212158
rect 679695 212130 679700 212186
rect 679756 212130 679806 212186
rect 679695 212128 679806 212130
rect 679695 212125 679761 212128
rect 41146 211534 41152 211598
rect 41216 211534 41222 211598
rect 140802 211596 140862 212078
rect 146127 211596 146193 211599
rect 140802 211594 146193 211596
rect 140802 211538 146132 211594
rect 146188 211538 146193 211594
rect 140802 211536 146193 211538
rect 146127 211533 146193 211536
rect 679695 211448 679761 211451
rect 679695 211446 679806 211448
rect 37314 210859 37374 211418
rect 679695 211390 679700 211446
rect 679756 211390 679806 211446
rect 679695 211385 679806 211390
rect 679746 211270 679806 211385
rect 639759 211004 639825 211007
rect 634464 211002 639825 211004
rect 634464 210946 639764 211002
rect 639820 210946 639825 211002
rect 634464 210944 639825 210946
rect 639759 210941 639825 210944
rect 37314 210854 37425 210859
rect 144015 210856 144081 210859
rect 37314 210798 37364 210854
rect 37420 210798 37425 210854
rect 37314 210796 37425 210798
rect 140832 210854 144081 210856
rect 140832 210798 144020 210854
rect 144076 210798 144081 210854
rect 140832 210796 144081 210798
rect 37359 210793 37425 210796
rect 144015 210793 144081 210796
rect 40770 210414 40830 210530
rect 40762 210350 40768 210414
rect 40832 210350 40838 210414
rect 674746 210054 674752 210118
rect 674816 210116 674822 210118
rect 679791 210116 679857 210119
rect 674816 210114 679857 210116
rect 674816 210058 679796 210114
rect 679852 210058 679857 210114
rect 674816 210056 679857 210058
rect 674816 210054 674822 210056
rect 679791 210053 679857 210056
rect 41922 209231 41982 209790
rect 41922 209226 42033 209231
rect 41922 209170 41972 209226
rect 42028 209170 42033 209226
rect 41922 209168 42033 209170
rect 41967 209165 42033 209168
rect 140802 209080 140862 209630
rect 144015 209080 144081 209083
rect 140802 209078 144081 209080
rect 140802 209022 144020 209078
rect 144076 209022 144081 209078
rect 140802 209020 144081 209022
rect 144015 209017 144081 209020
rect 42114 208343 42174 208902
rect 42063 208338 42174 208343
rect 42063 208282 42068 208338
rect 42124 208282 42174 208338
rect 42063 208280 42174 208282
rect 42063 208277 42129 208280
rect 42735 208118 42801 208121
rect 42336 208116 42801 208118
rect 42336 208060 42740 208116
rect 42796 208060 42801 208116
rect 42336 208058 42801 208060
rect 42735 208055 42801 208058
rect 140802 207896 140862 208384
rect 146223 207896 146289 207899
rect 140802 207894 146289 207896
rect 140802 207838 146228 207894
rect 146284 207838 146289 207894
rect 140802 207836 146289 207838
rect 146223 207833 146289 207836
rect 43023 207452 43089 207455
rect 42336 207450 43089 207452
rect 42336 207394 43028 207450
rect 43084 207394 43089 207450
rect 42336 207392 43089 207394
rect 43023 207389 43089 207392
rect 146799 207156 146865 207159
rect 140832 207154 146865 207156
rect 140832 207098 146804 207154
rect 146860 207098 146865 207154
rect 140832 207096 146865 207098
rect 146799 207093 146865 207096
rect 41730 206123 41790 206608
rect 676090 206206 676096 206270
rect 676160 206268 676166 206270
rect 676815 206268 676881 206271
rect 676160 206266 676881 206268
rect 676160 206210 676820 206266
rect 676876 206210 676881 206266
rect 676160 206208 676881 206210
rect 676160 206206 676166 206208
rect 676815 206205 676881 206208
rect 41679 206118 41790 206123
rect 146319 206120 146385 206123
rect 41679 206062 41684 206118
rect 41740 206062 41790 206118
rect 41679 206060 41790 206062
rect 140832 206118 146385 206120
rect 140832 206062 146324 206118
rect 146380 206062 146385 206118
rect 140832 206060 146385 206062
rect 41679 206057 41745 206060
rect 146319 206057 146385 206060
rect 43119 205824 43185 205827
rect 42336 205822 43185 205824
rect 42336 205766 43124 205822
rect 43180 205766 43185 205822
rect 42336 205764 43185 205766
rect 43119 205761 43185 205764
rect 42306 204640 42366 204980
rect 146799 204936 146865 204939
rect 140832 204934 146865 204936
rect 140832 204878 146804 204934
rect 146860 204878 146865 204934
rect 140832 204876 146865 204878
rect 146799 204873 146865 204876
rect 43023 204640 43089 204643
rect 42306 204638 43089 204640
rect 42306 204582 43028 204638
rect 43084 204582 43089 204638
rect 42306 204580 43089 204582
rect 43023 204577 43089 204580
rect 675759 204492 675825 204495
rect 676090 204492 676096 204494
rect 675759 204490 676096 204492
rect 675759 204434 675764 204490
rect 675820 204434 676096 204490
rect 675759 204432 676096 204434
rect 675759 204429 675825 204432
rect 676090 204430 676096 204432
rect 676160 204430 676166 204494
rect 42351 204344 42417 204347
rect 42306 204342 42417 204344
rect 42306 204286 42356 204342
rect 42412 204286 42417 204342
rect 42306 204281 42417 204286
rect 42306 204166 42366 204281
rect 140802 203456 140862 203646
rect 144975 203456 145041 203459
rect 140802 203454 145041 203456
rect 140802 203398 144980 203454
rect 145036 203398 145041 203454
rect 140802 203396 145041 203398
rect 144975 203393 145041 203396
rect 42351 202864 42417 202867
rect 42306 202862 42417 202864
rect 42306 202806 42356 202862
rect 42412 202806 42417 202862
rect 42306 202801 42417 202806
rect 200367 202864 200433 202867
rect 200943 202864 201009 202867
rect 200367 202862 204576 202864
rect 200367 202806 200372 202862
rect 200428 202806 200948 202862
rect 201004 202806 204576 202862
rect 200367 202804 204576 202806
rect 200367 202801 200433 202804
rect 200943 202801 201009 202804
rect 42306 202686 42366 202801
rect 146415 202420 146481 202423
rect 140832 202418 146481 202420
rect 140832 202362 146420 202418
rect 146476 202362 146481 202418
rect 140832 202360 146481 202362
rect 146415 202357 146481 202360
rect 674607 201680 674673 201683
rect 675514 201680 675520 201682
rect 674607 201678 675520 201680
rect 674607 201622 674612 201678
rect 674668 201622 675520 201678
rect 674607 201620 675520 201622
rect 674607 201617 674673 201620
rect 675514 201618 675520 201620
rect 675584 201618 675590 201682
rect 140802 200644 140862 201198
rect 144975 200644 145041 200647
rect 140802 200642 145041 200644
rect 140802 200586 144980 200642
rect 145036 200586 145041 200642
rect 140802 200584 145041 200586
rect 144975 200581 145041 200584
rect 675471 200054 675537 200055
rect 675471 200052 675520 200054
rect 675428 200050 675520 200052
rect 675428 199994 675476 200050
rect 675428 199992 675520 199994
rect 675471 199990 675520 199992
rect 675584 199990 675590 200054
rect 675471 199989 675537 199990
rect 140802 199460 140862 199948
rect 144399 199460 144465 199463
rect 675375 199462 675441 199463
rect 140802 199458 144465 199460
rect 140802 199402 144404 199458
rect 144460 199402 144465 199458
rect 140802 199400 144465 199402
rect 144399 199397 144465 199400
rect 675322 199398 675328 199462
rect 675392 199460 675441 199462
rect 675392 199458 675484 199460
rect 675436 199402 675484 199458
rect 675392 199400 675484 199402
rect 675392 199398 675441 199400
rect 675375 199397 675441 199398
rect 146703 198720 146769 198723
rect 140832 198718 146769 198720
rect 140832 198662 146708 198718
rect 146764 198662 146769 198718
rect 140832 198660 146769 198662
rect 146703 198657 146769 198660
rect 675130 198362 675136 198426
rect 675200 198424 675206 198426
rect 675471 198424 675537 198427
rect 675200 198422 675537 198424
rect 675200 198366 675476 198422
rect 675532 198366 675537 198422
rect 675200 198364 675537 198366
rect 675200 198362 675206 198364
rect 675471 198361 675537 198364
rect 41679 197684 41745 197687
rect 42490 197684 42496 197686
rect 41679 197682 42496 197684
rect 41679 197626 41684 197682
rect 41740 197626 42496 197682
rect 41679 197624 42496 197626
rect 41679 197621 41745 197624
rect 42490 197622 42496 197624
rect 42560 197622 42566 197686
rect 145263 197684 145329 197687
rect 140832 197682 145329 197684
rect 140832 197626 145268 197682
rect 145324 197626 145329 197682
rect 140832 197624 145329 197626
rect 145263 197621 145329 197624
rect 140802 196204 140862 196396
rect 144975 196204 145041 196207
rect 140802 196202 145041 196204
rect 140802 196146 144980 196202
rect 145036 196146 145041 196202
rect 140802 196144 145041 196146
rect 144975 196141 145041 196144
rect 42490 195698 42496 195762
rect 42560 195760 42566 195762
rect 42639 195760 42705 195763
rect 42560 195758 42705 195760
rect 42560 195702 42644 195758
rect 42700 195702 42705 195758
rect 42560 195700 42705 195702
rect 42560 195698 42566 195700
rect 42639 195697 42705 195700
rect 674938 195254 674944 195318
rect 675008 195316 675014 195318
rect 675471 195316 675537 195319
rect 675008 195314 675537 195316
rect 675008 195258 675476 195314
rect 675532 195258 675537 195314
rect 675008 195256 675537 195258
rect 675008 195254 675014 195256
rect 675471 195253 675537 195256
rect 140802 194724 140862 195212
rect 146799 194724 146865 194727
rect 140802 194722 146865 194724
rect 140802 194666 146804 194722
rect 146860 194666 146865 194722
rect 140802 194664 146865 194666
rect 146799 194661 146865 194664
rect 144591 193984 144657 193987
rect 140832 193982 144657 193984
rect 140832 193926 144596 193982
rect 144652 193926 144657 193982
rect 140832 193924 144657 193926
rect 144591 193921 144657 193924
rect 674554 193478 674560 193542
rect 674624 193540 674630 193542
rect 675375 193540 675441 193543
rect 674624 193538 675441 193540
rect 674624 193482 675380 193538
rect 675436 193482 675441 193538
rect 674624 193480 675441 193482
rect 674624 193478 674630 193480
rect 675375 193477 675441 193480
rect 675087 193244 675153 193247
rect 675514 193244 675520 193246
rect 675087 193242 675520 193244
rect 675087 193186 675092 193242
rect 675148 193186 675520 193242
rect 675087 193184 675520 193186
rect 675087 193181 675153 193184
rect 675514 193182 675520 193184
rect 675584 193182 675590 193246
rect 675183 193096 675249 193099
rect 675322 193096 675328 193098
rect 675183 193094 675328 193096
rect 675183 193038 675188 193094
rect 675244 193038 675328 193094
rect 675183 193036 675328 193038
rect 675183 193033 675249 193036
rect 675322 193034 675328 193036
rect 675392 193034 675398 193098
rect 140802 192208 140862 192766
rect 144303 192208 144369 192211
rect 140802 192206 144369 192208
rect 140802 192150 144308 192206
rect 144364 192150 144369 192206
rect 140802 192148 144369 192150
rect 144303 192145 144369 192148
rect 674362 191554 674368 191618
rect 674432 191616 674438 191618
rect 675375 191616 675441 191619
rect 674432 191614 675441 191616
rect 674432 191558 675380 191614
rect 675436 191558 675441 191614
rect 674432 191556 675441 191558
rect 674432 191554 674438 191556
rect 675375 191553 675441 191556
rect 140802 191024 140862 191512
rect 144879 191024 144945 191027
rect 140802 191022 144945 191024
rect 140802 190966 144884 191022
rect 144940 190966 144945 191022
rect 140802 190964 144945 190966
rect 144879 190961 144945 190964
rect 146511 190432 146577 190435
rect 140832 190430 146577 190432
rect 140832 190374 146516 190430
rect 146572 190374 146577 190430
rect 140832 190372 146577 190374
rect 146511 190369 146577 190372
rect 41146 190074 41152 190138
rect 41216 190136 41222 190138
rect 41775 190136 41841 190139
rect 41216 190134 41841 190136
rect 41216 190078 41780 190134
rect 41836 190078 41841 190134
rect 41216 190076 41841 190078
rect 41216 190074 41222 190076
rect 41775 190073 41841 190076
rect 146799 189248 146865 189251
rect 140832 189246 146865 189248
rect 140832 189190 146804 189246
rect 146860 189190 146865 189246
rect 140832 189188 146865 189190
rect 146799 189185 146865 189188
rect 41967 189102 42033 189103
rect 41914 189100 41920 189102
rect 41876 189040 41920 189100
rect 41984 189098 42033 189102
rect 42028 189042 42033 189098
rect 41914 189038 41920 189040
rect 41984 189038 42033 189042
rect 41967 189037 42033 189038
rect 41775 188362 41841 188363
rect 41722 188298 41728 188362
rect 41792 188360 41841 188362
rect 41792 188358 41884 188360
rect 41836 188302 41884 188358
rect 41792 188300 41884 188302
rect 41792 188298 41841 188300
rect 41775 188297 41841 188298
rect 140802 187472 140862 187960
rect 145167 187472 145233 187475
rect 140802 187470 145233 187472
rect 140802 187414 145172 187470
rect 145228 187414 145233 187470
rect 140802 187412 145233 187414
rect 145167 187409 145233 187412
rect 140802 186288 140862 186776
rect 146607 186288 146673 186291
rect 140802 186286 146673 186288
rect 140802 186230 146612 186286
rect 146668 186230 146673 186286
rect 140802 186228 146673 186230
rect 146607 186225 146673 186228
rect 40954 185930 40960 185994
rect 41024 185992 41030 185994
rect 41775 185992 41841 185995
rect 41024 185990 41841 185992
rect 41024 185934 41780 185990
rect 41836 185934 41841 185990
rect 41024 185932 41841 185934
rect 41024 185930 41030 185932
rect 41775 185929 41841 185932
rect 146799 185548 146865 185551
rect 140832 185546 146865 185548
rect 140832 185490 146804 185546
rect 146860 185490 146865 185546
rect 140832 185488 146865 185490
rect 146799 185485 146865 185488
rect 674415 184512 674481 184515
rect 674415 184510 674784 184512
rect 674415 184454 674420 184510
rect 674476 184454 674784 184510
rect 674415 184452 674784 184454
rect 674415 184449 674481 184452
rect 145071 184364 145137 184367
rect 140832 184362 145137 184364
rect 140832 184306 145076 184362
rect 145132 184306 145137 184362
rect 140832 184304 145137 184306
rect 145071 184301 145137 184304
rect 40570 184154 40576 184218
rect 40640 184216 40646 184218
rect 41775 184216 41841 184219
rect 40640 184214 41841 184216
rect 40640 184158 41780 184214
rect 41836 184158 41841 184214
rect 40640 184156 41841 184158
rect 40640 184154 40646 184156
rect 41775 184153 41841 184156
rect 674703 183920 674769 183923
rect 674703 183918 674814 183920
rect 674703 183862 674708 183918
rect 674764 183862 674814 183918
rect 674703 183857 674814 183862
rect 674754 183668 674814 183857
rect 40762 183562 40768 183626
rect 40832 183624 40838 183626
rect 41775 183624 41841 183627
rect 40832 183622 41841 183624
rect 40832 183566 41780 183622
rect 41836 183566 41841 183622
rect 40832 183564 41841 183566
rect 40832 183562 40838 183564
rect 41775 183561 41841 183564
rect 40378 182822 40384 182886
rect 40448 182884 40454 182886
rect 41775 182884 41841 182887
rect 40448 182882 41841 182884
rect 40448 182826 41780 182882
rect 41836 182826 41841 182882
rect 40448 182824 41841 182826
rect 40448 182822 40454 182824
rect 41775 182821 41841 182824
rect 140802 182736 140862 183224
rect 674415 182884 674481 182887
rect 674415 182882 674784 182884
rect 674415 182826 674420 182882
rect 674476 182826 674784 182882
rect 674415 182824 674784 182826
rect 674415 182821 674481 182824
rect 144687 182736 144753 182739
rect 140802 182734 144753 182736
rect 140802 182678 144692 182734
rect 144748 182678 144753 182734
rect 140802 182676 144753 182678
rect 144687 182673 144753 182676
rect 674170 182008 674176 182072
rect 674240 182070 674246 182072
rect 674240 182010 674784 182070
rect 674240 182008 674246 182010
rect 146799 181996 146865 181999
rect 140832 181994 146865 181996
rect 140832 181938 146804 181994
rect 146860 181938 146865 181994
rect 140832 181936 146865 181938
rect 146799 181933 146865 181936
rect 200847 181406 200913 181407
rect 200847 181402 200896 181406
rect 200960 181404 200966 181406
rect 200847 181346 200852 181402
rect 200847 181342 200896 181346
rect 200960 181344 201004 181404
rect 200960 181342 200966 181344
rect 200847 181341 200913 181342
rect 674170 181194 674176 181258
rect 674240 181256 674246 181258
rect 674240 181196 674784 181256
rect 674240 181194 674246 181196
rect 674746 180898 674752 180962
rect 674816 180898 674822 180962
rect 144879 180812 144945 180815
rect 140832 180810 144945 180812
rect 140832 180754 144884 180810
rect 144940 180754 144945 180810
rect 140832 180752 144945 180754
rect 144879 180749 144945 180752
rect 674362 180454 674368 180518
rect 674432 180516 674438 180518
rect 674754 180516 674814 180898
rect 674432 180486 674814 180516
rect 674432 180456 674784 180486
rect 674432 180454 674438 180456
rect 673978 179714 673984 179778
rect 674048 179776 674054 179778
rect 674048 179716 674784 179776
rect 674048 179714 674054 179716
rect 140802 179184 140862 179524
rect 144015 179184 144081 179187
rect 140802 179182 144081 179184
rect 140802 179126 144020 179182
rect 144076 179126 144081 179182
rect 140802 179124 144081 179126
rect 144015 179121 144081 179124
rect 676866 178743 676926 178858
rect 676866 178738 676977 178743
rect 676866 178682 676916 178738
rect 676972 178682 676977 178738
rect 676866 178680 676977 178682
rect 676911 178677 676977 178680
rect 140802 177852 140862 178340
rect 144687 177852 144753 177855
rect 140802 177850 144753 177852
rect 140802 177794 144692 177850
rect 144748 177794 144753 177850
rect 140802 177792 144753 177794
rect 144687 177789 144753 177792
rect 674754 177558 674814 178118
rect 674746 177494 674752 177558
rect 674816 177494 674822 177558
rect 31738 177050 31744 177114
rect 31808 177112 31814 177114
rect 42735 177112 42801 177115
rect 144495 177112 144561 177115
rect 31808 177110 42801 177112
rect 31808 177054 42740 177110
rect 42796 177054 42801 177110
rect 31808 177052 42801 177054
rect 140832 177110 144561 177112
rect 140832 177054 144500 177110
rect 144556 177054 144561 177110
rect 140832 177052 144561 177054
rect 31808 177050 31814 177052
rect 42735 177049 42801 177052
rect 144495 177049 144561 177052
rect 674511 177112 674577 177115
rect 674754 177112 674814 177230
rect 674511 177110 674814 177112
rect 674511 177054 674516 177110
rect 674572 177054 674814 177110
rect 674511 177052 674814 177054
rect 674511 177049 674577 177052
rect 676866 176227 676926 176490
rect 676815 176222 676926 176227
rect 676815 176166 676820 176222
rect 676876 176166 676926 176222
rect 676815 176164 676926 176166
rect 676815 176161 676881 176164
rect 144975 175928 145041 175931
rect 140832 175926 145041 175928
rect 140832 175870 144980 175926
rect 145036 175870 145041 175926
rect 140832 175868 145041 175870
rect 144975 175865 145041 175868
rect 677058 175635 677118 175750
rect 677007 175630 677118 175635
rect 677007 175574 677012 175630
rect 677068 175574 677118 175630
rect 677007 175572 677118 175574
rect 677007 175569 677073 175572
rect 140802 174300 140862 174788
rect 674554 174386 674560 174450
rect 674624 174448 674630 174450
rect 674754 174448 674814 175010
rect 674624 174388 674814 174448
rect 674624 174386 674630 174388
rect 144975 174300 145041 174303
rect 140802 174298 145041 174300
rect 140802 174242 144980 174298
rect 145036 174242 145041 174298
rect 140802 174240 145041 174242
rect 144975 174237 145041 174240
rect 675714 174007 675774 174122
rect 675663 174002 675774 174007
rect 675663 173946 675668 174002
rect 675724 173946 675774 174002
rect 675663 173944 675774 173946
rect 675663 173941 675729 173944
rect 144783 173560 144849 173563
rect 140832 173558 144849 173560
rect 140832 173502 144788 173558
rect 144844 173502 144849 173558
rect 140832 173500 144849 173502
rect 144783 173497 144849 173500
rect 674946 173119 675006 173382
rect 674895 173114 675006 173119
rect 674895 173058 674900 173114
rect 674956 173058 675006 173114
rect 674895 173056 675006 173058
rect 674895 173053 674961 173056
rect 674946 172379 675006 172494
rect 144399 172376 144465 172379
rect 140832 172374 144465 172376
rect 140832 172318 144404 172374
rect 144460 172318 144465 172374
rect 140832 172316 144465 172318
rect 674946 172374 675057 172379
rect 674946 172318 674996 172374
rect 675052 172318 675057 172374
rect 674946 172316 675057 172318
rect 144399 172313 144465 172316
rect 674991 172313 675057 172316
rect 674946 171342 675006 171754
rect 674938 171278 674944 171342
rect 675008 171278 675014 171342
rect 140802 170600 140862 171088
rect 674031 171044 674097 171047
rect 674031 171042 674784 171044
rect 674031 170986 674036 171042
rect 674092 170986 674784 171042
rect 674031 170984 674784 170986
rect 674031 170981 674097 170984
rect 144975 170600 145041 170603
rect 140802 170598 145041 170600
rect 140802 170542 144980 170598
rect 145036 170542 145041 170598
rect 140802 170540 145041 170542
rect 144975 170537 145041 170540
rect 675138 170011 675198 170200
rect 144591 170008 144657 170011
rect 140832 170006 144657 170008
rect 140832 169950 144596 170006
rect 144652 169950 144657 170006
rect 140832 169948 144657 169950
rect 144591 169945 144657 169948
rect 675087 170006 675198 170011
rect 675087 169950 675092 170006
rect 675148 169950 675198 170006
rect 675087 169948 675198 169950
rect 675087 169945 675153 169948
rect 674223 169416 674289 169419
rect 674223 169414 674784 169416
rect 674223 169358 674228 169414
rect 674284 169358 674784 169414
rect 674223 169356 674784 169358
rect 674223 169353 674289 169356
rect 144975 168676 145041 168679
rect 140832 168674 145041 168676
rect 140832 168618 144980 168674
rect 145036 168618 145041 168674
rect 140832 168616 145041 168618
rect 144975 168613 145041 168616
rect 674511 168380 674577 168383
rect 674754 168380 674814 168572
rect 674511 168378 674814 168380
rect 674511 168322 674516 168378
rect 674572 168322 674814 168378
rect 674511 168320 674814 168322
rect 674511 168317 674577 168320
rect 140802 167196 140862 167606
rect 674754 167347 674814 167758
rect 674703 167342 674814 167347
rect 674703 167286 674708 167342
rect 674764 167286 674814 167342
rect 674703 167284 674814 167286
rect 674703 167281 674769 167284
rect 144975 167196 145041 167199
rect 140802 167194 145041 167196
rect 140802 167138 144980 167194
rect 145036 167138 145041 167194
rect 140802 167136 145041 167138
rect 144975 167133 145041 167136
rect 200943 166902 201009 166903
rect 200890 166900 200896 166902
rect 200852 166840 200896 166900
rect 200960 166898 201009 166902
rect 642063 166900 642129 166903
rect 201004 166842 201009 166898
rect 200890 166838 200896 166840
rect 200960 166838 201009 166842
rect 634464 166898 642129 166900
rect 634464 166842 642068 166898
rect 642124 166842 642129 166898
rect 634464 166840 642129 166842
rect 200943 166837 201009 166838
rect 642063 166837 642129 166840
rect 674607 166752 674673 166755
rect 674754 166752 674814 166944
rect 674607 166750 674814 166752
rect 674607 166694 674612 166750
rect 674668 166694 674814 166750
rect 674607 166692 674814 166694
rect 674607 166689 674673 166692
rect 642159 166456 642225 166459
rect 634464 166454 642225 166456
rect 634464 166398 642164 166454
rect 642220 166398 642225 166454
rect 634464 166396 642225 166398
rect 642159 166393 642225 166396
rect 140802 165864 140862 166352
rect 144975 165864 145041 165867
rect 641487 165864 641553 165867
rect 140802 165862 145041 165864
rect 140802 165806 144980 165862
rect 145036 165806 145041 165862
rect 140802 165804 145041 165806
rect 634464 165862 641553 165864
rect 634464 165806 641492 165862
rect 641548 165806 641553 165862
rect 634464 165804 641553 165806
rect 144975 165801 145041 165804
rect 641487 165801 641553 165804
rect 674754 165719 674814 166278
rect 674703 165714 674814 165719
rect 674703 165658 674708 165714
rect 674764 165658 674814 165714
rect 674703 165656 674814 165658
rect 674703 165653 674769 165656
rect 140802 164680 140862 165158
rect 144015 164680 144081 164683
rect 140802 164678 144081 164680
rect 140802 164622 144020 164678
rect 144076 164622 144081 164678
rect 140802 164620 144081 164622
rect 144015 164617 144081 164620
rect 144303 163940 144369 163943
rect 140832 163938 144369 163940
rect 140832 163882 144308 163938
rect 144364 163882 144369 163938
rect 140832 163880 144369 163882
rect 144303 163877 144369 163880
rect 140802 162164 140862 162652
rect 144207 162164 144273 162167
rect 140802 162162 144273 162164
rect 140802 162106 144212 162162
rect 144268 162106 144273 162162
rect 140802 162104 144273 162106
rect 144207 162101 144273 162104
rect 144975 161572 145041 161575
rect 140832 161570 145041 161572
rect 140832 161514 144980 161570
rect 145036 161514 145041 161570
rect 140832 161512 145041 161514
rect 144975 161509 145041 161512
rect 675706 161362 675712 161426
rect 675776 161424 675782 161426
rect 677007 161424 677073 161427
rect 675776 161422 677073 161424
rect 675776 161366 677012 161422
rect 677068 161366 677073 161422
rect 675776 161364 677073 161366
rect 675776 161362 675782 161364
rect 677007 161361 677073 161364
rect 144303 160388 144369 160391
rect 140832 160386 144369 160388
rect 140832 160330 144308 160386
rect 144364 160330 144369 160386
rect 140832 160328 144369 160330
rect 144303 160325 144369 160328
rect 140802 158612 140862 159146
rect 144111 158612 144177 158615
rect 140802 158610 144177 158612
rect 140802 158554 144116 158610
rect 144172 158554 144177 158610
rect 140802 158552 144177 158554
rect 144111 158549 144177 158552
rect 140802 157428 140862 157916
rect 144495 157428 144561 157431
rect 140802 157426 144561 157428
rect 140802 157370 144500 157426
rect 144556 157370 144561 157426
rect 140802 157368 144561 157370
rect 144495 157365 144561 157368
rect 140802 156244 140862 156726
rect 144303 156244 144369 156247
rect 140802 156242 144369 156244
rect 140802 156186 144308 156242
rect 144364 156186 144369 156242
rect 140802 156184 144369 156186
rect 144303 156181 144369 156184
rect 144207 155504 144273 155507
rect 140832 155502 144273 155504
rect 140832 155446 144212 155502
rect 144268 155446 144273 155502
rect 140832 155444 144273 155446
rect 144207 155441 144273 155444
rect 675279 155210 675345 155211
rect 675279 155208 675328 155210
rect 675236 155206 675328 155208
rect 675236 155150 675284 155206
rect 675236 155148 675328 155150
rect 675279 155146 675328 155148
rect 675392 155146 675398 155210
rect 675279 155145 675345 155146
rect 675471 155062 675537 155063
rect 675471 155060 675520 155062
rect 675428 155058 675520 155060
rect 675428 155002 675476 155058
rect 675428 155000 675520 155002
rect 675471 154998 675520 155000
rect 675584 154998 675590 155062
rect 675471 154997 675537 154998
rect 140802 153728 140862 154278
rect 144303 153728 144369 153731
rect 140802 153726 144369 153728
rect 140802 153670 144308 153726
rect 144364 153670 144369 153726
rect 140802 153668 144369 153670
rect 144303 153665 144369 153668
rect 675759 153434 675825 153435
rect 675706 153370 675712 153434
rect 675776 153432 675825 153434
rect 675776 153430 675868 153432
rect 675820 153374 675868 153430
rect 675776 153372 675868 153374
rect 675776 153370 675825 153372
rect 675759 153369 675825 153370
rect 144495 153136 144561 153139
rect 140832 153134 144561 153136
rect 140832 153078 144500 153134
rect 144556 153078 144561 153134
rect 140832 153076 144561 153078
rect 144495 153073 144561 153076
rect 144495 151952 144561 151955
rect 140832 151950 144561 151952
rect 140832 151894 144500 151950
rect 144556 151894 144561 151950
rect 140832 151892 144561 151894
rect 144495 151889 144561 151892
rect 144303 150768 144369 150771
rect 140832 150766 144369 150768
rect 140832 150710 144308 150766
rect 144364 150710 144369 150766
rect 140832 150708 144369 150710
rect 144303 150705 144369 150708
rect 674938 150262 674944 150326
rect 675008 150324 675014 150326
rect 675471 150324 675537 150327
rect 675008 150322 675537 150324
rect 675008 150266 675476 150322
rect 675532 150266 675537 150322
rect 675008 150264 675537 150266
rect 675008 150262 675014 150264
rect 675471 150261 675537 150264
rect 640143 150028 640209 150031
rect 634464 150026 640209 150028
rect 634464 149970 640148 150026
rect 640204 149970 640209 150026
rect 634464 149968 640209 149970
rect 640143 149965 640209 149968
rect 140802 148992 140862 149480
rect 144207 148992 144273 148995
rect 140802 148990 144273 148992
rect 140802 148934 144212 148990
rect 144268 148934 144273 148990
rect 140802 148932 144273 148934
rect 144207 148929 144273 148932
rect 674746 148486 674752 148550
rect 674816 148548 674822 148550
rect 675471 148548 675537 148551
rect 674816 148546 675537 148548
rect 674816 148490 675476 148546
rect 675532 148490 675537 148546
rect 674816 148488 675537 148490
rect 674816 148486 674822 148488
rect 675471 148485 675537 148488
rect 140802 147808 140862 148294
rect 144303 147808 144369 147811
rect 140802 147806 144369 147808
rect 140802 147750 144308 147806
rect 144364 147750 144369 147806
rect 140802 147748 144369 147750
rect 144303 147745 144369 147748
rect 144495 147068 144561 147071
rect 140832 147066 144561 147068
rect 140832 147010 144500 147066
rect 144556 147010 144561 147066
rect 140832 147008 144561 147010
rect 144495 147005 144561 147008
rect 674554 146414 674560 146478
rect 674624 146476 674630 146478
rect 675375 146476 675441 146479
rect 674624 146474 675441 146476
rect 674624 146418 675380 146474
rect 675436 146418 675441 146474
rect 674624 146416 675441 146418
rect 674624 146414 674630 146416
rect 675375 146413 675441 146416
rect 140802 145292 140862 145846
rect 144303 145292 144369 145295
rect 140802 145290 144369 145292
rect 140802 145234 144308 145290
rect 144364 145234 144369 145290
rect 140802 145232 144369 145234
rect 144303 145229 144369 145232
rect 140802 144404 140862 144744
rect 144495 144404 144561 144407
rect 140802 144402 144561 144404
rect 140802 144346 144500 144402
rect 144556 144346 144561 144402
rect 140802 144344 144561 144346
rect 144495 144341 144561 144344
rect 144303 143516 144369 143519
rect 642159 143516 642225 143519
rect 140832 143514 144369 143516
rect 140832 143458 144308 143514
rect 144364 143458 144369 143514
rect 140832 143456 144369 143458
rect 634464 143514 642225 143516
rect 634464 143458 642164 143514
rect 642220 143458 642225 143514
rect 634464 143456 642225 143458
rect 144303 143453 144369 143456
rect 642159 143453 642225 143456
rect 674319 142778 674385 142779
rect 674319 142774 674368 142778
rect 674432 142776 674438 142778
rect 674319 142718 674324 142774
rect 674319 142714 674368 142718
rect 674432 142716 674476 142776
rect 674432 142714 674438 142716
rect 674319 142713 674385 142714
rect 144495 142332 144561 142335
rect 140832 142330 144561 142332
rect 140832 142274 144500 142330
rect 144556 142274 144561 142330
rect 140832 142272 144561 142274
rect 144495 142269 144561 142272
rect 140802 140556 140862 141044
rect 144303 140556 144369 140559
rect 140802 140554 144369 140556
rect 140802 140498 144308 140554
rect 144364 140498 144369 140554
rect 140802 140496 144369 140498
rect 144303 140493 144369 140496
rect 140802 139372 140862 139860
rect 144207 139372 144273 139375
rect 140802 139370 144273 139372
rect 140802 139314 144212 139370
rect 144268 139314 144273 139370
rect 140802 139312 144273 139314
rect 144207 139309 144273 139312
rect 674754 138783 674814 139342
rect 674703 138778 674814 138783
rect 674703 138722 674708 138778
rect 674764 138722 674814 138778
rect 674703 138720 674814 138722
rect 674703 138717 674769 138720
rect 144495 138632 144561 138635
rect 140832 138630 144561 138632
rect 140832 138574 144500 138630
rect 144556 138574 144561 138630
rect 140832 138572 144561 138574
rect 144495 138569 144561 138572
rect 674415 138484 674481 138487
rect 674415 138482 674784 138484
rect 674415 138426 674420 138482
rect 674476 138426 674784 138482
rect 674415 138424 674784 138426
rect 674415 138421 674481 138424
rect 140802 137004 140862 137492
rect 674754 137155 674814 137640
rect 674703 137150 674814 137155
rect 674703 137094 674708 137150
rect 674764 137094 674814 137150
rect 674703 137092 674814 137094
rect 674703 137089 674769 137092
rect 144207 137004 144273 137007
rect 140802 137002 144273 137004
rect 140802 136946 144212 137002
rect 144268 136946 144273 137002
rect 140802 136944 144273 136946
rect 144207 136941 144273 136944
rect 674170 136794 674176 136858
rect 674240 136856 674246 136858
rect 674240 136796 674784 136856
rect 674240 136794 674246 136796
rect 140802 135968 140862 136308
rect 144111 135968 144177 135971
rect 140802 135966 144177 135968
rect 140802 135910 144116 135966
rect 144172 135910 144177 135966
rect 140802 135908 144177 135910
rect 144111 135905 144177 135908
rect 674754 135527 674814 136012
rect 674703 135522 674814 135527
rect 674703 135466 674708 135522
rect 674764 135466 674814 135522
rect 674703 135464 674814 135466
rect 679695 135524 679761 135527
rect 679695 135522 679806 135524
rect 679695 135466 679700 135522
rect 679756 135466 679806 135522
rect 674703 135461 674769 135464
rect 679695 135461 679806 135466
rect 679746 135346 679806 135461
rect 144111 135080 144177 135083
rect 140832 135078 144177 135080
rect 140832 135022 144116 135078
rect 144172 135022 144177 135078
rect 140832 135020 144177 135022
rect 144111 135017 144177 135020
rect 673978 135018 673984 135082
rect 674048 135080 674054 135082
rect 674048 135020 674814 135080
rect 674048 135018 674054 135020
rect 674415 134562 674481 134565
rect 674754 134562 674814 135020
rect 674415 134560 674814 134562
rect 674415 134504 674420 134560
rect 674476 134532 674814 134560
rect 674476 134504 674784 134532
rect 674415 134502 674784 134504
rect 674415 134499 674481 134502
rect 144207 133896 144273 133899
rect 140832 133894 144273 133896
rect 140832 133838 144212 133894
rect 144268 133838 144273 133894
rect 140832 133836 144273 133838
rect 144207 133833 144273 133836
rect 675330 133455 675390 133718
rect 675279 133450 675390 133455
rect 675279 133394 675284 133450
rect 675340 133394 675390 133450
rect 675279 133392 675390 133394
rect 675279 133389 675345 133392
rect 144015 132712 144081 132715
rect 140832 132710 144081 132712
rect 140832 132654 144020 132710
rect 144076 132654 144081 132710
rect 140832 132652 144081 132654
rect 144015 132649 144081 132652
rect 674554 132502 674560 132566
rect 674624 132564 674630 132566
rect 674754 132564 674814 132904
rect 674624 132504 674814 132564
rect 674624 132502 674630 132504
rect 675138 131827 675198 132090
rect 675138 131822 675249 131827
rect 675138 131766 675188 131822
rect 675244 131766 675249 131822
rect 675138 131764 675249 131766
rect 675183 131761 675249 131764
rect 140802 130936 140862 131424
rect 674127 131232 674193 131235
rect 674127 131230 674784 131232
rect 674127 131174 674132 131230
rect 674188 131174 674784 131230
rect 674127 131172 674784 131174
rect 674127 131169 674193 131172
rect 144111 130936 144177 130939
rect 140802 130934 144177 130936
rect 140802 130878 144116 130934
rect 144172 130878 144177 130934
rect 140802 130876 144177 130878
rect 144111 130873 144177 130876
rect 674362 130578 674368 130642
rect 674432 130640 674438 130642
rect 674432 130580 674784 130640
rect 674432 130578 674438 130580
rect 144207 130196 144273 130199
rect 140832 130194 144273 130196
rect 140832 130138 144212 130194
rect 144268 130138 144273 130194
rect 140832 130136 144273 130138
rect 144207 130133 144273 130136
rect 674170 129690 674176 129754
rect 674240 129752 674246 129754
rect 674240 129692 674784 129752
rect 674240 129690 674246 129692
rect 140802 128568 140862 129118
rect 675138 128719 675198 128982
rect 675087 128714 675198 128719
rect 675087 128658 675092 128714
rect 675148 128658 675198 128714
rect 675087 128656 675198 128658
rect 675087 128653 675153 128656
rect 144111 128568 144177 128571
rect 140802 128566 144177 128568
rect 140802 128510 144116 128566
rect 144172 128510 144177 128566
rect 140802 128508 144177 128510
rect 144111 128505 144177 128508
rect 674415 128124 674481 128127
rect 674415 128122 674784 128124
rect 674415 128066 674420 128122
rect 674476 128066 674784 128122
rect 674415 128064 674784 128066
rect 674415 128061 674481 128064
rect 140802 127384 140862 127872
rect 144207 127384 144273 127387
rect 140802 127382 144273 127384
rect 140802 127326 144212 127382
rect 144268 127326 144273 127382
rect 140802 127324 144273 127326
rect 144207 127321 144273 127324
rect 674319 127384 674385 127387
rect 674319 127382 674784 127384
rect 674319 127326 674324 127382
rect 674380 127326 674784 127382
rect 674319 127324 674784 127326
rect 674319 127321 674385 127324
rect 200751 126792 200817 126795
rect 200943 126792 201009 126795
rect 200751 126790 201009 126792
rect 200751 126734 200756 126790
rect 200812 126734 200948 126790
rect 201004 126734 201009 126790
rect 200751 126732 201009 126734
rect 200751 126729 200817 126732
rect 200943 126729 201009 126732
rect 673359 126792 673425 126795
rect 675130 126792 675136 126794
rect 673359 126790 675136 126792
rect 673359 126734 673364 126790
rect 673420 126734 675136 126790
rect 673359 126732 675136 126734
rect 673359 126729 673425 126732
rect 675130 126730 675136 126732
rect 675200 126730 675206 126794
rect 144015 126644 144081 126647
rect 140832 126642 144081 126644
rect 140832 126586 144020 126642
rect 144076 126586 144081 126642
rect 140832 126584 144081 126586
rect 144015 126581 144081 126584
rect 674223 126496 674289 126499
rect 674223 126494 674784 126496
rect 674223 126438 674228 126494
rect 674284 126438 674784 126494
rect 674223 126436 674784 126438
rect 674223 126433 674289 126436
rect 674031 125904 674097 125907
rect 674031 125902 674784 125904
rect 674031 125846 674036 125902
rect 674092 125846 674784 125902
rect 674031 125844 674784 125846
rect 674031 125841 674097 125844
rect 144207 125460 144273 125463
rect 140832 125458 144273 125460
rect 140832 125402 144212 125458
rect 144268 125402 144273 125458
rect 140832 125400 144273 125402
rect 144207 125397 144273 125400
rect 31738 125250 31744 125314
rect 31808 125312 31814 125314
rect 31808 125252 36222 125312
rect 31808 125250 31814 125252
rect 36162 124986 36222 125252
rect 674946 124871 675006 124986
rect 674946 124866 675057 124871
rect 674946 124810 674996 124866
rect 675052 124810 675057 124866
rect 674946 124808 675057 124810
rect 674991 124805 675057 124808
rect 144111 124276 144177 124279
rect 140832 124274 144177 124276
rect 140832 124218 144116 124274
rect 144172 124218 144177 124274
rect 140832 124216 144177 124218
rect 144111 124213 144177 124216
rect 674946 123983 675006 124246
rect 674895 123978 675006 123983
rect 674895 123922 674900 123978
rect 674956 123922 675006 123978
rect 674895 123920 675006 123922
rect 674895 123917 674961 123920
rect 674511 123240 674577 123243
rect 674754 123240 674814 123358
rect 674511 123238 674814 123240
rect 674511 123182 674516 123238
rect 674572 123182 674814 123238
rect 674511 123180 674814 123182
rect 674511 123177 674577 123180
rect 140802 122500 140862 122988
rect 147471 122500 147537 122503
rect 140802 122498 147537 122500
rect 140802 122442 147476 122498
rect 147532 122442 147537 122498
rect 140802 122440 147537 122442
rect 147471 122437 147537 122440
rect 674754 122207 674814 122544
rect 674754 122202 674865 122207
rect 674754 122146 674804 122202
rect 674860 122146 674865 122202
rect 674754 122144 674865 122146
rect 674799 122141 674865 122144
rect 144207 121908 144273 121911
rect 140832 121906 144273 121908
rect 140832 121850 144212 121906
rect 144268 121850 144273 121906
rect 140832 121848 144273 121850
rect 144207 121845 144273 121848
rect 642063 121760 642129 121763
rect 634464 121758 642129 121760
rect 634464 121702 642068 121758
rect 642124 121702 642129 121758
rect 634464 121700 642129 121702
rect 642063 121697 642129 121700
rect 674607 121612 674673 121615
rect 674754 121612 674814 121730
rect 674607 121610 674814 121612
rect 674607 121554 674612 121610
rect 674668 121554 674814 121610
rect 674607 121552 674814 121554
rect 674607 121549 674673 121552
rect 674703 121316 674769 121319
rect 674703 121314 674814 121316
rect 674703 121258 674708 121314
rect 674764 121258 674814 121314
rect 674703 121253 674814 121258
rect 634434 121168 634494 121212
rect 642159 121168 642225 121171
rect 634434 121166 642225 121168
rect 634434 121110 642164 121166
rect 642220 121110 642225 121166
rect 634434 121108 642225 121110
rect 642159 121105 642225 121108
rect 674754 121064 674814 121253
rect 641391 120724 641457 120727
rect 634464 120722 641457 120724
rect 140802 120132 140862 120686
rect 634464 120666 641396 120722
rect 641452 120666 641457 120722
rect 634464 120664 641457 120666
rect 641391 120661 641457 120664
rect 144111 120132 144177 120135
rect 640719 120132 640785 120135
rect 140802 120130 144177 120132
rect 140802 120074 144116 120130
rect 144172 120074 144177 120130
rect 140802 120072 144177 120074
rect 634464 120130 640785 120132
rect 634464 120074 640724 120130
rect 640780 120074 640785 120130
rect 634464 120072 640785 120074
rect 144111 120069 144177 120072
rect 640719 120069 640785 120072
rect 140802 118948 140862 119436
rect 144015 118948 144081 118951
rect 140802 118946 144081 118948
rect 140802 118890 144020 118946
rect 144076 118890 144081 118946
rect 140802 118888 144081 118890
rect 144015 118885 144081 118888
rect 144207 118208 144273 118211
rect 140832 118206 144273 118208
rect 140832 118150 144212 118206
rect 144268 118150 144273 118206
rect 140832 118148 144273 118150
rect 144207 118145 144273 118148
rect 144111 117024 144177 117027
rect 140832 117022 144177 117024
rect 140832 116966 144116 117022
rect 144172 116966 144177 117022
rect 140832 116964 144177 116966
rect 144111 116961 144177 116964
rect 140802 115544 140862 115736
rect 144207 115544 144273 115547
rect 140802 115542 144273 115544
rect 140802 115486 144212 115542
rect 144268 115486 144273 115542
rect 140802 115484 144273 115486
rect 144207 115481 144273 115484
rect 140802 114212 140862 114700
rect 144111 114212 144177 114215
rect 140802 114210 144177 114212
rect 140802 114154 144116 114210
rect 144172 114154 144177 114210
rect 140802 114152 144177 114154
rect 144111 114149 144177 114152
rect 144207 113472 144273 113475
rect 140832 113470 144273 113472
rect 140832 113414 144212 113470
rect 144268 113414 144273 113470
rect 140832 113412 144273 113414
rect 144207 113409 144273 113412
rect 665199 112288 665265 112291
rect 665154 112286 665265 112288
rect 140802 111696 140862 112254
rect 665154 112230 665204 112286
rect 665260 112230 665265 112286
rect 665154 112225 665265 112230
rect 665154 112083 665214 112225
rect 144015 111696 144081 111699
rect 140802 111694 144081 111696
rect 140802 111638 144020 111694
rect 144076 111638 144081 111694
rect 140802 111636 144081 111638
rect 144015 111633 144081 111636
rect 665346 111252 665406 111718
rect 668175 111252 668241 111255
rect 665346 111250 668241 111252
rect 665346 111194 668180 111250
rect 668236 111194 668241 111250
rect 665346 111192 668241 111194
rect 668175 111189 668241 111192
rect 140802 110512 140862 111000
rect 665346 110808 665406 110996
rect 674895 110808 674961 110811
rect 675130 110808 675136 110810
rect 665346 110806 675136 110808
rect 665346 110750 674900 110806
rect 674956 110750 675136 110806
rect 665346 110748 675136 110750
rect 674895 110745 674961 110748
rect 675130 110746 675136 110748
rect 675200 110746 675206 110810
rect 144111 110512 144177 110515
rect 140802 110510 144177 110512
rect 140802 110454 144116 110510
rect 144172 110454 144177 110510
rect 140802 110452 144177 110454
rect 144111 110449 144177 110452
rect 675567 110070 675633 110071
rect 675514 110068 675520 110070
rect 675476 110008 675520 110068
rect 675584 110066 675633 110070
rect 675628 110010 675633 110066
rect 675514 110006 675520 110008
rect 675584 110006 675633 110010
rect 675567 110005 675633 110006
rect 140802 109772 140862 109806
rect 144207 109772 144273 109775
rect 140802 109770 144273 109772
rect 140802 109714 144212 109770
rect 144268 109714 144273 109770
rect 140802 109712 144273 109714
rect 144207 109709 144273 109712
rect 147567 108588 147633 108591
rect 140832 108586 147633 108588
rect 140832 108530 147572 108586
rect 147628 108530 147633 108586
rect 140832 108528 147633 108530
rect 147567 108525 147633 108528
rect 674362 108082 674368 108146
rect 674432 108144 674438 108146
rect 675375 108144 675441 108147
rect 674432 108142 675441 108144
rect 674432 108086 675380 108142
rect 675436 108086 675441 108142
rect 674432 108084 675441 108086
rect 674432 108082 674438 108084
rect 675375 108081 675441 108084
rect 140802 106960 140862 107300
rect 144207 106960 144273 106963
rect 140802 106958 144273 106960
rect 140802 106902 144212 106958
rect 144268 106902 144273 106958
rect 140802 106900 144273 106902
rect 144207 106897 144273 106900
rect 140802 105776 140862 106264
rect 144015 105776 144081 105779
rect 140802 105774 144081 105776
rect 140802 105718 144020 105774
rect 144076 105718 144081 105774
rect 140802 105716 144081 105718
rect 144015 105713 144081 105716
rect 144111 105036 144177 105039
rect 140832 105034 144177 105036
rect 140832 104978 144116 105034
rect 144172 104978 144177 105034
rect 140832 104976 144177 104978
rect 144111 104973 144177 104976
rect 144207 103852 144273 103855
rect 140832 103850 144273 103852
rect 140832 103794 144212 103850
rect 144268 103794 144273 103850
rect 140832 103792 144273 103794
rect 144207 103789 144273 103792
rect 674554 103198 674560 103262
rect 674624 103260 674630 103262
rect 675375 103260 675441 103263
rect 674624 103258 675441 103260
rect 674624 103202 675380 103258
rect 675436 103202 675441 103258
rect 674624 103200 675441 103202
rect 674624 103198 674630 103200
rect 675375 103197 675441 103200
rect 140802 102076 140862 102564
rect 144207 102076 144273 102079
rect 140802 102074 144273 102076
rect 140802 102018 144212 102074
rect 144268 102018 144273 102074
rect 140802 102016 144273 102018
rect 144207 102013 144273 102016
rect 674170 101422 674176 101486
rect 674240 101484 674246 101486
rect 675375 101484 675441 101487
rect 674240 101482 675441 101484
rect 674240 101426 675380 101482
rect 675436 101426 675441 101482
rect 674240 101424 675441 101426
rect 674240 101422 674246 101424
rect 675375 101421 675441 101424
rect 140802 100892 140862 101374
rect 147375 100892 147441 100895
rect 140802 100890 147441 100892
rect 140802 100834 147380 100890
rect 147436 100834 147441 100890
rect 140802 100832 147441 100834
rect 147375 100829 147441 100832
rect 144207 100152 144273 100155
rect 140832 100150 144273 100152
rect 140832 100094 144212 100150
rect 144268 100094 144273 100150
rect 140832 100092 144273 100094
rect 144207 100089 144273 100092
rect 140802 98524 140862 99012
rect 147279 98524 147345 98527
rect 140802 98522 147345 98524
rect 140802 98466 147284 98522
rect 147340 98466 147345 98522
rect 140802 98464 147345 98466
rect 147279 98461 147345 98464
rect 140802 97340 140862 97828
rect 144111 97340 144177 97343
rect 140802 97338 144177 97340
rect 140802 97282 144116 97338
rect 144172 97282 144177 97338
rect 140802 97280 144177 97282
rect 144111 97277 144177 97280
rect 144207 96600 144273 96603
rect 140832 96598 144273 96600
rect 140832 96542 144212 96598
rect 144268 96542 144273 96598
rect 140832 96540 144273 96542
rect 144207 96537 144273 96540
rect 144015 95416 144081 95419
rect 140832 95414 144081 95416
rect 140832 95358 144020 95414
rect 144076 95358 144081 95414
rect 140832 95356 144081 95358
rect 144015 95353 144081 95356
rect 140802 93640 140862 94128
rect 144207 93640 144273 93643
rect 140802 93638 144273 93640
rect 140802 93582 144212 93638
rect 144268 93582 144273 93638
rect 140802 93580 144273 93582
rect 144207 93577 144273 93580
rect 198831 93492 198897 93495
rect 198831 93490 204576 93492
rect 198831 93434 198836 93490
rect 198892 93434 204576 93490
rect 198831 93432 204576 93434
rect 198831 93429 198897 93432
rect 198927 93344 198993 93347
rect 198927 93342 204606 93344
rect 198927 93286 198932 93342
rect 198988 93286 204606 93342
rect 198927 93284 204606 93286
rect 198927 93281 198993 93284
rect 204546 92944 204606 93284
rect 140802 92308 140862 92942
rect 198735 92456 198801 92459
rect 198735 92454 204576 92456
rect 198735 92398 198740 92454
rect 198796 92398 204576 92454
rect 198735 92396 204576 92398
rect 198735 92393 198801 92396
rect 143919 92308 143985 92311
rect 140802 92306 143985 92308
rect 140802 92250 143924 92306
rect 143980 92250 143985 92306
rect 140802 92248 143985 92250
rect 143919 92245 143985 92248
rect 144111 91864 144177 91867
rect 140832 91862 144177 91864
rect 140832 91806 144116 91862
rect 144172 91806 144177 91862
rect 140832 91804 144177 91806
rect 144111 91801 144177 91804
rect 198735 91864 198801 91867
rect 198735 91862 204576 91864
rect 198735 91806 198740 91862
rect 198796 91806 204576 91862
rect 198735 91804 204576 91806
rect 198735 91801 198801 91804
rect 199119 91716 199185 91719
rect 199119 91714 204606 91716
rect 199119 91658 199124 91714
rect 199180 91658 204606 91714
rect 199119 91656 204606 91658
rect 199119 91653 199185 91656
rect 204546 91316 204606 91656
rect 198831 91124 198897 91127
rect 198831 91122 204606 91124
rect 198831 91066 198836 91122
rect 198892 91066 204606 91122
rect 198831 91064 204606 91066
rect 198831 91061 198897 91064
rect 204546 90798 204606 91064
rect 144207 90680 144273 90683
rect 140832 90678 144273 90680
rect 140832 90622 144212 90678
rect 144268 90622 144273 90678
rect 140832 90620 144273 90622
rect 144207 90617 144273 90620
rect 199023 90236 199089 90239
rect 199023 90234 204576 90236
rect 199023 90178 199028 90234
rect 199084 90178 204576 90234
rect 199023 90176 204576 90178
rect 199023 90173 199089 90176
rect 198927 90088 198993 90091
rect 198927 90086 204606 90088
rect 198927 90030 198932 90086
rect 198988 90030 204606 90086
rect 198927 90028 204606 90030
rect 198927 90025 198993 90028
rect 204546 89614 204606 90028
rect 140802 89348 140862 89392
rect 144207 89348 144273 89351
rect 140802 89346 144273 89348
rect 140802 89290 144212 89346
rect 144268 89290 144273 89346
rect 140802 89288 144273 89290
rect 144207 89285 144273 89288
rect 198735 89052 198801 89055
rect 204546 89052 204606 89170
rect 198735 89050 204606 89052
rect 198735 88994 198740 89050
rect 198796 88994 204606 89050
rect 198735 88992 204606 88994
rect 198735 88989 198801 88992
rect 198927 88608 198993 88611
rect 198927 88606 204576 88608
rect 198927 88550 198932 88606
rect 198988 88550 204576 88606
rect 198927 88548 204576 88550
rect 198927 88545 198993 88548
rect 199215 88460 199281 88463
rect 199215 88458 204606 88460
rect 199215 88402 199220 88458
rect 199276 88402 204606 88458
rect 199215 88400 204606 88402
rect 199215 88397 199281 88400
rect 144111 88164 144177 88167
rect 140832 88162 144177 88164
rect 140832 88106 144116 88162
rect 144172 88106 144177 88162
rect 140832 88104 144177 88106
rect 144111 88101 144177 88104
rect 204546 87986 204606 88400
rect 198831 87868 198897 87871
rect 198831 87866 204798 87868
rect 198831 87810 198836 87866
rect 198892 87810 204798 87866
rect 198831 87808 204798 87810
rect 198831 87805 198897 87808
rect 204738 87542 204798 87808
rect 144207 86980 144273 86983
rect 140832 86978 144273 86980
rect 140832 86922 144212 86978
rect 144268 86922 144273 86978
rect 140832 86920 144273 86922
rect 144207 86917 144273 86920
rect 199023 86980 199089 86983
rect 652623 86980 652689 86983
rect 199023 86978 204576 86980
rect 199023 86922 199028 86978
rect 199084 86922 204576 86978
rect 199023 86920 204576 86922
rect 652623 86978 656736 86980
rect 652623 86922 652628 86978
rect 652684 86922 656736 86978
rect 652623 86920 656736 86922
rect 199023 86917 199089 86920
rect 652623 86917 652689 86920
rect 204346 86622 204352 86686
rect 204416 86684 204422 86686
rect 204879 86684 204945 86687
rect 204416 86682 204945 86684
rect 204416 86626 204884 86682
rect 204940 86626 204945 86682
rect 204416 86624 204945 86626
rect 204416 86622 204422 86624
rect 204879 86621 204945 86624
rect 198831 86240 198897 86243
rect 204738 86240 204798 86358
rect 198831 86238 204798 86240
rect 198831 86182 198836 86238
rect 198892 86182 204798 86238
rect 198831 86180 204798 86182
rect 653583 86240 653649 86243
rect 653583 86238 656736 86240
rect 653583 86182 653588 86238
rect 653644 86182 656736 86238
rect 653583 86180 656736 86182
rect 198831 86177 198897 86180
rect 653583 86177 653649 86180
rect 198735 86092 198801 86095
rect 198735 86090 204798 86092
rect 198735 86034 198740 86090
rect 198796 86034 204798 86090
rect 198735 86032 204798 86034
rect 198735 86029 198801 86032
rect 204738 85914 204798 86032
rect 140802 85204 140862 85692
rect 663426 85651 663486 86210
rect 663375 85646 663486 85651
rect 663375 85590 663380 85646
rect 663436 85590 663486 85646
rect 663375 85588 663486 85590
rect 663375 85585 663441 85588
rect 198927 85352 198993 85355
rect 653487 85352 653553 85355
rect 198927 85350 204576 85352
rect 198927 85294 198932 85350
rect 198988 85294 204576 85350
rect 198927 85292 204576 85294
rect 653487 85350 656736 85352
rect 653487 85294 653492 85350
rect 653548 85294 656736 85350
rect 653487 85292 656736 85294
rect 198927 85289 198993 85292
rect 653487 85289 653553 85292
rect 144111 85204 144177 85207
rect 140802 85202 144177 85204
rect 140802 85146 144116 85202
rect 144172 85146 144177 85202
rect 140802 85144 144177 85146
rect 144111 85141 144177 85144
rect 199119 85056 199185 85059
rect 199119 85054 204606 85056
rect 199119 84998 199124 85054
rect 199180 84998 204606 85054
rect 199119 84996 204606 84998
rect 199119 84993 199185 84996
rect 204546 84730 204606 84996
rect 663618 84763 663678 85322
rect 663567 84758 663678 84763
rect 663567 84702 663572 84758
rect 663628 84702 663678 84758
rect 663567 84700 663678 84702
rect 663567 84697 663633 84700
rect 199023 84612 199089 84615
rect 199023 84610 204798 84612
rect 199023 84554 199028 84610
rect 199084 84554 204798 84610
rect 199023 84552 204798 84554
rect 199023 84549 199089 84552
rect 140802 83872 140862 84508
rect 204738 84286 204798 84552
rect 653679 84316 653745 84319
rect 653679 84314 656736 84316
rect 653679 84258 653684 84314
rect 653740 84258 656736 84314
rect 653679 84256 656736 84258
rect 653679 84253 653745 84256
rect 663234 84023 663294 84582
rect 663234 84018 663345 84023
rect 663234 83962 663284 84018
rect 663340 83962 663345 84018
rect 663234 83960 663345 83962
rect 663279 83957 663345 83960
rect 146895 83872 146961 83875
rect 140802 83870 146961 83872
rect 140802 83814 146900 83870
rect 146956 83814 146961 83870
rect 140802 83812 146961 83814
rect 146895 83809 146961 83812
rect 199215 83724 199281 83727
rect 199215 83722 204576 83724
rect 199215 83666 199220 83722
rect 199276 83666 204576 83722
rect 199215 83664 204576 83666
rect 199215 83661 199281 83664
rect 144111 83428 144177 83431
rect 140832 83426 144177 83428
rect 140832 83370 144116 83426
rect 144172 83370 144177 83426
rect 140832 83368 144177 83370
rect 144111 83365 144177 83368
rect 653583 83428 653649 83431
rect 653583 83426 656736 83428
rect 653583 83370 653588 83426
rect 653644 83370 656736 83426
rect 653583 83368 656736 83370
rect 653583 83365 653649 83368
rect 198735 83280 198801 83283
rect 198735 83278 204606 83280
rect 198735 83222 198740 83278
rect 198796 83222 204606 83278
rect 198735 83220 204606 83222
rect 198735 83217 198801 83220
rect 204546 83102 204606 83220
rect 200751 82984 200817 82987
rect 200751 82982 204798 82984
rect 200751 82926 200756 82982
rect 200812 82926 204798 82982
rect 200751 82924 204798 82926
rect 200751 82921 200817 82924
rect 204738 82658 204798 82924
rect 663426 82839 663486 83398
rect 663426 82834 663537 82839
rect 663426 82778 663476 82834
rect 663532 82778 663537 82834
rect 663426 82776 663537 82778
rect 663471 82773 663537 82776
rect 653679 82688 653745 82691
rect 653679 82686 656736 82688
rect 653679 82630 653684 82686
rect 653740 82630 656736 82686
rect 653679 82628 656736 82630
rect 653679 82625 653745 82628
rect 146991 82244 147057 82247
rect 140832 82242 147057 82244
rect 140832 82186 146996 82242
rect 147052 82186 147057 82242
rect 140832 82184 147057 82186
rect 146991 82181 147057 82184
rect 663234 82099 663294 82658
rect 199503 82096 199569 82099
rect 199503 82094 204576 82096
rect 199503 82038 199508 82094
rect 199564 82038 204576 82094
rect 199503 82036 204576 82038
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 199503 82033 199569 82036
rect 663279 82033 663345 82036
rect 198831 81800 198897 81803
rect 198831 81798 204606 81800
rect 198831 81742 198836 81798
rect 198892 81742 204606 81798
rect 198831 81740 204606 81742
rect 198831 81737 198897 81740
rect 204546 81474 204606 81740
rect 198927 81356 198993 81359
rect 198927 81354 204606 81356
rect 198927 81298 198932 81354
rect 198988 81298 204606 81354
rect 198927 81296 204606 81298
rect 198927 81293 198993 81296
rect 146895 81060 146961 81063
rect 140832 81058 146961 81060
rect 140832 81002 146900 81058
rect 146956 81002 146961 81058
rect 140832 81000 146961 81002
rect 146895 80997 146961 81000
rect 204546 80956 204606 81296
rect 662415 81208 662481 81211
rect 663042 81208 663102 81770
rect 662415 81206 663102 81208
rect 662415 81150 662420 81206
rect 662476 81150 663102 81206
rect 662415 81148 663102 81150
rect 662415 81145 662481 81148
rect 198735 80468 198801 80471
rect 198735 80466 204576 80468
rect 198735 80410 198740 80466
rect 198796 80410 204576 80466
rect 198735 80408 204576 80410
rect 198735 80405 198801 80408
rect 198735 79876 198801 79879
rect 198735 79874 204576 79876
rect 198735 79818 198740 79874
rect 198796 79818 204576 79874
rect 198735 79816 204576 79818
rect 198735 79813 198801 79816
rect 144111 79728 144177 79731
rect 140832 79726 144177 79728
rect 140832 79670 144116 79726
rect 144172 79670 144177 79726
rect 140832 79668 144177 79670
rect 144111 79665 144177 79668
rect 198831 79728 198897 79731
rect 198831 79726 204606 79728
rect 198831 79670 198836 79726
rect 198892 79670 204606 79726
rect 198831 79668 204606 79670
rect 198831 79665 198897 79668
rect 204546 79328 204606 79668
rect 198927 78840 198993 78843
rect 198927 78838 204576 78840
rect 198927 78782 198932 78838
rect 198988 78782 204576 78838
rect 198927 78780 204576 78782
rect 198927 78777 198993 78780
rect 144207 78544 144273 78547
rect 140832 78542 144273 78544
rect 140832 78486 144212 78542
rect 144268 78486 144273 78542
rect 140832 78484 144273 78486
rect 144207 78481 144273 78484
rect 199023 78248 199089 78251
rect 199023 78246 204576 78248
rect 199023 78190 199028 78246
rect 199084 78190 204576 78246
rect 199023 78188 204576 78190
rect 199023 78185 199089 78188
rect 198735 77656 198801 77659
rect 204546 77656 204606 77700
rect 198735 77654 204606 77656
rect 198735 77598 198740 77654
rect 198796 77598 204606 77654
rect 198735 77596 204606 77598
rect 198735 77593 198801 77596
rect 144207 77360 144273 77363
rect 140832 77358 144273 77360
rect 140832 77302 144212 77358
rect 144268 77302 144273 77358
rect 140832 77300 144273 77302
rect 144207 77297 144273 77300
rect 198735 77212 198801 77215
rect 198735 77210 204576 77212
rect 198735 77154 198740 77210
rect 198796 77154 204576 77210
rect 198735 77152 204576 77154
rect 198735 77149 198801 77152
rect 198927 76620 198993 76623
rect 198927 76618 204576 76620
rect 198927 76562 198932 76618
rect 198988 76562 204576 76618
rect 198927 76560 204576 76562
rect 198927 76557 198993 76560
rect 198831 76472 198897 76475
rect 198831 76470 204606 76472
rect 198831 76414 198836 76470
rect 198892 76414 204606 76470
rect 198831 76412 204606 76414
rect 198831 76409 198897 76412
rect 140802 75880 140862 76214
rect 204546 76072 204606 76412
rect 144207 75880 144273 75883
rect 140802 75878 144273 75880
rect 140802 75822 144212 75878
rect 144268 75822 144273 75878
rect 140802 75820 144273 75822
rect 144207 75817 144273 75820
rect 199023 75584 199089 75587
rect 642159 75584 642225 75587
rect 199023 75582 204576 75584
rect 199023 75526 199028 75582
rect 199084 75526 204576 75582
rect 199023 75524 204576 75526
rect 634464 75582 642225 75584
rect 634464 75526 642164 75582
rect 642220 75526 642225 75582
rect 634464 75524 642225 75526
rect 199023 75521 199089 75524
rect 642159 75521 642225 75524
rect 146895 74992 146961 74995
rect 140832 74990 146961 74992
rect 140832 74934 146900 74990
rect 146956 74934 146961 74990
rect 140832 74932 146961 74934
rect 146895 74929 146961 74932
rect 199119 74992 199185 74995
rect 199119 74990 204576 74992
rect 199119 74934 199124 74990
rect 199180 74934 204576 74990
rect 199119 74932 204576 74934
rect 199119 74929 199185 74932
rect 198735 74548 198801 74551
rect 198735 74546 204606 74548
rect 198735 74490 198740 74546
rect 198796 74490 204606 74546
rect 198735 74488 204606 74490
rect 198735 74485 198801 74488
rect 204546 74444 204606 74488
rect 198927 73956 198993 73959
rect 198927 73954 204576 73956
rect 198927 73898 198932 73954
rect 198988 73898 204576 73954
rect 198927 73896 204576 73898
rect 198927 73893 198993 73896
rect 143919 73808 143985 73811
rect 140832 73806 143985 73808
rect 140832 73750 143924 73806
rect 143980 73750 143985 73806
rect 140832 73748 143985 73750
rect 143919 73745 143985 73748
rect 198831 73364 198897 73367
rect 198831 73362 204576 73364
rect 198831 73306 198836 73362
rect 198892 73306 204576 73362
rect 198831 73304 204576 73306
rect 198831 73301 198897 73304
rect 199023 73216 199089 73219
rect 199023 73214 204606 73216
rect 199023 73158 199028 73214
rect 199084 73158 204606 73214
rect 199023 73156 204606 73158
rect 199023 73153 199089 73156
rect 204546 72816 204606 73156
rect 140802 72180 140862 72520
rect 199119 72328 199185 72331
rect 199119 72326 204576 72328
rect 199119 72270 199124 72326
rect 199180 72270 204576 72326
rect 199119 72268 204576 72270
rect 199119 72265 199185 72268
rect 143919 72180 143985 72183
rect 140802 72178 143985 72180
rect 140802 72122 143924 72178
rect 143980 72122 143985 72178
rect 140802 72120 143985 72122
rect 143919 72117 143985 72120
rect 198735 71736 198801 71739
rect 198735 71734 204576 71736
rect 198735 71678 198740 71734
rect 198796 71678 204576 71734
rect 198735 71676 204576 71678
rect 198735 71673 198801 71676
rect 200751 71588 200817 71591
rect 200751 71586 204606 71588
rect 200751 71530 200756 71586
rect 200812 71530 204606 71586
rect 200751 71528 204606 71530
rect 200751 71525 200817 71528
rect 146991 71292 147057 71295
rect 140832 71290 147057 71292
rect 140832 71234 146996 71290
rect 147052 71234 147057 71290
rect 140832 71232 147057 71234
rect 146991 71229 147057 71232
rect 204546 71188 204606 71528
rect 199599 70996 199665 70999
rect 199599 70994 204606 70996
rect 199599 70938 199604 70994
rect 199660 70938 204606 70994
rect 199599 70936 204606 70938
rect 199599 70933 199665 70936
rect 204546 70670 204606 70936
rect 146895 70108 146961 70111
rect 140832 70106 146961 70108
rect 140832 70050 146900 70106
rect 146956 70050 146961 70106
rect 140832 70048 146961 70050
rect 146895 70045 146961 70048
rect 198831 70108 198897 70111
rect 198831 70106 204576 70108
rect 198831 70050 198836 70106
rect 198892 70050 204576 70106
rect 198831 70048 204576 70050
rect 198831 70045 198897 70048
rect 198927 69960 198993 69963
rect 198927 69958 204606 69960
rect 198927 69902 198932 69958
rect 198988 69902 204606 69958
rect 198927 69900 204606 69902
rect 198927 69897 198993 69900
rect 204546 69486 204606 69900
rect 140802 68332 140862 68968
rect 198831 68924 198897 68927
rect 204546 68924 204606 69042
rect 198831 68922 204606 68924
rect 198831 68866 198836 68922
rect 198892 68866 204606 68922
rect 198831 68864 204606 68866
rect 198831 68861 198897 68864
rect 199023 68480 199089 68483
rect 199023 68478 204576 68480
rect 199023 68422 199028 68478
rect 199084 68422 204576 68478
rect 199023 68420 204576 68422
rect 199023 68417 199089 68420
rect 143823 68332 143889 68335
rect 140802 68330 143889 68332
rect 140802 68274 143828 68330
rect 143884 68274 143889 68330
rect 140802 68272 143889 68274
rect 143823 68269 143889 68272
rect 198735 68332 198801 68335
rect 198735 68330 204606 68332
rect 198735 68274 198740 68330
rect 198796 68274 204606 68330
rect 198735 68272 204606 68274
rect 198735 68269 198801 68272
rect 204546 67858 204606 68272
rect 140802 67148 140862 67782
rect 198927 67740 198993 67743
rect 198927 67738 204798 67740
rect 198927 67682 198932 67738
rect 198988 67682 204798 67738
rect 198927 67680 204798 67682
rect 198927 67677 198993 67680
rect 204738 67414 204798 67680
rect 143919 67148 143985 67151
rect 140802 67146 143985 67148
rect 140802 67090 143924 67146
rect 143980 67090 143985 67146
rect 140802 67088 143985 67090
rect 143919 67085 143985 67088
rect 143919 66852 143985 66855
rect 140610 66850 143985 66852
rect 140610 66794 143924 66850
rect 143980 66794 143985 66850
rect 140610 66792 143985 66794
rect 140610 66600 140670 66792
rect 143919 66789 143985 66792
rect 199119 66852 199185 66855
rect 199119 66850 204576 66852
rect 199119 66794 199124 66850
rect 199180 66794 204576 66850
rect 199119 66792 204576 66794
rect 199119 66789 199185 66792
rect 198927 66112 198993 66115
rect 204738 66112 204798 66230
rect 198927 66110 204798 66112
rect 198927 66054 198932 66110
rect 198988 66054 204798 66110
rect 198927 66052 204798 66054
rect 198927 66049 198993 66052
rect 198735 65964 198801 65967
rect 198735 65962 204798 65964
rect 198735 65906 198740 65962
rect 198796 65906 204798 65962
rect 198735 65904 204798 65906
rect 198735 65901 198801 65904
rect 204738 65786 204798 65904
rect 140802 64780 140862 65334
rect 198831 65224 198897 65227
rect 198831 65222 204576 65224
rect 198831 65166 198836 65222
rect 198892 65166 204576 65222
rect 198831 65164 204576 65166
rect 198831 65161 198897 65164
rect 199023 64928 199089 64931
rect 199023 64926 204606 64928
rect 199023 64870 199028 64926
rect 199084 64870 204606 64926
rect 199023 64868 204606 64870
rect 199023 64865 199089 64868
rect 143919 64780 143985 64783
rect 140802 64778 143985 64780
rect 140802 64722 143924 64778
rect 143980 64722 143985 64778
rect 140802 64720 143985 64722
rect 143919 64717 143985 64720
rect 204546 64602 204606 64868
rect 199119 64484 199185 64487
rect 199119 64482 204798 64484
rect 199119 64426 199124 64482
rect 199180 64426 204798 64482
rect 199119 64424 204798 64426
rect 199119 64421 199185 64424
rect 146895 64188 146961 64191
rect 140832 64186 146961 64188
rect 140832 64130 146900 64186
rect 146956 64130 146961 64186
rect 204738 64158 204798 64424
rect 140832 64128 146961 64130
rect 146895 64125 146961 64128
rect 199215 63596 199281 63599
rect 199215 63594 204576 63596
rect 199215 63538 199220 63594
rect 199276 63538 204576 63594
rect 199215 63536 204576 63538
rect 199215 63533 199281 63536
rect 198735 63152 198801 63155
rect 198735 63150 204606 63152
rect 198735 63094 198740 63150
rect 198796 63094 204606 63150
rect 198735 63092 204606 63094
rect 198735 63089 198801 63092
rect 204546 62974 204606 63092
rect 198831 62856 198897 62859
rect 198831 62854 204798 62856
rect 140802 62264 140862 62826
rect 198831 62798 198836 62854
rect 198892 62798 204798 62854
rect 198831 62796 204798 62798
rect 198831 62793 198897 62796
rect 204738 62530 204798 62796
rect 146991 62264 147057 62267
rect 140802 62262 147057 62264
rect 140802 62206 146996 62262
rect 147052 62206 147057 62262
rect 140802 62204 147057 62206
rect 146991 62201 147057 62204
rect 204015 62264 204081 62267
rect 204154 62264 204160 62266
rect 204015 62262 204160 62264
rect 204015 62206 204020 62262
rect 204076 62206 204160 62262
rect 204015 62204 204160 62206
rect 204015 62201 204081 62204
rect 204154 62202 204160 62204
rect 204224 62202 204230 62266
rect 198927 61968 198993 61971
rect 198927 61966 204576 61968
rect 198927 61910 198932 61966
rect 198988 61910 204576 61966
rect 198927 61908 204576 61910
rect 198927 61905 198993 61908
rect 140802 61228 140862 61790
rect 199023 61672 199089 61675
rect 199023 61670 204606 61672
rect 199023 61614 199028 61670
rect 199084 61614 204606 61670
rect 199023 61612 204606 61614
rect 199023 61609 199089 61612
rect 204546 61346 204606 61612
rect 641007 61376 641073 61379
rect 634434 61374 641073 61376
rect 634434 61318 641012 61374
rect 641068 61318 641073 61374
rect 634434 61316 641073 61318
rect 146895 61228 146961 61231
rect 140802 61226 146961 61228
rect 140802 61170 146900 61226
rect 146956 61170 146961 61226
rect 140802 61168 146961 61170
rect 146895 61165 146961 61168
rect 199119 61228 199185 61231
rect 199119 61226 204606 61228
rect 199119 61170 199124 61226
rect 199180 61170 204606 61226
rect 199119 61168 204606 61170
rect 199119 61165 199185 61168
rect 204546 60828 204606 61168
rect 634434 60828 634494 61316
rect 641007 61313 641073 61316
rect 198735 60340 198801 60343
rect 640143 60340 640209 60343
rect 198735 60338 204576 60340
rect 198735 60282 198740 60338
rect 198796 60282 204576 60338
rect 198735 60280 204576 60282
rect 634464 60338 640209 60340
rect 634464 60282 640148 60338
rect 640204 60282 640209 60338
rect 634464 60280 640209 60282
rect 198735 60277 198801 60280
rect 640143 60277 640209 60280
rect 198831 59748 198897 59751
rect 641583 59748 641649 59751
rect 198831 59746 204576 59748
rect 198831 59690 198836 59746
rect 198892 59690 204576 59746
rect 198831 59688 204576 59690
rect 634464 59746 641649 59748
rect 634464 59690 641588 59746
rect 641644 59690 641649 59746
rect 634464 59688 641649 59690
rect 198831 59685 198897 59688
rect 641583 59685 641649 59688
rect 198927 59600 198993 59603
rect 641391 59600 641457 59603
rect 198927 59598 204606 59600
rect 198927 59542 198932 59598
rect 198988 59542 204606 59598
rect 198927 59540 204606 59542
rect 198927 59537 198993 59540
rect 204546 59200 204606 59540
rect 634434 59598 641457 59600
rect 634434 59542 641396 59598
rect 641452 59542 641457 59598
rect 634434 59540 641457 59542
rect 634434 59200 634494 59540
rect 641391 59537 641457 59540
rect 204687 58862 204753 58863
rect 204687 58858 204736 58862
rect 204800 58860 204806 58862
rect 204687 58802 204692 58858
rect 204687 58798 204736 58802
rect 204800 58800 204844 58860
rect 204800 58798 204806 58800
rect 204687 58797 204753 58798
rect 640815 58712 640881 58715
rect 634464 58710 640881 58712
rect 204546 58419 204606 58682
rect 634464 58654 640820 58710
rect 640876 58654 640881 58710
rect 634464 58652 640881 58654
rect 640815 58649 640881 58652
rect 204546 58414 204657 58419
rect 204546 58358 204596 58414
rect 204652 58358 204657 58414
rect 204546 58356 204657 58358
rect 204591 58353 204657 58356
rect 204399 58120 204465 58123
rect 641199 58120 641265 58123
rect 204399 58118 204576 58120
rect 204399 58062 204404 58118
rect 204460 58062 204576 58118
rect 204399 58060 204576 58062
rect 634464 58118 641265 58120
rect 634464 58062 641204 58118
rect 641260 58062 641265 58118
rect 634464 58060 641265 58062
rect 204399 58057 204465 58060
rect 641199 58057 641265 58060
rect 204546 57235 204606 57572
rect 634434 57528 634494 57572
rect 640911 57528 640977 57531
rect 634434 57526 640977 57528
rect 634434 57470 640916 57526
rect 640972 57470 640977 57526
rect 634434 57468 640977 57470
rect 640911 57465 640977 57468
rect 204495 57230 204606 57235
rect 204495 57174 204500 57230
rect 204556 57174 204606 57230
rect 204495 57172 204606 57174
rect 204495 57169 204561 57172
rect 641295 57084 641361 57087
rect 634464 57082 641361 57084
rect 204930 56790 204990 57054
rect 634464 57026 641300 57082
rect 641356 57026 641361 57082
rect 634464 57024 641361 57026
rect 641295 57021 641361 57024
rect 204922 56726 204928 56790
rect 204992 56726 204998 56790
rect 641103 56492 641169 56495
rect 634464 56490 641169 56492
rect 204738 56199 204798 56462
rect 634464 56434 641108 56490
rect 641164 56434 641169 56490
rect 634464 56432 641169 56434
rect 641103 56429 641169 56432
rect 641679 56344 641745 56347
rect 204687 56194 204798 56199
rect 204687 56138 204692 56194
rect 204748 56138 204798 56194
rect 204687 56136 204798 56138
rect 634434 56342 641745 56344
rect 634434 56286 641684 56342
rect 641740 56286 641745 56342
rect 634434 56284 641745 56286
rect 204687 56133 204753 56136
rect 634434 55944 634494 56284
rect 641679 56281 641745 56284
rect 201327 55604 201393 55607
rect 204546 55604 204606 55944
rect 201327 55602 204606 55604
rect 201327 55546 201332 55602
rect 201388 55546 204606 55602
rect 201327 55544 204606 55546
rect 201327 55541 201393 55544
rect 640719 55456 640785 55459
rect 634464 55454 640785 55456
rect 204738 55163 204798 55426
rect 634464 55398 640724 55454
rect 640780 55398 640785 55454
rect 634464 55396 640785 55398
rect 640719 55393 640785 55396
rect 204738 55158 204849 55163
rect 204738 55102 204788 55158
rect 204844 55102 204849 55158
rect 204738 55100 204849 55102
rect 204783 55097 204849 55100
rect 641487 54864 641553 54867
rect 634464 54862 641553 54864
rect 204930 54719 204990 54834
rect 634464 54806 641492 54862
rect 641548 54806 641553 54862
rect 634464 54804 641553 54806
rect 641487 54801 641553 54804
rect 143919 54716 143985 54719
rect 144207 54716 144273 54719
rect 143919 54714 144273 54716
rect 143919 54658 143924 54714
rect 143980 54658 144212 54714
rect 144268 54658 144273 54714
rect 143919 54656 144273 54658
rect 204930 54714 205041 54719
rect 204930 54658 204980 54714
rect 205036 54658 205041 54714
rect 204930 54656 205041 54658
rect 143919 54653 143985 54656
rect 144207 54653 144273 54656
rect 204975 54653 205041 54656
rect 206074 54654 206080 54718
rect 206144 54716 206150 54718
rect 206144 54656 215022 54716
rect 206144 54654 206150 54656
rect 204879 54568 204945 54571
rect 204879 54566 210558 54568
rect 204879 54510 204884 54566
rect 204940 54510 210558 54566
rect 204879 54508 210558 54510
rect 204879 54505 204945 54508
rect 206266 54358 206272 54422
rect 206336 54420 206342 54422
rect 206336 54360 210414 54420
rect 206336 54358 206342 54360
rect 210354 54275 210414 54360
rect 207418 54210 207424 54274
rect 207488 54272 207494 54274
rect 207488 54212 208830 54272
rect 207488 54210 207494 54212
rect 207994 54062 208000 54126
rect 208064 54124 208070 54126
rect 208527 54124 208593 54127
rect 208064 54122 208593 54124
rect 208064 54066 208532 54122
rect 208588 54066 208593 54122
rect 208064 54064 208593 54066
rect 208770 54124 208830 54212
rect 210351 54270 210417 54275
rect 210351 54214 210356 54270
rect 210412 54214 210417 54270
rect 210351 54209 210417 54214
rect 210498 54272 210558 54508
rect 214962 54275 215022 54656
rect 635343 54420 635409 54423
rect 627138 54418 635409 54420
rect 627138 54362 635348 54418
rect 635404 54362 635409 54418
rect 627138 54360 635409 54362
rect 627138 54275 627198 54360
rect 635343 54357 635409 54360
rect 214767 54272 214833 54275
rect 210498 54270 214833 54272
rect 210498 54214 214772 54270
rect 214828 54214 214833 54270
rect 210498 54212 214833 54214
rect 214767 54209 214833 54212
rect 214959 54270 215025 54275
rect 214959 54214 214964 54270
rect 215020 54214 215025 54270
rect 214959 54209 215025 54214
rect 627087 54270 627198 54275
rect 627087 54214 627092 54270
rect 627148 54214 627198 54270
rect 627087 54212 627198 54214
rect 629583 54272 629649 54275
rect 635055 54272 635121 54275
rect 629583 54270 635121 54272
rect 629583 54214 629588 54270
rect 629644 54214 635060 54270
rect 635116 54214 635121 54270
rect 629583 54212 635121 54214
rect 627087 54209 627153 54212
rect 629583 54209 629649 54212
rect 635055 54209 635121 54212
rect 212559 54124 212625 54127
rect 208770 54122 212625 54124
rect 208770 54066 212564 54122
rect 212620 54066 212625 54122
rect 208770 54064 212625 54066
rect 208064 54062 208070 54064
rect 208527 54061 208593 54064
rect 212559 54061 212625 54064
rect 632943 54124 633009 54127
rect 636399 54124 636465 54127
rect 632943 54122 636465 54124
rect 632943 54066 632948 54122
rect 633004 54066 636404 54122
rect 636460 54066 636465 54122
rect 632943 54064 636465 54066
rect 632943 54061 633009 54064
rect 636399 54061 636465 54064
rect 207610 53914 207616 53978
rect 207680 53976 207686 53978
rect 208143 53976 208209 53979
rect 207680 53974 208209 53976
rect 207680 53918 208148 53974
rect 208204 53918 208209 53974
rect 207680 53916 208209 53918
rect 207680 53914 207686 53916
rect 208143 53913 208209 53916
rect 628527 53976 628593 53979
rect 634863 53976 634929 53979
rect 628527 53974 634929 53976
rect 628527 53918 628532 53974
rect 628588 53918 634868 53974
rect 634924 53918 634929 53974
rect 628527 53916 634929 53918
rect 628527 53913 628593 53916
rect 634863 53913 634929 53916
rect 204730 53766 204736 53830
rect 204800 53828 204806 53830
rect 210735 53828 210801 53831
rect 204800 53826 210801 53828
rect 204800 53770 210740 53826
rect 210796 53770 210801 53826
rect 204800 53768 210801 53770
rect 204800 53766 204806 53768
rect 210735 53765 210801 53768
rect 630639 53828 630705 53831
rect 636303 53828 636369 53831
rect 630639 53826 636369 53828
rect 630639 53770 630644 53826
rect 630700 53770 636308 53826
rect 636364 53770 636369 53826
rect 630639 53768 636369 53770
rect 630639 53765 630705 53768
rect 636303 53765 636369 53768
rect 206650 53618 206656 53682
rect 206720 53680 206726 53682
rect 206720 53646 207150 53680
rect 206720 53641 207153 53646
rect 206720 53620 207092 53641
rect 206720 53618 206726 53620
rect 207087 53585 207092 53620
rect 207148 53585 207153 53641
rect 207087 53580 207153 53585
rect 203535 53532 203601 53535
rect 206703 53532 206769 53535
rect 203535 53530 206769 53532
rect 203535 53474 203540 53530
rect 203596 53474 206708 53530
rect 206764 53474 206769 53530
rect 203535 53472 206769 53474
rect 203535 53469 203601 53472
rect 206703 53469 206769 53472
rect 207226 53470 207232 53534
rect 207296 53532 207302 53534
rect 207567 53532 207633 53535
rect 207296 53530 207633 53532
rect 207296 53474 207572 53530
rect 207628 53474 207633 53530
rect 207296 53472 207633 53474
rect 207296 53470 207302 53472
rect 207567 53469 207633 53472
rect 207802 53470 207808 53534
rect 207872 53532 207878 53534
rect 209007 53532 209073 53535
rect 207872 53530 209073 53532
rect 207872 53474 209012 53530
rect 209068 53474 209073 53530
rect 207872 53472 209073 53474
rect 207872 53470 207878 53472
rect 209007 53469 209073 53472
rect 212559 53532 212625 53535
rect 214479 53532 214545 53535
rect 212559 53530 214545 53532
rect 212559 53474 212564 53530
rect 212620 53474 214484 53530
rect 214540 53474 214545 53530
rect 212559 53472 214545 53474
rect 212559 53469 212625 53472
rect 214479 53469 214545 53472
rect 202863 53384 202929 53387
rect 206895 53384 206961 53387
rect 202863 53382 206961 53384
rect 202863 53326 202868 53382
rect 202924 53326 206900 53382
rect 206956 53326 206961 53382
rect 202863 53324 206961 53326
rect 202863 53321 202929 53324
rect 206895 53321 206961 53324
rect 207034 53322 207040 53386
rect 207104 53384 207110 53386
rect 209295 53384 209361 53387
rect 207104 53382 209361 53384
rect 207104 53326 209300 53382
rect 209356 53326 209361 53382
rect 207104 53324 209361 53326
rect 207104 53322 207110 53324
rect 209295 53321 209361 53324
rect 204922 53174 204928 53238
rect 204992 53236 204998 53238
rect 471034 53236 471040 53238
rect 204992 53176 471040 53236
rect 204992 53174 204998 53176
rect 471034 53174 471040 53176
rect 471104 53174 471110 53238
rect 204303 53088 204369 53091
rect 205839 53088 205905 53091
rect 204303 53086 205905 53088
rect 204303 53030 204308 53086
rect 204364 53030 205844 53086
rect 205900 53030 205905 53086
rect 204303 53028 205905 53030
rect 204303 53025 204369 53028
rect 205839 53025 205905 53028
rect 206703 53088 206769 53091
rect 218319 53088 218385 53091
rect 206703 53086 218385 53088
rect 206703 53030 206708 53086
rect 206764 53030 218324 53086
rect 218380 53030 218385 53086
rect 206703 53028 218385 53030
rect 206703 53025 206769 53028
rect 218319 53025 218385 53028
rect 203919 52940 203985 52943
rect 213711 52940 213777 52943
rect 203919 52938 213777 52940
rect 203919 52882 203924 52938
rect 203980 52882 213716 52938
rect 213772 52882 213777 52938
rect 203919 52880 213777 52882
rect 203919 52877 203985 52880
rect 213711 52877 213777 52880
rect 203055 52792 203121 52795
rect 220527 52792 220593 52795
rect 203055 52790 220593 52792
rect 203055 52734 203060 52790
rect 203116 52734 220532 52790
rect 220588 52734 220593 52790
rect 203055 52732 220593 52734
rect 203055 52729 203121 52732
rect 220527 52729 220593 52732
rect 203151 52644 203217 52647
rect 220239 52644 220305 52647
rect 203151 52642 220305 52644
rect 203151 52586 203156 52642
rect 203212 52586 220244 52642
rect 220300 52586 220305 52642
rect 203151 52584 220305 52586
rect 203151 52581 203217 52584
rect 220239 52581 220305 52584
rect 204154 52434 204160 52498
rect 204224 52496 204230 52498
rect 218031 52496 218097 52499
rect 204224 52494 218097 52496
rect 204224 52438 218036 52494
rect 218092 52438 218097 52494
rect 204224 52436 218097 52438
rect 204224 52434 204230 52436
rect 218031 52433 218097 52436
rect 207855 52348 207921 52351
rect 208186 52348 208192 52350
rect 207855 52346 208192 52348
rect 207855 52290 207860 52346
rect 207916 52290 208192 52346
rect 207855 52288 208192 52290
rect 207855 52285 207921 52288
rect 208186 52286 208192 52288
rect 208256 52286 208262 52350
rect 205647 52200 205713 52203
rect 632698 52200 632704 52202
rect 205647 52198 632704 52200
rect 205647 52142 205652 52198
rect 205708 52142 632704 52198
rect 205647 52140 632704 52142
rect 205647 52137 205713 52140
rect 632698 52138 632704 52140
rect 632768 52138 632774 52202
rect 206799 52052 206865 52055
rect 632890 52052 632896 52054
rect 206799 52050 632896 52052
rect 206799 51994 206804 52050
rect 206860 51994 632896 52050
rect 206799 51992 632896 51994
rect 206799 51989 206865 51992
rect 632890 51990 632896 51992
rect 632960 51990 632966 52054
rect 204346 51842 204352 51906
rect 204416 51904 204422 51906
rect 204687 51904 204753 51907
rect 204416 51902 204753 51904
rect 204416 51846 204692 51902
rect 204748 51846 204753 51902
rect 204416 51844 204753 51846
rect 204416 51842 204422 51844
rect 204687 51841 204753 51844
rect 214959 51904 215025 51907
rect 633274 51904 633280 51906
rect 214959 51902 633280 51904
rect 214959 51846 214964 51902
rect 215020 51846 633280 51902
rect 214959 51844 633280 51846
rect 214959 51841 215025 51844
rect 633274 51842 633280 51844
rect 633344 51842 633350 51906
rect 218223 51756 218289 51759
rect 632506 51756 632512 51758
rect 218223 51754 632512 51756
rect 218223 51698 218228 51754
rect 218284 51698 632512 51754
rect 218223 51696 632512 51698
rect 218223 51693 218289 51696
rect 632506 51694 632512 51696
rect 632576 51694 632582 51758
rect 145594 51250 145600 51314
rect 145664 51312 145670 51314
rect 242991 51312 243057 51315
rect 145664 51310 243057 51312
rect 145664 51254 242996 51310
rect 243052 51254 243057 51310
rect 145664 51252 243057 51254
rect 145664 51250 145670 51252
rect 242991 51249 243057 51252
rect 145978 51102 145984 51166
rect 146048 51164 146054 51166
rect 239823 51164 239889 51167
rect 146048 51162 239889 51164
rect 146048 51106 239828 51162
rect 239884 51106 239889 51162
rect 146048 51104 239889 51106
rect 146048 51102 146054 51104
rect 239823 51101 239889 51104
rect 145786 50954 145792 51018
rect 145856 51016 145862 51018
rect 242031 51016 242097 51019
rect 145856 51014 242097 51016
rect 145856 50958 242036 51014
rect 242092 50958 242097 51014
rect 145856 50956 242097 50958
rect 145856 50954 145862 50956
rect 242031 50953 242097 50956
rect 145402 50806 145408 50870
rect 145472 50868 145478 50870
rect 244143 50868 244209 50871
rect 145472 50866 244209 50868
rect 145472 50810 244148 50866
rect 244204 50810 244209 50866
rect 145472 50808 244209 50810
rect 145472 50806 145478 50808
rect 244143 50805 244209 50808
rect 264879 50424 264945 50427
rect 632314 50424 632320 50426
rect 264879 50422 632320 50424
rect 264879 50366 264884 50422
rect 264940 50366 632320 50422
rect 264879 50364 632320 50366
rect 264879 50361 264945 50364
rect 632314 50362 632320 50364
rect 632384 50362 632390 50426
rect 217455 48944 217521 48947
rect 632122 48944 632128 48946
rect 217455 48942 632128 48944
rect 217455 48886 217460 48942
rect 217516 48886 632128 48942
rect 217455 48884 632128 48886
rect 217455 48881 217521 48884
rect 632122 48882 632128 48884
rect 632192 48882 632198 48946
rect 217071 48796 217137 48799
rect 633466 48796 633472 48798
rect 217071 48794 633472 48796
rect 217071 48738 217076 48794
rect 217132 48738 633472 48794
rect 217071 48736 633472 48738
rect 217071 48733 217137 48736
rect 633466 48734 633472 48736
rect 633536 48734 633542 48798
rect 148239 48648 148305 48651
rect 243759 48648 243825 48651
rect 148239 48646 243825 48648
rect 148239 48590 148244 48646
rect 148300 48590 243764 48646
rect 243820 48590 243825 48646
rect 148239 48588 243825 48590
rect 148239 48585 148305 48588
rect 243759 48585 243825 48588
rect 148431 48500 148497 48503
rect 243375 48500 243441 48503
rect 148431 48498 243441 48500
rect 148431 48442 148436 48498
rect 148492 48442 243380 48498
rect 243436 48442 243441 48498
rect 148431 48440 243441 48442
rect 148431 48437 148497 48440
rect 243375 48437 243441 48440
rect 148623 48352 148689 48355
rect 242415 48352 242481 48355
rect 148623 48350 242481 48352
rect 148623 48294 148628 48350
rect 148684 48294 242420 48350
rect 242476 48294 242481 48350
rect 148623 48292 242481 48294
rect 148623 48289 148689 48292
rect 242415 48289 242481 48292
rect 149199 48204 149265 48207
rect 239343 48204 239409 48207
rect 149199 48202 239409 48204
rect 149199 48146 149204 48202
rect 149260 48146 239348 48202
rect 239404 48146 239409 48202
rect 149199 48144 239409 48146
rect 149199 48141 149265 48144
rect 239343 48141 239409 48144
rect 149391 48056 149457 48059
rect 238575 48056 238641 48059
rect 149391 48054 238641 48056
rect 149391 47998 149396 48054
rect 149452 47998 238580 48054
rect 238636 47998 238641 48054
rect 149391 47996 238641 47998
rect 149391 47993 149457 47996
rect 238575 47993 238641 47996
rect 149583 47908 149649 47911
rect 236751 47908 236817 47911
rect 149583 47906 236817 47908
rect 149583 47850 149588 47906
rect 149644 47850 236756 47906
rect 236812 47850 236817 47906
rect 149583 47848 236817 47850
rect 149583 47845 149649 47848
rect 236751 47845 236817 47848
rect 148047 47760 148113 47763
rect 241551 47760 241617 47763
rect 148047 47758 241617 47760
rect 148047 47702 148052 47758
rect 148108 47702 241556 47758
rect 241612 47702 241617 47758
rect 148047 47700 241617 47702
rect 148047 47697 148113 47700
rect 241551 47697 241617 47700
rect 148815 47612 148881 47615
rect 240207 47612 240273 47615
rect 148815 47610 240273 47612
rect 148815 47554 148820 47610
rect 148876 47554 240212 47610
rect 240268 47554 240273 47610
rect 148815 47552 240273 47554
rect 148815 47549 148881 47552
rect 240207 47549 240273 47552
rect 161295 46724 161361 46727
rect 181359 46724 181425 46727
rect 161295 46722 181425 46724
rect 161295 46666 161300 46722
rect 161356 46666 181364 46722
rect 181420 46666 181425 46722
rect 161295 46664 181425 46666
rect 161295 46661 161361 46664
rect 181359 46661 181425 46664
rect 207951 46576 208017 46579
rect 208527 46576 208593 46579
rect 207951 46574 208593 46576
rect 207951 46518 207956 46574
rect 208012 46518 208532 46574
rect 208588 46518 208593 46574
rect 207951 46516 208593 46518
rect 207951 46513 208017 46516
rect 208527 46513 208593 46516
rect 207855 46428 207921 46431
rect 209679 46428 209745 46431
rect 207855 46426 209745 46428
rect 207855 46370 207860 46426
rect 207916 46370 209684 46426
rect 209740 46370 209745 46426
rect 207855 46368 209745 46370
rect 207855 46365 207921 46368
rect 209679 46365 209745 46368
rect 206223 45540 206289 45543
rect 302458 45540 302464 45542
rect 206223 45538 302464 45540
rect 206223 45482 206228 45538
rect 206284 45482 302464 45538
rect 206223 45480 302464 45482
rect 206223 45477 206289 45480
rect 302458 45478 302464 45480
rect 302528 45478 302534 45542
rect 205071 45392 205137 45395
rect 305338 45392 305344 45394
rect 205071 45390 305344 45392
rect 205071 45334 205076 45390
rect 205132 45334 305344 45390
rect 205071 45332 305344 45334
rect 205071 45329 205137 45332
rect 305338 45330 305344 45332
rect 305408 45330 305414 45394
rect 206127 45244 206193 45247
rect 356986 45244 356992 45246
rect 206127 45242 356992 45244
rect 206127 45186 206132 45242
rect 206188 45186 356992 45242
rect 206127 45184 356992 45186
rect 206127 45181 206193 45184
rect 356986 45182 356992 45184
rect 357056 45182 357062 45246
rect 205455 45096 205521 45099
rect 360058 45096 360064 45098
rect 205455 45094 360064 45096
rect 205455 45038 205460 45094
rect 205516 45038 360064 45094
rect 205455 45036 360064 45038
rect 205455 45033 205521 45036
rect 360058 45034 360064 45036
rect 360128 45034 360134 45098
rect 205743 44948 205809 44951
rect 362938 44948 362944 44950
rect 205743 44946 362944 44948
rect 205743 44890 205748 44946
rect 205804 44890 362944 44946
rect 205743 44888 362944 44890
rect 205743 44885 205809 44888
rect 362938 44886 362944 44888
rect 363008 44886 363014 44950
rect 206319 44800 206385 44803
rect 465615 44800 465681 44803
rect 206319 44798 465681 44800
rect 206319 44742 206324 44798
rect 206380 44742 465620 44798
rect 465676 44742 465681 44798
rect 206319 44740 465681 44742
rect 206319 44737 206385 44740
rect 465615 44737 465681 44740
rect 208815 44652 208881 44655
rect 521583 44652 521649 44655
rect 208815 44650 521649 44652
rect 208815 44594 208820 44650
rect 208876 44594 521588 44650
rect 521644 44594 521649 44650
rect 208815 44592 521649 44594
rect 208815 44589 208881 44592
rect 521583 44589 521649 44592
rect 302511 43322 302577 43323
rect 302458 43320 302464 43322
rect 302420 43260 302464 43320
rect 302528 43318 302577 43322
rect 302572 43262 302577 43318
rect 302458 43258 302464 43260
rect 302528 43258 302577 43262
rect 305338 43258 305344 43322
rect 305408 43320 305414 43322
rect 306735 43320 306801 43323
rect 305408 43318 306801 43320
rect 305408 43262 306740 43318
rect 306796 43262 306801 43318
rect 305408 43260 306801 43262
rect 305408 43258 305414 43260
rect 302511 43257 302577 43258
rect 306735 43257 306801 43260
rect 360058 43258 360064 43322
rect 360128 43320 360134 43322
rect 361743 43320 361809 43323
rect 360128 43318 361809 43320
rect 360128 43262 361748 43318
rect 361804 43262 361809 43318
rect 360128 43260 361809 43262
rect 360128 43258 360134 43260
rect 361743 43257 361809 43260
rect 362938 43258 362944 43322
rect 363008 43320 363014 43322
rect 364911 43320 364977 43323
rect 363008 43318 364977 43320
rect 363008 43262 364916 43318
rect 364972 43262 364977 43318
rect 363008 43260 364977 43262
rect 363008 43258 363014 43260
rect 364911 43257 364977 43260
rect 356986 43110 356992 43174
rect 357056 43172 357062 43174
rect 357135 43172 357201 43175
rect 357056 43170 357201 43172
rect 357056 43114 357140 43170
rect 357196 43114 357201 43170
rect 357056 43112 357201 43114
rect 357056 43110 357062 43112
rect 357135 43109 357201 43112
rect 523887 43172 523953 43175
rect 529263 43172 529329 43175
rect 523887 43170 529329 43172
rect 523887 43114 523892 43170
rect 523948 43114 529268 43170
rect 529324 43114 529329 43170
rect 523887 43112 529329 43114
rect 523887 43109 523953 43112
rect 529263 43109 529329 43112
rect 408879 42136 408945 42139
rect 416271 42136 416337 42139
rect 471087 42138 471153 42139
rect 471034 42136 471040 42138
rect 408879 42134 416337 42136
rect 408879 42078 408884 42134
rect 408940 42078 416276 42134
rect 416332 42078 416337 42134
rect 408879 42076 416337 42078
rect 470996 42076 471040 42136
rect 471104 42134 471153 42138
rect 471148 42078 471153 42134
rect 408879 42073 408945 42076
rect 416271 42073 416337 42076
rect 471034 42074 471040 42076
rect 471104 42074 471153 42078
rect 471087 42073 471153 42074
rect 521199 42136 521265 42139
rect 525903 42136 525969 42139
rect 521199 42134 525969 42136
rect 521199 42078 521204 42134
rect 521260 42078 525908 42134
rect 525964 42078 525969 42134
rect 521199 42076 525969 42078
rect 521199 42073 521265 42076
rect 525903 42073 525969 42076
rect 187599 41840 187665 41843
rect 189946 41840 189952 41842
rect 187599 41838 189952 41840
rect 187599 41782 187604 41838
rect 187660 41782 189952 41838
rect 187599 41780 189952 41782
rect 187599 41777 187665 41780
rect 189946 41778 189952 41780
rect 190016 41778 190022 41842
rect 194319 41840 194385 41843
rect 194938 41840 194944 41842
rect 194319 41838 194944 41840
rect 194319 41782 194324 41838
rect 194380 41782 194944 41838
rect 194319 41780 194944 41782
rect 194319 41777 194385 41780
rect 194938 41778 194944 41780
rect 195008 41778 195014 41842
rect 406287 41840 406353 41843
rect 410799 41840 410865 41843
rect 518511 41842 518577 41843
rect 518458 41840 518464 41842
rect 406287 41838 410865 41840
rect 406287 41782 406292 41838
rect 406348 41782 410804 41838
rect 410860 41782 410865 41838
rect 406287 41780 410865 41782
rect 518420 41780 518464 41840
rect 518528 41838 518577 41842
rect 518572 41782 518577 41838
rect 406287 41777 406353 41780
rect 410799 41777 410865 41780
rect 518458 41778 518464 41780
rect 518528 41778 518577 41782
rect 518511 41777 518577 41778
rect 189946 40742 189952 40806
rect 190016 40804 190022 40806
rect 204879 40804 204945 40807
rect 190016 40802 204945 40804
rect 190016 40746 204884 40802
rect 204940 40746 204945 40802
rect 190016 40744 204945 40746
rect 190016 40742 190022 40744
rect 204879 40741 204945 40744
rect 512559 40804 512625 40807
rect 518266 40804 518272 40806
rect 512559 40802 518272 40804
rect 512559 40746 512564 40802
rect 512620 40746 518272 40802
rect 512559 40744 518272 40746
rect 512559 40741 512625 40744
rect 518266 40742 518272 40744
rect 518336 40742 518342 40806
rect 194938 40594 194944 40658
rect 195008 40656 195014 40658
rect 613455 40656 613521 40659
rect 195008 40654 613521 40656
rect 195008 40598 613460 40654
rect 613516 40598 613521 40654
rect 195008 40596 613521 40598
rect 195008 40594 195014 40596
rect 613455 40593 613521 40596
rect 138159 40212 138225 40215
rect 138159 40210 141822 40212
rect 138159 40154 138164 40210
rect 138220 40154 141822 40210
rect 138159 40152 141822 40154
rect 138159 40149 138225 40152
rect 141762 39886 141822 40152
<< via3 >>
rect 385984 996082 386048 996146
rect 385984 995490 386048 995554
rect 294784 993566 294848 993630
rect 294784 992086 294848 992150
rect 40576 968702 40640 968766
rect 675520 967518 675584 967582
rect 41728 967134 41792 967138
rect 41728 967078 41780 967134
rect 41780 967078 41792 967134
rect 41728 967074 41792 967078
rect 674560 965594 674624 965658
rect 675904 965594 675968 965658
rect 40384 965002 40448 965066
rect 674752 964854 674816 964918
rect 40768 963966 40832 964030
rect 40960 963374 41024 963438
rect 41152 962782 41216 962846
rect 674944 962782 675008 962846
rect 674368 962486 674432 962550
rect 41536 962190 41600 962254
rect 42880 962190 42944 962254
rect 675328 962250 675392 962254
rect 675328 962194 675380 962250
rect 675380 962194 675392 962250
rect 675328 962190 675392 962194
rect 43072 962042 43136 962106
rect 676672 961450 676736 961514
rect 675520 961066 675584 961070
rect 675520 961010 675532 961066
rect 675532 961010 675584 961066
rect 675520 961006 675584 961010
rect 675712 960178 675776 960182
rect 675712 960122 675724 960178
rect 675724 960122 675776 960178
rect 675712 960118 675776 960122
rect 41344 959674 41408 959738
rect 41920 959142 41984 959146
rect 41920 959086 41932 959142
rect 41932 959086 41984 959142
rect 41920 959082 41984 959086
rect 42112 958402 42176 958406
rect 42112 958346 42124 958402
rect 42124 958346 42176 958402
rect 42112 958342 42176 958346
rect 42304 957750 42368 957814
rect 676480 957602 676544 957666
rect 42496 956122 42560 956186
rect 675136 955974 675200 956038
rect 677056 953458 677120 953522
rect 676864 953310 676928 953374
rect 674752 940878 674816 940942
rect 674560 938806 674624 938870
rect 674944 938362 675008 938426
rect 675904 935846 675968 935910
rect 674368 934662 674432 934726
rect 675328 934514 675392 934578
rect 675136 933626 675200 933690
rect 676480 932590 676544 932654
rect 676672 931850 676736 931914
rect 677056 931406 677120 931470
rect 676864 930222 676928 930286
rect 42880 907134 42944 907198
rect 42688 903286 42752 903350
rect 42496 902990 42560 903054
rect 41728 902250 41792 902314
rect 42304 900622 42368 900686
rect 41536 899734 41600 899798
rect 40576 899142 40640 899206
rect 42112 897514 42176 897578
rect 41920 896626 41984 896690
rect 40384 895590 40448 895654
rect 40960 894998 41024 895062
rect 41344 894406 41408 894470
rect 41152 893518 41216 893582
rect 40768 892482 40832 892546
rect 42880 887154 42944 887218
rect 674368 876350 674432 876414
rect 676672 876350 676736 876414
rect 674752 876202 674816 876266
rect 675712 875758 675776 875822
rect 674944 873982 675008 874046
rect 674560 873390 674624 873454
rect 674176 872798 674240 872862
rect 675520 872414 675584 872418
rect 675520 872358 675572 872414
rect 675572 872358 675584 872414
rect 675520 872354 675584 872358
rect 675328 869898 675392 869902
rect 675328 869842 675380 869898
rect 675380 869842 675392 869898
rect 675328 869838 675392 869842
rect 675136 866878 675200 866942
rect 42304 866434 42368 866498
rect 42880 866434 42944 866498
rect 675520 864718 675584 864722
rect 675520 864662 675532 864718
rect 675532 864662 675584 864718
rect 675520 864658 675584 864662
rect 42688 864214 42752 864278
rect 42688 864066 42752 864130
rect 675712 862942 675776 862946
rect 675712 862886 675724 862942
rect 675724 862886 675776 862942
rect 675712 862882 675776 862886
rect 42496 858146 42560 858210
rect 43264 857998 43328 858062
rect 42688 852670 42752 852734
rect 40000 842606 40064 842670
rect 43072 840978 43136 841042
rect 43072 840682 43136 840746
rect 42880 830914 42944 830978
rect 43264 830914 43328 830978
rect 40000 827570 40064 827574
rect 40000 827514 40012 827570
rect 40012 827514 40064 827570
rect 40000 827510 40064 827514
rect 40768 818334 40832 818398
rect 41344 802054 41408 802118
rect 41536 801906 41600 801970
rect 42688 800426 42752 800490
rect 41728 800338 41792 800342
rect 41728 800282 41780 800338
rect 41780 800282 41792 800338
rect 41728 800278 41792 800282
rect 42112 800338 42176 800342
rect 42112 800282 42124 800338
rect 42124 800282 42176 800338
rect 42112 800278 42176 800282
rect 42304 800042 42368 800046
rect 42304 799986 42316 800042
rect 42316 799986 42368 800042
rect 42304 799982 42368 799986
rect 42304 797910 42368 797974
rect 42688 794862 42752 794866
rect 42688 794806 42740 794862
rect 42740 794806 42752 794862
rect 42688 794802 42752 794806
rect 41728 794270 41792 794274
rect 41728 794214 41780 794270
rect 41780 794214 41792 794270
rect 41728 794210 41792 794214
rect 41728 794062 41792 794126
rect 43072 794062 43136 794126
rect 42112 792138 42176 792202
rect 41536 791842 41600 791906
rect 41344 791694 41408 791758
rect 41728 791162 41792 791166
rect 41728 791106 41780 791162
rect 41780 791106 41792 791162
rect 41728 791102 41792 791106
rect 41920 790954 41984 791018
rect 42496 790954 42560 791018
rect 676288 787846 676352 787910
rect 673984 787402 674048 787466
rect 675904 786662 675968 786726
rect 676096 784146 676160 784210
rect 676480 781926 676544 781990
rect 677056 780446 677120 780510
rect 677056 777486 677120 777550
rect 676864 777338 676928 777402
rect 40768 775118 40832 775182
rect 676864 773046 676928 773110
rect 677824 773046 677888 773110
rect 676864 772898 676928 772962
rect 677248 772898 677312 772962
rect 677248 772602 677312 772666
rect 42304 763130 42368 763194
rect 42304 762686 42368 762750
rect 674752 762390 674816 762454
rect 42112 761798 42176 761862
rect 675520 761650 675584 761714
rect 674368 760244 674432 760308
rect 40960 760170 41024 760234
rect 674944 760022 675008 760086
rect 40384 759578 40448 759642
rect 675328 759134 675392 759198
rect 41152 758542 41216 758606
rect 675712 758542 675776 758606
rect 676672 757358 676736 757422
rect 42304 757062 42368 757126
rect 674560 756914 674624 756978
rect 674176 755434 674240 755498
rect 675136 755286 675200 755350
rect 41152 754842 41216 754906
rect 677248 754398 677312 754462
rect 42304 754250 42368 754314
rect 676864 753806 676928 753870
rect 677824 752918 677888 752982
rect 42688 751882 42752 751946
rect 42688 751646 42752 751650
rect 42688 751590 42740 751646
rect 42740 751590 42752 751646
rect 42688 751586 42752 751590
rect 41728 748686 41792 748690
rect 41728 748630 41780 748686
rect 41780 748630 41792 748686
rect 41728 748626 41792 748630
rect 41920 747354 41984 747358
rect 41920 747298 41972 747354
rect 41972 747298 41984 747354
rect 41920 747294 41984 747298
rect 40384 747146 40448 747210
rect 40960 746850 41024 746914
rect 674368 743298 674432 743362
rect 676672 741670 676736 741734
rect 674176 741374 674240 741438
rect 675520 740398 675584 740402
rect 675520 740342 675532 740398
rect 675532 740342 675584 740398
rect 675520 740338 675584 740342
rect 674752 739302 674816 739366
rect 675328 738622 675392 738626
rect 675328 738566 675380 738622
rect 675380 738566 675392 738622
rect 675328 738562 675392 738566
rect 676480 736638 676544 736702
rect 675712 734478 675776 734482
rect 675712 734422 675724 734478
rect 675724 734422 675776 734478
rect 675712 734418 675776 734422
rect 41728 733826 41792 733890
rect 40576 733086 40640 733150
rect 40768 733086 40832 733150
rect 676864 732494 676928 732558
rect 41152 732198 41216 732262
rect 41344 729534 41408 729598
rect 40960 726278 41024 726342
rect 42496 721542 42560 721606
rect 43072 721394 43136 721458
rect 675904 717065 675968 717129
rect 41728 716126 41792 716130
rect 41728 716070 41780 716126
rect 41780 716070 41792 716126
rect 41728 716066 41792 716070
rect 676288 715770 676352 715834
rect 42112 713994 42176 714058
rect 42304 713846 42368 713910
rect 673984 712070 674048 712134
rect 676096 711922 676160 711986
rect 42880 711834 42944 711838
rect 42880 711778 42932 711834
rect 42932 711778 42944 711834
rect 42880 711774 42944 711778
rect 42112 711686 42176 711690
rect 42112 711630 42124 711686
rect 42124 711630 42176 711686
rect 42112 711626 42176 711630
rect 42688 711626 42752 711690
rect 41536 711330 41600 711394
rect 42688 711182 42752 711246
rect 41728 711034 41792 711098
rect 42304 711034 42368 711098
rect 43072 708518 43136 708582
rect 677056 708370 677120 708434
rect 42880 707778 42944 707842
rect 42496 707334 42560 707398
rect 41920 706506 41984 706510
rect 41920 706450 41972 706506
rect 41972 706450 41984 706506
rect 41920 706446 41984 706450
rect 41728 704966 41792 705030
rect 41536 704670 41600 704734
rect 42112 704138 42176 704142
rect 42112 704082 42124 704138
rect 42124 704082 42176 704138
rect 42112 704078 42176 704082
rect 41344 703634 41408 703698
rect 40960 703486 41024 703550
rect 675136 697862 675200 697926
rect 673984 697270 674048 697334
rect 674944 696826 675008 696890
rect 676096 694754 676160 694818
rect 674560 694606 674624 694670
rect 675904 693422 675968 693486
rect 41536 692682 41600 692746
rect 676480 691646 676544 691710
rect 40576 689574 40640 689638
rect 41152 689574 41216 689638
rect 676672 689278 676736 689342
rect 676672 689130 676736 689194
rect 42112 688686 42176 688750
rect 677056 688242 677120 688306
rect 41152 686318 41216 686382
rect 677056 685578 677120 685642
rect 42496 684838 42560 684902
rect 40960 683210 41024 683274
rect 42880 682914 42944 682978
rect 676288 679658 676352 679722
rect 42304 678326 42368 678390
rect 41344 674834 41408 674838
rect 41344 674778 41396 674834
rect 41396 674778 41408 674834
rect 41344 674774 41408 674778
rect 676288 672258 676352 672322
rect 41728 670926 41792 670990
rect 42688 670986 42752 670990
rect 42688 670930 42700 670986
rect 42700 670930 42752 670986
rect 42688 670926 42752 670930
rect 43072 670986 43136 670990
rect 43072 670930 43084 670986
rect 43084 670930 43136 670986
rect 43072 670926 43136 670930
rect 674368 670038 674432 670102
rect 675520 669742 675584 669806
rect 42496 668914 42560 668918
rect 42496 668858 42548 668914
rect 42548 668858 42560 668914
rect 42496 668854 42560 668858
rect 41728 668470 41792 668474
rect 41728 668414 41780 668470
rect 41780 668414 41792 668470
rect 41728 668410 41792 668414
rect 42304 668262 42368 668326
rect 674176 666930 674240 666994
rect 674752 666634 674816 666698
rect 42880 666546 42944 666550
rect 42880 666490 42932 666546
rect 42932 666490 42944 666546
rect 42880 666486 42944 666490
rect 675328 665894 675392 665958
rect 41344 665746 41408 665810
rect 41344 665598 41408 665662
rect 43072 665302 43136 665366
rect 675712 664266 675776 664330
rect 677248 663526 677312 663590
rect 42688 663378 42752 663442
rect 676864 662342 676928 662406
rect 41344 661306 41408 661370
rect 41728 661366 41792 661370
rect 41728 661310 41780 661366
rect 41780 661310 41792 661366
rect 41728 661306 41792 661310
rect 41920 661070 41984 661074
rect 41920 661014 41932 661070
rect 41932 661014 41984 661070
rect 41920 661010 41984 661014
rect 40960 660862 41024 660926
rect 675712 659382 675776 659446
rect 676672 659382 676736 659446
rect 675520 659234 675584 659298
rect 676480 659234 676544 659298
rect 41152 656126 41216 656190
rect 675520 652722 675584 652786
rect 675520 652634 675584 652638
rect 675520 652578 675532 652634
rect 675532 652578 675584 652634
rect 675520 652574 675584 652578
rect 674752 652130 674816 652194
rect 675328 651006 675392 651010
rect 675328 650950 675340 651006
rect 675340 650950 675392 651006
rect 675328 650946 675392 650950
rect 676288 649614 676352 649678
rect 673984 648430 674048 648494
rect 676480 648430 676544 648494
rect 674176 648282 674240 648346
rect 42112 646654 42176 646718
rect 40576 646358 40640 646422
rect 674368 645470 674432 645534
rect 675904 645026 675968 645090
rect 676864 644878 676928 644942
rect 40768 643102 40832 643166
rect 675136 641918 675200 641982
rect 675712 640734 675776 640798
rect 676672 640734 676736 640798
rect 676480 640438 676544 640502
rect 676480 640290 676544 640354
rect 40960 639994 41024 640058
rect 674752 639846 674816 639910
rect 674944 639402 675008 639466
rect 675136 638514 675200 638578
rect 674368 637774 674432 637838
rect 42880 635850 42944 635914
rect 41536 635110 41600 635174
rect 676864 634962 676928 635026
rect 42496 634370 42560 634434
rect 676096 633246 676160 633250
rect 676096 633190 676108 633246
rect 676108 633190 676160 633246
rect 676096 633186 676160 633190
rect 674176 630374 674240 630438
rect 676864 630374 676928 630438
rect 676096 630078 676160 630142
rect 676672 630138 676736 630142
rect 676672 630082 676724 630138
rect 676724 630082 676736 630138
rect 676672 630078 676736 630082
rect 41344 627710 41408 627774
rect 42304 627562 42368 627626
rect 42112 627414 42176 627478
rect 674752 627266 674816 627330
rect 41344 625194 41408 625258
rect 673984 624958 674048 624962
rect 673984 624902 674036 624958
rect 674036 624902 674048 624958
rect 673984 624898 674048 624902
rect 42112 624454 42176 624518
rect 41536 624306 41600 624370
rect 42112 624306 42176 624370
rect 42496 622086 42560 622150
rect 674560 621642 674624 621706
rect 42112 620962 42176 620966
rect 42112 620906 42124 620962
rect 42124 620906 42176 620962
rect 42112 620902 42176 620906
rect 676672 620902 676736 620966
rect 42304 620754 42368 620818
rect 41728 619186 41792 619190
rect 41728 619130 41780 619186
rect 41780 619130 41792 619186
rect 41728 619126 41792 619130
rect 674176 618830 674240 618894
rect 41920 618298 41984 618302
rect 41920 618242 41932 618298
rect 41932 618242 41984 618298
rect 41920 618238 41984 618242
rect 42880 618298 42944 618302
rect 42880 618242 42892 618298
rect 42892 618242 42944 618298
rect 42880 618238 42944 618242
rect 40768 618090 40832 618154
rect 677056 617794 677120 617858
rect 40960 617646 41024 617710
rect 674368 607730 674432 607794
rect 674560 607434 674624 607498
rect 675712 606458 675776 606462
rect 675712 606402 675724 606458
rect 675724 606402 675776 606458
rect 675712 606398 675776 606402
rect 673984 604918 674048 604982
rect 674176 604770 674240 604834
rect 40576 603882 40640 603946
rect 42112 603142 42176 603206
rect 675904 600182 675968 600246
rect 40576 599886 40640 599950
rect 674944 599146 675008 599210
rect 676096 599146 676160 599210
rect 40960 596778 41024 596842
rect 676672 595298 676736 595362
rect 676096 593374 676160 593438
rect 43072 586566 43136 586630
rect 42496 584998 42560 585002
rect 42496 584942 42548 584998
rect 42548 584942 42560 584998
rect 42496 584938 42560 584942
rect 41344 584494 41408 584558
rect 41536 584346 41600 584410
rect 42880 584406 42944 584410
rect 42880 584350 42932 584406
rect 42932 584350 42944 584406
rect 42880 584346 42944 584350
rect 42304 584198 42368 584262
rect 673984 584494 674048 584558
rect 674176 584554 674240 584558
rect 674176 584498 674228 584554
rect 674228 584498 674240 584554
rect 674176 584494 674240 584498
rect 673984 584050 674048 584114
rect 676864 581830 676928 581894
rect 675328 581682 675392 581746
rect 42304 581238 42368 581302
rect 676480 581238 676544 581302
rect 675520 580350 675584 580414
rect 676288 579610 676352 579674
rect 42880 578338 42944 578342
rect 42880 578282 42932 578338
rect 42932 578282 42944 578338
rect 42880 578278 42944 578282
rect 674944 578130 675008 578194
rect 675136 578130 675200 578194
rect 43072 577598 43136 577602
rect 43072 577542 43084 577598
rect 43084 577542 43136 577598
rect 43072 577538 43136 577542
rect 674752 577242 674816 577306
rect 41536 577094 41600 577158
rect 42496 577006 42560 577010
rect 42496 576950 42508 577006
rect 42508 576950 42560 577006
rect 42496 576946 42560 576950
rect 41920 575082 41984 575086
rect 41920 575026 41932 575082
rect 41932 575026 41984 575082
rect 41920 575022 41984 575026
rect 41728 574934 41792 574938
rect 41728 574878 41780 574934
rect 41780 574878 41792 574934
rect 41728 574874 41792 574878
rect 40960 573986 41024 574050
rect 41344 573838 41408 573902
rect 40576 573246 40640 573310
rect 675520 567326 675584 567390
rect 674944 562886 675008 562950
rect 674176 561702 674240 561766
rect 675136 561554 675200 561618
rect 42112 560962 42176 561026
rect 674752 558890 674816 558954
rect 676288 557706 676352 557770
rect 40576 556670 40640 556734
rect 40960 553562 41024 553626
rect 676864 547050 676928 547114
rect 42688 541278 42752 541342
rect 42112 541130 42176 541194
rect 43072 540982 43136 541046
rect 42112 538970 42176 538974
rect 42112 538914 42124 538970
rect 42124 538914 42176 538970
rect 42112 538910 42176 538914
rect 42688 538614 42752 538678
rect 675520 538318 675584 538382
rect 675712 536986 675776 537050
rect 43072 536838 43136 536902
rect 676672 536246 676736 536310
rect 674368 534840 674432 534904
rect 673984 534026 674048 534090
rect 675904 533730 675968 533794
rect 676096 532694 676160 532758
rect 40960 532546 41024 532610
rect 40576 532250 40640 532314
rect 674560 532250 674624 532314
rect 41728 531718 41792 531722
rect 41728 531662 41780 531718
rect 41780 531662 41792 531718
rect 41728 531658 41792 531662
rect 41920 531274 41984 531278
rect 41920 531218 41932 531274
rect 41932 531218 41984 531274
rect 41920 531214 41984 531218
rect 675136 492734 675200 492798
rect 674944 491402 675008 491466
rect 674176 487702 674240 487766
rect 674752 487406 674816 487470
rect 676288 484002 676352 484066
rect 673984 475270 674048 475334
rect 42112 432646 42176 432710
rect 40576 431906 40640 431970
rect 40960 430722 41024 430786
rect 40768 429390 40832 429454
rect 41344 428354 41408 428418
rect 41536 427614 41600 427678
rect 41152 426282 41216 426346
rect 40384 425098 40448 425162
rect 41728 419030 41792 419094
rect 42304 419030 42368 419094
rect 676672 411986 676736 411990
rect 676672 411930 676684 411986
rect 676684 411930 676736 411986
rect 676672 411926 676736 411930
rect 41536 406006 41600 406070
rect 673984 405858 674048 405922
rect 675328 405266 675392 405330
rect 676672 405266 676736 405330
rect 41728 404290 41792 404294
rect 41728 404234 41780 404290
rect 41780 404234 41792 404290
rect 41728 404230 41792 404234
rect 42304 404230 42368 404294
rect 41536 403786 41600 403850
rect 42688 403786 42752 403850
rect 674176 403490 674240 403554
rect 40384 402454 40448 402518
rect 41344 402010 41408 402074
rect 674560 400530 674624 400594
rect 674368 400382 674432 400446
rect 40960 400086 41024 400150
rect 41152 399494 41216 399558
rect 40768 398754 40832 398818
rect 42112 390170 42176 390234
rect 42496 389430 42560 389494
rect 40576 388542 40640 388606
rect 40960 387506 41024 387570
rect 40768 386026 40832 386090
rect 41344 385138 41408 385202
rect 41536 384398 41600 384462
rect 41152 383066 41216 383130
rect 42112 381882 42176 381946
rect 674560 378774 674624 378838
rect 675520 374482 675584 374546
rect 674176 373890 674240 373954
rect 674368 371966 674432 372030
rect 675712 371522 675776 371586
rect 40576 368710 40640 368774
rect 42112 368710 42176 368774
rect 41728 368562 41792 368626
rect 42112 368414 42176 368478
rect 41920 368266 41984 368330
rect 42304 368266 42368 368330
rect 41728 363086 41792 363150
rect 40384 362938 40448 363002
rect 41536 362790 41600 362854
rect 674176 361384 674240 361448
rect 42304 360866 42368 360930
rect 673984 360718 674048 360782
rect 41728 360630 41792 360634
rect 41728 360574 41780 360630
rect 41780 360574 41792 360630
rect 41728 360570 41792 360574
rect 42688 360570 42752 360634
rect 675328 360126 675392 360190
rect 675904 360126 675968 360190
rect 42112 359446 42176 359450
rect 42112 359390 42124 359446
rect 42124 359390 42176 359446
rect 42112 359386 42176 359390
rect 41344 358646 41408 358710
rect 674368 358202 674432 358266
rect 40960 356870 41024 356934
rect 41152 356426 41216 356490
rect 40768 355538 40832 355602
rect 674752 355390 674816 355454
rect 674560 354502 674624 354566
rect 675136 351394 675200 351458
rect 42496 346806 42560 346870
rect 42112 346066 42176 346130
rect 41344 345918 41408 345982
rect 42304 345918 42368 345982
rect 674944 345474 675008 345538
rect 40768 344290 40832 344354
rect 40960 342810 41024 342874
rect 42496 342662 42560 342726
rect 43072 342662 43136 342726
rect 41344 341922 41408 341986
rect 41536 341182 41600 341246
rect 41152 339850 41216 339914
rect 40384 338666 40448 338730
rect 41920 335558 41984 335622
rect 675520 335174 675584 335178
rect 675520 335118 675532 335174
rect 675532 335118 675584 335174
rect 675520 335114 675584 335118
rect 675328 333782 675392 333846
rect 674752 333486 674816 333550
rect 675136 330526 675200 330590
rect 675520 329490 675584 329554
rect 674368 328306 674432 328370
rect 674560 326826 674624 326890
rect 41536 319722 41600 319786
rect 41536 318686 41600 318750
rect 43072 318686 43136 318750
rect 41728 318006 41792 318010
rect 41728 317950 41780 318006
rect 41780 317950 41792 318006
rect 41728 317946 41792 317950
rect 41920 317414 41984 317418
rect 41920 317358 41932 317414
rect 41932 317358 41984 317414
rect 41920 317354 41984 317358
rect 674176 317206 674240 317270
rect 674176 316392 674240 316456
rect 40384 316022 40448 316086
rect 674944 315874 675008 315938
rect 674368 315726 674432 315790
rect 41344 315578 41408 315642
rect 675904 315134 675968 315198
rect 673984 314838 674048 314902
rect 41728 313802 41792 313866
rect 43072 313802 43136 313866
rect 40768 313654 40832 313718
rect 41152 313210 41216 313274
rect 674752 312618 674816 312682
rect 40960 312322 41024 312386
rect 674560 309510 674624 309574
rect 674944 306402 675008 306466
rect 40576 302702 40640 302766
rect 42112 302702 42176 302766
rect 42304 302702 42368 302766
rect 40960 301074 41024 301138
rect 40768 299594 40832 299658
rect 41344 298706 41408 298770
rect 41536 298706 41600 298770
rect 42496 298706 42560 298770
rect 41536 297966 41600 298030
rect 41152 296634 41216 296698
rect 40384 295450 40448 295514
rect 675520 290182 675584 290186
rect 675520 290126 675532 290182
rect 675532 290126 675584 290182
rect 675520 290122 675584 290126
rect 675328 289590 675392 289594
rect 675328 289534 675380 289590
rect 675380 289534 675392 289590
rect 675328 289530 675392 289534
rect 674944 285238 675008 285302
rect 42304 283670 42368 283674
rect 42304 283614 42316 283670
rect 42316 283614 42368 283670
rect 42304 283610 42368 283614
rect 674752 283610 674816 283674
rect 41920 282278 41984 282342
rect 42496 282278 42560 282342
rect 674752 282278 674816 282342
rect 674560 281834 674624 281898
rect 42304 281538 42368 281602
rect 41536 276506 41600 276570
rect 41920 274790 41984 274794
rect 41920 274734 41972 274790
rect 41972 274734 41984 274790
rect 41920 274730 41984 274734
rect 41728 273990 41792 274054
rect 43072 273990 43136 274054
rect 287872 273842 287936 273906
rect 674752 273546 674816 273610
rect 674944 273546 675008 273610
rect 40384 272806 40448 272870
rect 674752 272718 674816 272722
rect 674752 272662 674804 272718
rect 674804 272662 674816 272718
rect 674752 272658 674816 272662
rect 41344 272362 41408 272426
rect 674176 272214 674240 272278
rect 675904 270882 675968 270946
rect 674368 270734 674432 270798
rect 40960 270586 41024 270650
rect 442240 270586 442304 270650
rect 450688 270586 450752 270650
rect 446464 270438 446528 270502
rect 449536 270438 449600 270502
rect 443584 270290 443648 270354
rect 41152 269994 41216 270058
rect 443008 270142 443072 270206
rect 442048 269994 442112 270058
rect 673984 269846 674048 269910
rect 449728 269698 449792 269762
rect 445696 269402 445760 269466
rect 40768 269106 40832 269170
rect 290368 268958 290432 269022
rect 447232 268958 447296 269022
rect 290176 268810 290240 268874
rect 452224 269254 452288 269318
rect 290752 268662 290816 268726
rect 290560 268514 290624 268578
rect 452416 269106 452480 269170
rect 674752 268514 674816 268578
rect 449344 268366 449408 268430
rect 443392 268218 443456 268282
rect 446656 268070 446720 268134
rect 675712 268070 675776 268134
rect 284800 267774 284864 267838
rect 289984 267626 290048 267690
rect 284416 267478 284480 267542
rect 292864 267330 292928 267394
rect 289216 267182 289280 267246
rect 284992 266146 285056 266210
rect 284032 265998 284096 266062
rect 674560 265406 674624 265470
rect 674368 265110 674432 265174
rect 42112 264814 42176 264878
rect 287680 264814 287744 264878
rect 289024 263334 289088 263398
rect 291520 263038 291584 263102
rect 289792 262890 289856 262954
rect 287488 262150 287552 262214
rect 675328 262150 675392 262214
rect 40576 259486 40640 259550
rect 443200 259042 443264 259106
rect 442624 258894 442688 258958
rect 442816 258746 442880 258810
rect 446848 258598 446912 258662
rect 451072 258450 451136 258514
rect 446080 258302 446144 258366
rect 40384 257858 40448 257922
rect 289600 257414 289664 257478
rect 290752 257414 290816 257478
rect 441472 257266 441536 257330
rect 674944 257266 675008 257330
rect 675520 257266 675584 257330
rect 351424 257178 351488 257182
rect 351424 257122 351476 257178
rect 351476 257122 351488 257178
rect 351424 257118 351488 257122
rect 448384 257118 448448 257182
rect 445120 256970 445184 257034
rect 287104 256822 287168 256886
rect 445312 256822 445376 256886
rect 443776 256674 443840 256738
rect 292096 256526 292160 256590
rect 447808 256526 447872 256590
rect 40576 256378 40640 256442
rect 286912 256378 286976 256442
rect 286720 256230 286784 256294
rect 448768 256230 448832 256294
rect 676672 256230 676736 256294
rect 290752 256082 290816 256146
rect 443008 256082 443072 256146
rect 448960 256082 449024 256146
rect 290944 255934 291008 255998
rect 337216 255934 337280 255998
rect 446656 255934 446720 255998
rect 291328 255786 291392 255850
rect 351424 255786 351488 255850
rect 448576 255786 448640 255850
rect 40960 255638 41024 255702
rect 291712 255638 291776 255702
rect 452992 255638 453056 255702
rect 673984 255638 674048 255702
rect 291904 255490 291968 255554
rect 448192 255490 448256 255554
rect 292288 255342 292352 255406
rect 453760 255342 453824 255406
rect 292672 255194 292736 255258
rect 293056 255046 293120 255110
rect 453184 255194 453248 255258
rect 204928 254898 204992 254962
rect 293248 254898 293312 254962
rect 453376 255046 453440 255110
rect 454144 254898 454208 254962
rect 41344 254750 41408 254814
rect 204736 254750 204800 254814
rect 449920 254750 449984 254814
rect 284224 254602 284288 254666
rect 337600 254602 337664 254666
rect 287296 254454 287360 254518
rect 453952 254602 454016 254666
rect 441856 254454 441920 254518
rect 444160 254454 444224 254518
rect 293440 254158 293504 254222
rect 442432 254306 442496 254370
rect 444352 254306 444416 254370
rect 447616 254306 447680 254370
rect 444544 254158 444608 254222
rect 448000 254158 448064 254222
rect 288064 254010 288128 254074
rect 443968 254010 444032 254074
rect 451264 254010 451328 254074
rect 452608 253862 452672 253926
rect 288256 253714 288320 253778
rect 288448 253566 288512 253630
rect 452800 253714 452864 253778
rect 441664 253566 441728 253630
rect 442624 253566 442688 253630
rect 445888 253566 445952 253630
rect 40768 253418 40832 253482
rect 288832 253418 288896 253482
rect 444928 253418 444992 253482
rect 450112 253418 450176 253482
rect 283072 253270 283136 253334
rect 292480 253270 292544 253334
rect 444736 253270 444800 253334
rect 450496 253270 450560 253334
rect 286528 252974 286592 253038
rect 288640 252974 288704 253038
rect 289408 253034 289472 253038
rect 289408 252978 289460 253034
rect 289460 252978 289472 253034
rect 289408 252974 289472 252978
rect 291136 252974 291200 253038
rect 450880 253122 450944 253186
rect 442624 252974 442688 253038
rect 443584 252974 443648 253038
rect 446272 253034 446336 253038
rect 446272 252978 446284 253034
rect 446284 252978 446336 253034
rect 446272 252974 446336 252978
rect 447424 252974 447488 253038
rect 453568 252974 453632 253038
rect 41152 252382 41216 252446
rect 208384 252086 208448 252150
rect 207424 251938 207488 252002
rect 145408 250606 145472 250670
rect 674752 249570 674816 249634
rect 283072 248890 283136 248894
rect 283072 248834 283124 248890
rect 283124 248834 283136 248890
rect 283072 248830 283136 248834
rect 288640 248830 288704 248894
rect 288640 248682 288704 248746
rect 284800 248534 284864 248598
rect 284032 248386 284096 248450
rect 284800 248386 284864 248450
rect 285760 248090 285824 248154
rect 284992 247942 285056 248006
rect 40576 247794 40640 247858
rect 41536 247646 41600 247710
rect 284800 247350 284864 247414
rect 285760 247262 285824 247266
rect 285760 247206 285812 247262
rect 285812 247206 285824 247262
rect 285760 247202 285824 247206
rect 284416 246906 284480 246970
rect 288640 246610 288704 246674
rect 284224 245722 284288 245786
rect 674944 244982 675008 245046
rect 675328 245042 675392 245046
rect 675328 244986 675340 245042
rect 675340 244986 675392 245042
rect 675328 244982 675392 244986
rect 675520 244746 675584 244750
rect 675520 244690 675532 244746
rect 675532 244690 675584 244746
rect 675520 244686 675584 244690
rect 145600 244390 145664 244454
rect 674560 243502 674624 243566
rect 286528 242170 286592 242234
rect 288640 242170 288704 242234
rect 145792 240838 145856 240902
rect 42304 240690 42368 240754
rect 287488 239506 287552 239570
rect 289408 239506 289472 239570
rect 290176 239506 290240 239570
rect 290944 239566 291008 239570
rect 290944 239510 290956 239566
rect 290956 239510 291008 239566
rect 290944 239506 291008 239510
rect 291136 239566 291200 239570
rect 291136 239510 291188 239566
rect 291188 239510 291200 239566
rect 291136 239506 291200 239510
rect 291328 239566 291392 239570
rect 291328 239510 291380 239566
rect 291380 239510 291392 239566
rect 291328 239506 291392 239510
rect 291712 239506 291776 239570
rect 291904 239566 291968 239570
rect 291904 239510 291956 239566
rect 291956 239510 291968 239566
rect 291904 239506 291968 239510
rect 292288 239566 292352 239570
rect 292288 239510 292340 239566
rect 292340 239510 292352 239566
rect 292288 239506 292352 239510
rect 292672 239566 292736 239570
rect 292672 239510 292724 239566
rect 292724 239510 292736 239566
rect 292672 239506 292736 239510
rect 293056 239566 293120 239570
rect 293056 239510 293108 239566
rect 293108 239510 293120 239566
rect 293056 239506 293120 239510
rect 288640 239358 288704 239422
rect 290752 239358 290816 239422
rect 293248 239358 293312 239422
rect 442624 239506 442688 239570
rect 446272 239506 446336 239570
rect 441088 239358 441152 239422
rect 442432 239358 442496 239422
rect 443968 239358 444032 239422
rect 444352 239418 444416 239422
rect 444352 239362 444364 239418
rect 444364 239362 444416 239418
rect 444352 239358 444416 239362
rect 445312 239418 445376 239422
rect 445312 239362 445324 239418
rect 445324 239362 445376 239418
rect 445312 239358 445376 239362
rect 447808 239358 447872 239422
rect 450112 239358 450176 239422
rect 292864 239210 292928 239274
rect 443584 239210 443648 239274
rect 444160 239270 444224 239274
rect 444160 239214 444172 239270
rect 444172 239214 444224 239270
rect 444160 239210 444224 239214
rect 445120 239210 445184 239274
rect 447616 239210 447680 239274
rect 448768 239210 448832 239274
rect 290560 239062 290624 239126
rect 450304 239062 450368 239126
rect 291520 238914 291584 238978
rect 442240 238914 442304 238978
rect 442432 238914 442496 238978
rect 445888 238914 445952 238978
rect 674752 238914 674816 238978
rect 442048 238766 442112 238830
rect 442624 238766 442688 238830
rect 448960 238766 449024 238830
rect 287872 238618 287936 238682
rect 447040 238618 447104 238682
rect 675712 238678 675776 238682
rect 675712 238622 675724 238678
rect 675724 238622 675776 238678
rect 675712 238618 675776 238622
rect 400576 238470 400640 238534
rect 447232 238470 447296 238534
rect 445696 238322 445760 238386
rect 292096 238174 292160 238238
rect 445504 237878 445568 237942
rect 450688 237730 450752 237794
rect 293440 237582 293504 237646
rect 446656 237582 446720 237646
rect 447232 237582 447296 237646
rect 448192 237582 448256 237646
rect 444544 237434 444608 237498
rect 286912 237286 286976 237350
rect 441664 237286 441728 237350
rect 442816 237286 442880 237350
rect 449920 237138 449984 237202
rect 399232 237050 399296 237054
rect 399232 236994 399244 237050
rect 399244 236994 399296 237050
rect 399232 236990 399296 236994
rect 446080 236990 446144 237054
rect 400576 236842 400640 236906
rect 411328 236842 411392 236906
rect 444736 236842 444800 236906
rect 674368 236842 674432 236906
rect 145984 236694 146048 236758
rect 442432 236694 442496 236758
rect 444928 236546 444992 236610
rect 292480 236398 292544 236462
rect 290368 236102 290432 236166
rect 443584 236162 443648 236166
rect 443584 236106 443636 236162
rect 443636 236106 443648 236162
rect 443584 236102 443648 236106
rect 289600 235954 289664 236018
rect 289792 235806 289856 235870
rect 289984 235658 290048 235722
rect 289024 235510 289088 235574
rect 289216 235362 289280 235426
rect 287680 235066 287744 235130
rect 42304 234770 42368 234834
rect 441088 234178 441152 234242
rect 451264 233882 451328 233946
rect 448000 233734 448064 233798
rect 442816 233586 442880 233650
rect 443008 233438 443072 233502
rect 41344 233290 41408 233354
rect 446080 232698 446144 232762
rect 450880 232698 450944 232762
rect 287104 232106 287168 232170
rect 288448 231958 288512 232022
rect 288832 231810 288896 231874
rect 443392 232106 443456 232170
rect 41728 231722 41792 231726
rect 41728 231666 41780 231722
rect 41780 231666 41792 231722
rect 41728 231662 41792 231666
rect 41920 231574 41984 231578
rect 41920 231518 41932 231574
rect 41932 231518 41984 231574
rect 41920 231514 41984 231518
rect 442624 230774 442688 230838
rect 204928 230390 204992 230394
rect 204928 230334 204940 230390
rect 204940 230334 204992 230390
rect 204928 230330 204992 230334
rect 207424 230330 207488 230394
rect 208384 230390 208448 230394
rect 208384 230334 208436 230390
rect 208436 230334 208448 230390
rect 208384 230330 208448 230334
rect 288256 230330 288320 230394
rect 441856 230330 441920 230394
rect 443584 230390 443648 230394
rect 443584 230334 443636 230390
rect 443636 230334 443648 230390
rect 443584 230330 443648 230334
rect 204736 230182 204800 230246
rect 41152 229738 41216 229802
rect 286720 229146 286784 229210
rect 40960 228998 41024 229062
rect 287296 228998 287360 229062
rect 288064 228850 288128 228914
rect 413248 228110 413312 228174
rect 441280 227962 441344 228026
rect 443776 227814 443840 227878
rect 207616 227666 207680 227730
rect 40576 227518 40640 227582
rect 41536 227518 41600 227582
rect 443200 227370 443264 227434
rect 40384 227222 40448 227286
rect 419200 226926 419264 226990
rect 452224 227222 452288 227286
rect 675904 227222 675968 227286
rect 453184 227074 453248 227138
rect 453952 226926 454016 226990
rect 40768 226778 40832 226842
rect 208000 226778 208064 226842
rect 452992 226778 453056 226842
rect 207808 226690 207872 226694
rect 207808 226634 207820 226690
rect 207820 226634 207872 226690
rect 207808 226630 207872 226634
rect 419008 226630 419072 226694
rect 419200 226630 419264 226694
rect 448384 226630 448448 226694
rect 208192 226542 208256 226546
rect 208192 226486 208204 226542
rect 208204 226486 208256 226542
rect 208192 226482 208256 226486
rect 452416 226482 452480 226546
rect 40576 225890 40640 225954
rect 446848 226334 446912 226398
rect 452800 226334 452864 226398
rect 453376 226186 453440 226250
rect 674176 226186 674240 226250
rect 453568 226038 453632 226102
rect 419200 225742 419264 225806
rect 454144 225742 454208 225806
rect 676672 225742 676736 225806
rect 447424 225594 447488 225658
rect 451072 225446 451136 225510
rect 452608 225298 452672 225362
rect 449728 225150 449792 225214
rect 453760 225002 453824 225066
rect 388672 224766 388736 224770
rect 388672 224710 388724 224766
rect 388724 224710 388736 224766
rect 388672 224706 388736 224710
rect 391744 224766 391808 224770
rect 391744 224710 391756 224766
rect 391756 224710 391808 224766
rect 391744 224706 391808 224710
rect 447232 224854 447296 224918
rect 448576 224706 448640 224770
rect 673984 224706 674048 224770
rect 429184 224262 429248 224326
rect 429376 224262 429440 224326
rect 207040 223966 207104 224030
rect 206656 223818 206720 223882
rect 207424 223818 207488 223882
rect 206272 223670 206336 223734
rect 349312 223818 349376 223882
rect 359680 223818 359744 223882
rect 362752 223878 362816 223882
rect 362752 223822 362764 223878
rect 362764 223822 362816 223878
rect 362752 223818 362816 223822
rect 388672 223878 388736 223882
rect 388672 223822 388724 223878
rect 388724 223822 388736 223878
rect 388672 223818 388736 223822
rect 391744 223878 391808 223882
rect 391744 223822 391756 223878
rect 391756 223822 391808 223878
rect 391744 223818 391808 223822
rect 302464 223522 302528 223586
rect 380032 223522 380096 223586
rect 400192 223966 400256 224030
rect 405568 223818 405632 223882
rect 405952 223818 406016 223882
rect 429568 223878 429632 223882
rect 429568 223822 429620 223878
rect 429620 223822 429632 223878
rect 413056 223670 413120 223734
rect 413248 223670 413312 223734
rect 428992 223670 429056 223734
rect 429568 223818 429632 223822
rect 439552 223966 439616 224030
rect 440128 223966 440192 224030
rect 440896 224026 440960 224030
rect 440896 223970 440948 224026
rect 440948 223970 440960 224026
rect 440896 223966 440960 223970
rect 449536 223818 449600 223882
rect 429568 223522 429632 223586
rect 450496 223522 450560 223586
rect 400192 223374 400256 223438
rect 206848 222930 206912 222994
rect 302464 223078 302528 223142
rect 380032 223078 380096 223142
rect 380272 223078 380336 223142
rect 400192 223078 400256 223142
rect 427648 223374 427712 223438
rect 429376 223374 429440 223438
rect 446464 223374 446528 223438
rect 413056 223226 413120 223290
rect 417472 223226 417536 223290
rect 417664 223226 417728 223290
rect 446080 223226 446144 223290
rect 359680 222930 359744 222994
rect 439552 222930 439616 222994
rect 447808 222930 447872 222994
rect 633472 224114 633536 224178
rect 632512 223966 632576 224030
rect 632704 223966 632768 224030
rect 632128 223818 632192 223882
rect 632320 223878 632384 223882
rect 632320 223822 632372 223878
rect 632372 223822 632384 223878
rect 632320 223818 632384 223822
rect 632896 223818 632960 223882
rect 633280 223818 633344 223882
rect 362752 222782 362816 222846
rect 440128 222782 440192 222846
rect 207232 222634 207296 222698
rect 349312 222634 349376 222698
rect 440896 222634 440960 222698
rect 674560 222486 674624 222550
rect 675328 221006 675392 221070
rect 675136 220118 675200 220182
rect 674368 219970 674432 220034
rect 674944 216270 675008 216334
rect 40576 214642 40640 214706
rect 40384 213162 40448 213226
rect 40960 212422 41024 212486
rect 41152 211534 41216 211598
rect 40768 210350 40832 210414
rect 674752 210054 674816 210118
rect 676096 206206 676160 206270
rect 676096 204430 676160 204494
rect 675520 201618 675584 201682
rect 675520 200050 675584 200054
rect 675520 199994 675532 200050
rect 675532 199994 675584 200050
rect 675520 199990 675584 199994
rect 675328 199458 675392 199462
rect 675328 199402 675380 199458
rect 675380 199402 675392 199458
rect 675328 199398 675392 199402
rect 675136 198362 675200 198426
rect 42496 197622 42560 197686
rect 42496 195698 42560 195762
rect 674944 195254 675008 195318
rect 674560 193478 674624 193542
rect 675520 193182 675584 193246
rect 675328 193034 675392 193098
rect 674368 191554 674432 191618
rect 41152 190074 41216 190138
rect 41920 189098 41984 189102
rect 41920 189042 41972 189098
rect 41972 189042 41984 189098
rect 41920 189038 41984 189042
rect 41728 188358 41792 188362
rect 41728 188302 41780 188358
rect 41780 188302 41792 188358
rect 41728 188298 41792 188302
rect 40960 185930 41024 185994
rect 40576 184154 40640 184218
rect 40768 183562 40832 183626
rect 40384 182822 40448 182886
rect 674176 182008 674240 182072
rect 200896 181402 200960 181406
rect 200896 181346 200908 181402
rect 200908 181346 200960 181402
rect 200896 181342 200960 181346
rect 674176 181194 674240 181258
rect 674752 180898 674816 180962
rect 674368 180454 674432 180518
rect 673984 179714 674048 179778
rect 674752 177494 674816 177558
rect 31744 177050 31808 177114
rect 674560 174386 674624 174450
rect 674944 171278 675008 171342
rect 200896 166898 200960 166902
rect 200896 166842 200948 166898
rect 200948 166842 200960 166898
rect 200896 166838 200960 166842
rect 675712 161362 675776 161426
rect 675328 155206 675392 155210
rect 675328 155150 675340 155206
rect 675340 155150 675392 155206
rect 675328 155146 675392 155150
rect 675520 155058 675584 155062
rect 675520 155002 675532 155058
rect 675532 155002 675584 155058
rect 675520 154998 675584 155002
rect 675712 153430 675776 153434
rect 675712 153374 675764 153430
rect 675764 153374 675776 153430
rect 675712 153370 675776 153374
rect 674944 150262 675008 150326
rect 674752 148486 674816 148550
rect 674560 146414 674624 146478
rect 674368 142774 674432 142778
rect 674368 142718 674380 142774
rect 674380 142718 674432 142774
rect 674368 142714 674432 142718
rect 674176 136794 674240 136858
rect 673984 135018 674048 135082
rect 674560 132502 674624 132566
rect 674368 130578 674432 130642
rect 674176 129690 674240 129754
rect 675136 126730 675200 126794
rect 31744 125250 31808 125314
rect 675136 110746 675200 110810
rect 675520 110066 675584 110070
rect 675520 110010 675572 110066
rect 675572 110010 675584 110066
rect 675520 110006 675584 110010
rect 674368 108082 674432 108146
rect 674560 103198 674624 103262
rect 674176 101422 674240 101486
rect 204352 86622 204416 86686
rect 204160 62202 204224 62266
rect 204736 58858 204800 58862
rect 204736 58802 204748 58858
rect 204748 58802 204800 58858
rect 204736 58798 204800 58802
rect 204928 56726 204992 56790
rect 206080 54654 206144 54718
rect 206272 54358 206336 54422
rect 207424 54210 207488 54274
rect 208000 54062 208064 54126
rect 207616 53914 207680 53978
rect 204736 53766 204800 53830
rect 206656 53618 206720 53682
rect 207232 53470 207296 53534
rect 207808 53470 207872 53534
rect 207040 53322 207104 53386
rect 204928 53174 204992 53238
rect 471040 53174 471104 53238
rect 204160 52434 204224 52498
rect 208192 52286 208256 52350
rect 632704 52138 632768 52202
rect 632896 51990 632960 52054
rect 204352 51842 204416 51906
rect 633280 51842 633344 51906
rect 632512 51694 632576 51758
rect 145600 51250 145664 51314
rect 145984 51102 146048 51166
rect 145792 50954 145856 51018
rect 145408 50806 145472 50870
rect 632320 50362 632384 50426
rect 632128 48882 632192 48946
rect 633472 48734 633536 48798
rect 302464 45478 302528 45542
rect 305344 45330 305408 45394
rect 356992 45182 357056 45246
rect 360064 45034 360128 45098
rect 362944 44886 363008 44950
rect 302464 43318 302528 43322
rect 302464 43262 302516 43318
rect 302516 43262 302528 43318
rect 302464 43258 302528 43262
rect 305344 43258 305408 43322
rect 360064 43258 360128 43322
rect 362944 43258 363008 43322
rect 356992 43110 357056 43174
rect 471040 42134 471104 42138
rect 471040 42078 471092 42134
rect 471092 42078 471104 42134
rect 471040 42074 471104 42078
rect 189952 41778 190016 41842
rect 194944 41778 195008 41842
rect 518464 41838 518528 41842
rect 518464 41782 518516 41838
rect 518516 41782 518528 41838
rect 518464 41778 518528 41782
rect 189952 40742 190016 40806
rect 518272 40742 518336 40806
rect 194944 40594 195008 40658
<< metal4 >>
rect 385983 996146 386049 996147
rect 385983 996082 385984 996146
rect 386048 996082 386049 996146
rect 385983 996081 386049 996082
rect 385986 995555 386046 996081
rect 385983 995554 386049 995555
rect 385983 995490 385984 995554
rect 386048 995490 386049 995554
rect 385983 995489 386049 995490
rect 294783 993630 294849 993631
rect 294783 993566 294784 993630
rect 294848 993566 294849 993630
rect 294783 993565 294849 993566
rect 294786 992151 294846 993565
rect 294783 992150 294849 992151
rect 294783 992086 294784 992150
rect 294848 992086 294849 992150
rect 294783 992085 294849 992086
rect 40575 968766 40641 968767
rect 40575 968702 40576 968766
rect 40640 968702 40641 968766
rect 40575 968701 40641 968702
rect 40383 965066 40449 965067
rect 40383 965002 40384 965066
rect 40448 965002 40449 965066
rect 40383 965001 40449 965002
rect 40386 895655 40446 965001
rect 40578 899207 40638 968701
rect 675519 967582 675585 967583
rect 675519 967518 675520 967582
rect 675584 967518 675585 967582
rect 675519 967517 675585 967518
rect 41727 967138 41793 967139
rect 41727 967074 41728 967138
rect 41792 967074 41793 967138
rect 41727 967073 41793 967074
rect 40767 964030 40833 964031
rect 40767 963966 40768 964030
rect 40832 963966 40833 964030
rect 40767 963965 40833 963966
rect 40575 899206 40641 899207
rect 40575 899142 40576 899206
rect 40640 899142 40641 899206
rect 40575 899141 40641 899142
rect 40383 895654 40449 895655
rect 40383 895590 40384 895654
rect 40448 895590 40449 895654
rect 40383 895589 40449 895590
rect 40770 892547 40830 963965
rect 40959 963438 41025 963439
rect 40959 963374 40960 963438
rect 41024 963374 41025 963438
rect 40959 963373 41025 963374
rect 40962 895063 41022 963373
rect 41151 962846 41217 962847
rect 41151 962782 41152 962846
rect 41216 962782 41217 962846
rect 41151 962781 41217 962782
rect 40959 895062 41025 895063
rect 40959 894998 40960 895062
rect 41024 894998 41025 895062
rect 40959 894997 41025 894998
rect 41154 893583 41214 962781
rect 41535 962254 41601 962255
rect 41535 962190 41536 962254
rect 41600 962190 41601 962254
rect 41535 962189 41601 962190
rect 41343 959738 41409 959739
rect 41343 959674 41344 959738
rect 41408 959674 41409 959738
rect 41343 959673 41409 959674
rect 41346 894471 41406 959673
rect 41538 899799 41598 962189
rect 41730 902315 41790 967073
rect 674559 965658 674625 965659
rect 674559 965594 674560 965658
rect 674624 965594 674625 965658
rect 674559 965593 674625 965594
rect 674367 962550 674433 962551
rect 674367 962486 674368 962550
rect 674432 962486 674433 962550
rect 674367 962485 674433 962486
rect 42879 962254 42945 962255
rect 42879 962190 42880 962254
rect 42944 962190 42945 962254
rect 42879 962189 42945 962190
rect 41919 959146 41985 959147
rect 41919 959082 41920 959146
rect 41984 959082 41985 959146
rect 41919 959081 41985 959082
rect 41727 902314 41793 902315
rect 41727 902250 41728 902314
rect 41792 902250 41793 902314
rect 41727 902249 41793 902250
rect 41535 899798 41601 899799
rect 41535 899734 41536 899798
rect 41600 899734 41601 899798
rect 41535 899733 41601 899734
rect 41922 896691 41982 959081
rect 42111 958406 42177 958407
rect 42111 958342 42112 958406
rect 42176 958342 42177 958406
rect 42111 958341 42177 958342
rect 42114 897579 42174 958341
rect 42303 957814 42369 957815
rect 42303 957750 42304 957814
rect 42368 957750 42369 957814
rect 42303 957749 42369 957750
rect 42306 900687 42366 957749
rect 42495 956186 42561 956187
rect 42495 956122 42496 956186
rect 42560 956122 42561 956186
rect 42495 956121 42561 956122
rect 42498 903055 42558 956121
rect 42882 907199 42942 962189
rect 43071 962106 43137 962107
rect 43071 962042 43072 962106
rect 43136 962042 43137 962106
rect 43071 962041 43137 962042
rect 42879 907198 42945 907199
rect 42879 907134 42880 907198
rect 42944 907134 42945 907198
rect 42879 907133 42945 907134
rect 42687 903350 42753 903351
rect 42687 903286 42688 903350
rect 42752 903286 42753 903350
rect 42687 903285 42753 903286
rect 42495 903054 42561 903055
rect 42495 902990 42496 903054
rect 42560 902990 42561 903054
rect 42495 902989 42561 902990
rect 42303 900686 42369 900687
rect 42303 900622 42304 900686
rect 42368 900622 42369 900686
rect 42303 900621 42369 900622
rect 42111 897578 42177 897579
rect 42111 897514 42112 897578
rect 42176 897514 42177 897578
rect 42111 897513 42177 897514
rect 41919 896690 41985 896691
rect 41919 896626 41920 896690
rect 41984 896626 41985 896690
rect 41919 896625 41985 896626
rect 41343 894470 41409 894471
rect 41343 894406 41344 894470
rect 41408 894406 41409 894470
rect 41343 894405 41409 894406
rect 41151 893582 41217 893583
rect 41151 893518 41152 893582
rect 41216 893518 41217 893582
rect 41151 893517 41217 893518
rect 40767 892546 40833 892547
rect 40767 892482 40768 892546
rect 40832 892482 40833 892546
rect 40767 892481 40833 892482
rect 42690 884145 42750 903285
rect 42879 887218 42945 887219
rect 42879 887154 42880 887218
rect 42944 887154 42945 887218
rect 42879 887153 42945 887154
rect 42498 884085 42750 884145
rect 42498 874155 42558 884085
rect 42498 874095 42750 874155
rect 42303 866498 42369 866499
rect 42303 866434 42304 866498
rect 42368 866434 42369 866498
rect 42303 866433 42369 866434
rect 42306 864165 42366 866433
rect 42690 864279 42750 874095
rect 42882 866499 42942 887153
rect 42879 866498 42945 866499
rect 42879 866434 42880 866498
rect 42944 866434 42945 866498
rect 42879 866433 42945 866434
rect 42687 864278 42753 864279
rect 42687 864214 42688 864278
rect 42752 864214 42753 864278
rect 42687 864213 42753 864214
rect 42306 864105 42558 864165
rect 42498 858211 42558 864105
rect 42687 864130 42753 864131
rect 42687 864066 42688 864130
rect 42752 864066 42753 864130
rect 42687 864065 42753 864066
rect 42495 858210 42561 858211
rect 42495 858146 42496 858210
rect 42560 858146 42561 858210
rect 42495 858145 42561 858146
rect 42690 852735 42750 864065
rect 42687 852734 42753 852735
rect 42687 852670 42688 852734
rect 42752 852670 42753 852734
rect 42687 852669 42753 852670
rect 39999 842670 40065 842671
rect 39999 842606 40000 842670
rect 40064 842606 40065 842670
rect 39999 842605 40065 842606
rect 40002 827575 40062 842605
rect 43074 841043 43134 962041
rect 674370 934727 674430 962485
rect 674562 938871 674622 965593
rect 674751 964918 674817 964919
rect 674751 964854 674752 964918
rect 674816 964854 674817 964918
rect 674751 964853 674817 964854
rect 674754 940943 674814 964853
rect 674943 962846 675009 962847
rect 674943 962782 674944 962846
rect 675008 962782 675009 962846
rect 674943 962781 675009 962782
rect 674751 940942 674817 940943
rect 674751 940878 674752 940942
rect 674816 940878 674817 940942
rect 674751 940877 674817 940878
rect 674559 938870 674625 938871
rect 674559 938806 674560 938870
rect 674624 938806 674625 938870
rect 674559 938805 674625 938806
rect 674946 938427 675006 962781
rect 675327 962254 675393 962255
rect 675327 962190 675328 962254
rect 675392 962190 675393 962254
rect 675327 962189 675393 962190
rect 675135 956038 675201 956039
rect 675135 955974 675136 956038
rect 675200 955974 675201 956038
rect 675135 955973 675201 955974
rect 674943 938426 675009 938427
rect 674943 938362 674944 938426
rect 675008 938362 675009 938426
rect 674943 938361 675009 938362
rect 674367 934726 674433 934727
rect 674367 934662 674368 934726
rect 674432 934662 674433 934726
rect 674367 934661 674433 934662
rect 675138 933691 675198 955973
rect 675330 934579 675390 962189
rect 675522 961071 675582 967517
rect 675903 965658 675969 965659
rect 675903 965594 675904 965658
rect 675968 965594 675969 965658
rect 675903 965593 675969 965594
rect 675519 961070 675585 961071
rect 675519 961006 675520 961070
rect 675584 961006 675585 961070
rect 675519 961005 675585 961006
rect 675327 934578 675393 934579
rect 675327 934514 675328 934578
rect 675392 934514 675393 934578
rect 675327 934513 675393 934514
rect 675135 933690 675201 933691
rect 675135 933626 675136 933690
rect 675200 933626 675201 933690
rect 675135 933625 675201 933626
rect 674367 876414 674433 876415
rect 674367 876350 674368 876414
rect 674432 876350 674433 876414
rect 674367 876349 674433 876350
rect 674175 872862 674241 872863
rect 674175 872798 674176 872862
rect 674240 872798 674241 872862
rect 674175 872797 674241 872798
rect 43263 858062 43329 858063
rect 43263 857998 43264 858062
rect 43328 857998 43329 858062
rect 43263 857997 43329 857998
rect 43071 841042 43137 841043
rect 43071 840978 43072 841042
rect 43136 840978 43137 841042
rect 43071 840977 43137 840978
rect 43071 840746 43137 840747
rect 43071 840682 43072 840746
rect 43136 840682 43137 840746
rect 43071 840681 43137 840682
rect 42879 830978 42945 830979
rect 42879 830914 42880 830978
rect 42944 830914 42945 830978
rect 42879 830913 42945 830914
rect 39999 827574 40065 827575
rect 39999 827510 40000 827574
rect 40064 827510 40065 827574
rect 39999 827509 40065 827510
rect 40767 818398 40833 818399
rect 40767 818334 40768 818398
rect 40832 818334 40833 818398
rect 40767 818333 40833 818334
rect 40770 775183 40830 818333
rect 42882 804225 42942 830913
rect 42690 804165 42942 804225
rect 42690 803559 42750 804165
rect 42498 803499 42750 803559
rect 41343 802118 41409 802119
rect 41343 802054 41344 802118
rect 41408 802054 41409 802118
rect 41343 802053 41409 802054
rect 41346 791759 41406 802053
rect 41535 801970 41601 801971
rect 41535 801906 41536 801970
rect 41600 801906 41601 801970
rect 41535 801905 41601 801906
rect 41538 791907 41598 801905
rect 41727 800342 41793 800343
rect 41727 800278 41728 800342
rect 41792 800278 41793 800342
rect 41727 800277 41793 800278
rect 42111 800342 42177 800343
rect 42111 800278 42112 800342
rect 42176 800278 42177 800342
rect 42111 800277 42177 800278
rect 41730 794275 41790 800277
rect 41727 794274 41793 794275
rect 41727 794210 41728 794274
rect 41792 794210 41793 794274
rect 41727 794209 41793 794210
rect 41727 794126 41793 794127
rect 41727 794062 41728 794126
rect 41792 794062 41793 794126
rect 41727 794061 41793 794062
rect 41535 791906 41601 791907
rect 41535 791842 41536 791906
rect 41600 791842 41601 791906
rect 41535 791841 41601 791842
rect 41343 791758 41409 791759
rect 41343 791694 41344 791758
rect 41408 791694 41409 791758
rect 41343 791693 41409 791694
rect 41730 791167 41790 794061
rect 42114 792203 42174 800277
rect 42303 800046 42369 800047
rect 42303 799982 42304 800046
rect 42368 799982 42369 800046
rect 42303 799981 42369 799982
rect 42306 797975 42366 799981
rect 42303 797974 42369 797975
rect 42303 797910 42304 797974
rect 42368 797910 42369 797974
rect 42303 797909 42369 797910
rect 42111 792202 42177 792203
rect 42111 792138 42112 792202
rect 42176 792138 42177 792202
rect 42111 792137 42177 792138
rect 41727 791166 41793 791167
rect 41727 791102 41728 791166
rect 41792 791102 41793 791166
rect 41727 791101 41793 791102
rect 40767 775182 40833 775183
rect 40767 775118 40768 775182
rect 40832 775118 40833 775182
rect 40767 775117 40833 775118
rect 40383 759642 40449 759643
rect 40383 759578 40384 759642
rect 40448 759578 40449 759642
rect 40383 759577 40449 759578
rect 40386 747211 40446 759577
rect 40383 747210 40449 747211
rect 40383 747146 40384 747210
rect 40448 747146 40449 747210
rect 40383 747145 40449 747146
rect 40770 733151 40830 775117
rect 40959 760234 41025 760235
rect 40959 760170 40960 760234
rect 41024 760170 41025 760234
rect 40959 760169 41025 760170
rect 40962 746915 41022 760169
rect 41151 758606 41217 758607
rect 41151 758542 41152 758606
rect 41216 758542 41217 758606
rect 41151 758541 41217 758542
rect 41154 754907 41214 758541
rect 41151 754906 41217 754907
rect 41151 754842 41152 754906
rect 41216 754842 41217 754906
rect 41151 754841 41217 754842
rect 41730 748947 41790 791101
rect 42498 791019 42558 803499
rect 42687 800490 42753 800491
rect 42687 800426 42688 800490
rect 42752 800426 42753 800490
rect 42687 800425 42753 800426
rect 42690 794867 42750 800425
rect 42687 794866 42753 794867
rect 42687 794802 42688 794866
rect 42752 794802 42753 794866
rect 42687 794801 42753 794802
rect 43074 794127 43134 840681
rect 43266 830979 43326 857997
rect 43263 830978 43329 830979
rect 43263 830914 43264 830978
rect 43328 830914 43329 830978
rect 43263 830913 43329 830914
rect 43071 794126 43137 794127
rect 43071 794062 43072 794126
rect 43136 794062 43137 794126
rect 43071 794061 43137 794062
rect 41919 791018 41985 791019
rect 41919 790954 41920 791018
rect 41984 790954 41985 791018
rect 41919 790953 41985 790954
rect 42495 791018 42561 791019
rect 42495 790954 42496 791018
rect 42560 790954 42561 791018
rect 42495 790953 42561 790954
rect 41922 762267 41982 790953
rect 673983 787466 674049 787467
rect 673983 787402 673984 787466
rect 674048 787402 674049 787466
rect 673983 787401 674049 787402
rect 42303 763194 42369 763195
rect 42303 763130 42304 763194
rect 42368 763130 42369 763194
rect 42303 763129 42369 763130
rect 42306 762751 42366 763129
rect 42303 762750 42369 762751
rect 42303 762686 42304 762750
rect 42368 762686 42369 762750
rect 42303 762685 42369 762686
rect 41922 762207 42558 762267
rect 42111 761862 42177 761863
rect 42111 761798 42112 761862
rect 42176 761798 42177 761862
rect 42111 761797 42177 761798
rect 41538 748887 41790 748947
rect 40959 746914 41025 746915
rect 40959 746850 40960 746914
rect 41024 746850 41025 746914
rect 40959 746849 41025 746850
rect 40575 733150 40641 733151
rect 40575 733086 40576 733150
rect 40640 733086 40641 733150
rect 40575 733085 40641 733086
rect 40767 733150 40833 733151
rect 40767 733086 40768 733150
rect 40832 733086 40833 733150
rect 40767 733085 40833 733086
rect 40578 689639 40638 733085
rect 41151 732262 41217 732263
rect 41151 732198 41152 732262
rect 41216 732198 41217 732262
rect 41151 732197 41217 732198
rect 40959 726342 41025 726343
rect 40959 726278 40960 726342
rect 41024 726278 41025 726342
rect 40959 726277 41025 726278
rect 40962 703551 41022 726277
rect 40959 703550 41025 703551
rect 40959 703486 40960 703550
rect 41024 703486 41025 703550
rect 40959 703485 41025 703486
rect 41154 689639 41214 732197
rect 41343 729598 41409 729599
rect 41343 729534 41344 729598
rect 41408 729534 41409 729598
rect 41343 729533 41409 729534
rect 41346 703699 41406 729533
rect 41538 711395 41598 748887
rect 41730 748691 41790 748887
rect 41727 748690 41793 748691
rect 41727 748626 41728 748690
rect 41792 748626 41793 748690
rect 41727 748625 41793 748626
rect 42114 748281 42174 761797
rect 42303 757126 42369 757127
rect 42303 757062 42304 757126
rect 42368 757062 42369 757126
rect 42303 757061 42369 757062
rect 42306 754315 42366 757061
rect 42303 754314 42369 754315
rect 42303 754250 42304 754314
rect 42368 754250 42369 754314
rect 42303 754249 42369 754250
rect 41730 748221 42174 748281
rect 41730 733891 41790 748221
rect 42498 747615 42558 762207
rect 42687 751946 42753 751947
rect 42687 751882 42688 751946
rect 42752 751882 42753 751946
rect 42687 751881 42753 751882
rect 42690 751651 42750 751881
rect 42687 751650 42753 751651
rect 42687 751586 42688 751650
rect 42752 751586 42753 751650
rect 42687 751585 42753 751586
rect 41922 747555 42558 747615
rect 41922 747359 41982 747555
rect 41919 747358 41985 747359
rect 41919 747294 41920 747358
rect 41984 747294 41985 747358
rect 41919 747293 41985 747294
rect 41727 733890 41793 733891
rect 41727 733826 41728 733890
rect 41792 733826 41793 733890
rect 41727 733825 41793 733826
rect 41727 716130 41793 716131
rect 41727 716066 41728 716130
rect 41792 716066 41793 716130
rect 41727 716065 41793 716066
rect 41730 711651 41790 716065
rect 41730 711591 41838 711651
rect 41535 711394 41601 711395
rect 41535 711330 41536 711394
rect 41600 711330 41601 711394
rect 41535 711329 41601 711330
rect 41778 711244 41838 711591
rect 41922 711392 41982 747293
rect 42495 721606 42561 721607
rect 42495 721542 42496 721606
rect 42560 721542 42561 721606
rect 42495 721541 42561 721542
rect 42111 714058 42177 714059
rect 42111 713994 42112 714058
rect 42176 713994 42177 714058
rect 42111 713993 42177 713994
rect 42114 711691 42174 713993
rect 42303 713910 42369 713911
rect 42303 713846 42304 713910
rect 42368 713846 42369 713910
rect 42303 713845 42369 713846
rect 42111 711690 42177 711691
rect 42111 711626 42112 711690
rect 42176 711626 42177 711690
rect 42111 711625 42177 711626
rect 41922 711332 42222 711392
rect 42162 711244 42222 711332
rect 41778 711184 41982 711244
rect 41727 711098 41793 711099
rect 41727 711034 41728 711098
rect 41792 711034 41793 711098
rect 41727 711033 41793 711034
rect 41730 705031 41790 711033
rect 41922 706511 41982 711184
rect 42114 711184 42222 711244
rect 41919 706510 41985 706511
rect 41919 706446 41920 706510
rect 41984 706446 41985 706510
rect 41919 706445 41985 706446
rect 41727 705030 41793 705031
rect 41727 704966 41728 705030
rect 41792 704966 41793 705030
rect 41727 704965 41793 704966
rect 41535 704734 41601 704735
rect 41535 704670 41536 704734
rect 41600 704670 41601 704734
rect 41535 704669 41601 704670
rect 41343 703698 41409 703699
rect 41343 703634 41344 703698
rect 41408 703634 41409 703698
rect 41343 703633 41409 703634
rect 41538 692747 41598 704669
rect 42114 704143 42174 711184
rect 42306 711099 42366 713845
rect 42303 711098 42369 711099
rect 42303 711034 42304 711098
rect 42368 711034 42369 711098
rect 42303 711033 42369 711034
rect 42498 707399 42558 721541
rect 43071 721458 43137 721459
rect 43071 721394 43072 721458
rect 43136 721394 43137 721458
rect 43071 721393 43137 721394
rect 42879 711838 42945 711839
rect 42879 711774 42880 711838
rect 42944 711774 42945 711838
rect 42879 711773 42945 711774
rect 42687 711690 42753 711691
rect 42687 711626 42688 711690
rect 42752 711626 42753 711690
rect 42687 711625 42753 711626
rect 42690 711247 42750 711625
rect 42687 711246 42753 711247
rect 42687 711182 42688 711246
rect 42752 711182 42753 711246
rect 42687 711181 42753 711182
rect 42882 707843 42942 711773
rect 43074 708583 43134 721393
rect 673986 712135 674046 787401
rect 674178 755499 674238 872797
rect 674370 760309 674430 876349
rect 674751 876266 674817 876267
rect 674751 876202 674752 876266
rect 674816 876202 674817 876266
rect 674751 876201 674817 876202
rect 674559 873454 674625 873455
rect 674559 873390 674560 873454
rect 674624 873390 674625 873454
rect 674559 873389 674625 873390
rect 674367 760308 674433 760309
rect 674367 760244 674368 760308
rect 674432 760244 674433 760308
rect 674367 760243 674433 760244
rect 674562 756979 674622 873389
rect 674754 762455 674814 876201
rect 674943 874046 675009 874047
rect 674943 873982 674944 874046
rect 675008 873982 675009 874046
rect 674943 873981 675009 873982
rect 674751 762454 674817 762455
rect 674751 762390 674752 762454
rect 674816 762390 674817 762454
rect 674751 762389 674817 762390
rect 674946 760087 675006 873981
rect 675522 872419 675582 961005
rect 675711 960182 675777 960183
rect 675711 960118 675712 960182
rect 675776 960118 675777 960182
rect 675711 960117 675777 960118
rect 675714 875823 675774 960117
rect 675906 935911 675966 965593
rect 676671 961514 676737 961515
rect 676671 961450 676672 961514
rect 676736 961450 676737 961514
rect 676671 961449 676737 961450
rect 676479 957666 676545 957667
rect 676479 957602 676480 957666
rect 676544 957602 676545 957666
rect 676479 957601 676545 957602
rect 675903 935910 675969 935911
rect 675903 935846 675904 935910
rect 675968 935846 675969 935910
rect 675903 935845 675969 935846
rect 676482 932655 676542 957601
rect 676479 932654 676545 932655
rect 676479 932590 676480 932654
rect 676544 932590 676545 932654
rect 676479 932589 676545 932590
rect 676674 931915 676734 961449
rect 677055 953522 677121 953523
rect 677055 953458 677056 953522
rect 677120 953458 677121 953522
rect 677055 953457 677121 953458
rect 676863 953374 676929 953375
rect 676863 953310 676864 953374
rect 676928 953310 676929 953374
rect 676863 953309 676929 953310
rect 676671 931914 676737 931915
rect 676671 931850 676672 931914
rect 676736 931850 676737 931914
rect 676671 931849 676737 931850
rect 676866 930287 676926 953309
rect 677058 931471 677118 953457
rect 677055 931470 677121 931471
rect 677055 931406 677056 931470
rect 677120 931406 677121 931470
rect 677055 931405 677121 931406
rect 676863 930286 676929 930287
rect 676863 930222 676864 930286
rect 676928 930222 676929 930286
rect 676863 930221 676929 930222
rect 676671 876414 676737 876415
rect 676671 876350 676672 876414
rect 676736 876350 676737 876414
rect 676671 876349 676737 876350
rect 675711 875822 675777 875823
rect 675711 875758 675712 875822
rect 675776 875758 675777 875822
rect 675711 875757 675777 875758
rect 675519 872418 675585 872419
rect 675519 872354 675520 872418
rect 675584 872354 675585 872418
rect 675519 872353 675585 872354
rect 675327 869902 675393 869903
rect 675327 869838 675328 869902
rect 675392 869838 675393 869902
rect 675327 869837 675393 869838
rect 675135 866942 675201 866943
rect 675135 866878 675136 866942
rect 675200 866878 675201 866942
rect 675135 866877 675201 866878
rect 674943 760086 675009 760087
rect 674943 760022 674944 760086
rect 675008 760022 675009 760086
rect 674943 760021 675009 760022
rect 674559 756978 674625 756979
rect 674559 756914 674560 756978
rect 674624 756914 674625 756978
rect 674559 756913 674625 756914
rect 674175 755498 674241 755499
rect 674175 755434 674176 755498
rect 674240 755434 674241 755498
rect 674175 755433 674241 755434
rect 675138 755351 675198 866877
rect 675330 759199 675390 869837
rect 675519 864722 675585 864723
rect 675519 864658 675520 864722
rect 675584 864658 675585 864722
rect 675519 864657 675585 864658
rect 675522 761715 675582 864657
rect 675711 862946 675777 862947
rect 675711 862882 675712 862946
rect 675776 862882 675777 862946
rect 675711 862881 675777 862882
rect 675519 761714 675585 761715
rect 675519 761650 675520 761714
rect 675584 761650 675585 761714
rect 675519 761649 675585 761650
rect 675327 759198 675393 759199
rect 675327 759134 675328 759198
rect 675392 759134 675393 759198
rect 675327 759133 675393 759134
rect 675714 758607 675774 862881
rect 676287 787910 676353 787911
rect 676287 787846 676288 787910
rect 676352 787846 676353 787910
rect 676287 787845 676353 787846
rect 675903 786726 675969 786727
rect 675903 786662 675904 786726
rect 675968 786662 675969 786726
rect 675903 786661 675969 786662
rect 675711 758606 675777 758607
rect 675711 758542 675712 758606
rect 675776 758542 675777 758606
rect 675711 758541 675777 758542
rect 675135 755350 675201 755351
rect 675135 755286 675136 755350
rect 675200 755286 675201 755350
rect 675135 755285 675201 755286
rect 674367 743362 674433 743363
rect 674367 743298 674368 743362
rect 674432 743298 674433 743362
rect 674367 743297 674433 743298
rect 674175 741438 674241 741439
rect 674175 741374 674176 741438
rect 674240 741374 674241 741438
rect 674175 741373 674241 741374
rect 673983 712134 674049 712135
rect 673983 712070 673984 712134
rect 674048 712070 674049 712134
rect 673983 712069 674049 712070
rect 43071 708582 43137 708583
rect 43071 708518 43072 708582
rect 43136 708518 43137 708582
rect 43071 708517 43137 708518
rect 42879 707842 42945 707843
rect 42879 707778 42880 707842
rect 42944 707778 42945 707842
rect 42879 707777 42945 707778
rect 42495 707398 42561 707399
rect 42495 707334 42496 707398
rect 42560 707334 42561 707398
rect 42495 707333 42561 707334
rect 42111 704142 42177 704143
rect 42111 704078 42112 704142
rect 42176 704078 42177 704142
rect 42111 704077 42177 704078
rect 41535 692746 41601 692747
rect 41535 692682 41536 692746
rect 41600 692682 41601 692746
rect 41535 692681 41601 692682
rect 42114 691671 42174 704077
rect 673983 697334 674049 697335
rect 673983 697270 673984 697334
rect 674048 697270 674049 697334
rect 673983 697269 674049 697270
rect 41346 691611 42174 691671
rect 40575 689638 40641 689639
rect 40575 689574 40576 689638
rect 40640 689574 40641 689638
rect 40575 689573 40641 689574
rect 41151 689638 41217 689639
rect 41151 689574 41152 689638
rect 41216 689574 41217 689638
rect 41151 689573 41217 689574
rect 40578 646423 40638 689573
rect 41151 686382 41217 686383
rect 41151 686318 41152 686382
rect 41216 686318 41217 686382
rect 41151 686317 41217 686318
rect 40959 683274 41025 683275
rect 40959 683210 40960 683274
rect 41024 683210 41025 683274
rect 40959 683209 41025 683210
rect 40962 660927 41022 683209
rect 40959 660926 41025 660927
rect 40959 660862 40960 660926
rect 41024 660862 41025 660926
rect 40959 660861 41025 660862
rect 41154 656191 41214 686317
rect 41346 675021 41406 691611
rect 42111 688750 42177 688751
rect 42111 688686 42112 688750
rect 42176 688686 42177 688750
rect 42111 688685 42177 688686
rect 41346 674961 41598 675021
rect 41343 674838 41409 674839
rect 41343 674774 41344 674838
rect 41408 674774 41409 674838
rect 41343 674773 41409 674774
rect 41346 665811 41406 674773
rect 41343 665810 41409 665811
rect 41343 665746 41344 665810
rect 41408 665746 41409 665810
rect 41343 665745 41409 665746
rect 41343 665662 41409 665663
rect 41343 665598 41344 665662
rect 41408 665598 41409 665662
rect 41343 665597 41409 665598
rect 41346 661371 41406 665597
rect 41538 661701 41598 674961
rect 41727 670990 41793 670991
rect 41727 670926 41728 670990
rect 41792 670926 41793 670990
rect 41727 670925 41793 670926
rect 41730 668475 41790 670925
rect 41727 668474 41793 668475
rect 41727 668410 41728 668474
rect 41792 668410 41793 668474
rect 41727 668409 41793 668410
rect 41538 661641 41982 661701
rect 41343 661370 41409 661371
rect 41343 661306 41344 661370
rect 41408 661306 41409 661370
rect 41343 661305 41409 661306
rect 41727 661370 41793 661371
rect 41727 661306 41728 661370
rect 41792 661306 41793 661370
rect 41727 661305 41793 661306
rect 41151 656190 41217 656191
rect 41151 656126 41152 656190
rect 41216 656126 41217 656190
rect 41151 656125 41217 656126
rect 40575 646422 40641 646423
rect 40575 646358 40576 646422
rect 40640 646358 40641 646422
rect 40575 646357 40641 646358
rect 40578 603947 40638 646357
rect 40767 643166 40833 643167
rect 40767 643102 40768 643166
rect 40832 643102 40833 643166
rect 40767 643101 40833 643102
rect 40770 618155 40830 643101
rect 40959 640058 41025 640059
rect 40959 639994 40960 640058
rect 41024 639994 41025 640058
rect 40959 639993 41025 639994
rect 40767 618154 40833 618155
rect 40767 618090 40768 618154
rect 40832 618090 40833 618154
rect 40767 618089 40833 618090
rect 40962 617711 41022 639993
rect 41535 635174 41601 635175
rect 41535 635110 41536 635174
rect 41600 635110 41601 635174
rect 41535 635109 41601 635110
rect 41343 627774 41409 627775
rect 41343 627710 41344 627774
rect 41408 627710 41409 627774
rect 41343 627709 41409 627710
rect 41346 625259 41406 627709
rect 41343 625258 41409 625259
rect 41343 625194 41344 625258
rect 41408 625194 41409 625258
rect 41343 625193 41409 625194
rect 41538 624371 41598 635109
rect 41535 624370 41601 624371
rect 41535 624306 41536 624370
rect 41600 624306 41601 624370
rect 41535 624305 41601 624306
rect 41730 619191 41790 661305
rect 41922 661075 41982 661641
rect 41919 661074 41985 661075
rect 41919 661010 41920 661074
rect 41984 661010 41985 661074
rect 41919 661009 41985 661010
rect 41727 619190 41793 619191
rect 41727 619126 41728 619190
rect 41792 619126 41793 619190
rect 41727 619125 41793 619126
rect 40959 617710 41025 617711
rect 40959 617646 40960 617710
rect 41024 617646 41025 617710
rect 40959 617645 41025 617646
rect 40575 603946 40641 603947
rect 40575 603882 40576 603946
rect 40640 603882 40641 603946
rect 40575 603881 40641 603882
rect 40575 599950 40641 599951
rect 40575 599886 40576 599950
rect 40640 599886 40641 599950
rect 40575 599885 40641 599886
rect 40578 573311 40638 599885
rect 40959 596842 41025 596843
rect 40959 596778 40960 596842
rect 41024 596778 41025 596842
rect 40959 596777 41025 596778
rect 40962 574051 41022 596777
rect 41343 584558 41409 584559
rect 41343 584494 41344 584558
rect 41408 584494 41409 584558
rect 41343 584493 41409 584494
rect 40959 574050 41025 574051
rect 40959 573986 40960 574050
rect 41024 573986 41025 574050
rect 40959 573985 41025 573986
rect 41346 573903 41406 584493
rect 41535 584410 41601 584411
rect 41535 584346 41536 584410
rect 41600 584346 41601 584410
rect 41535 584345 41601 584346
rect 41538 577159 41598 584345
rect 41535 577158 41601 577159
rect 41535 577094 41536 577158
rect 41600 577094 41601 577158
rect 41535 577093 41601 577094
rect 41730 574939 41790 619125
rect 41922 618303 41982 661009
rect 42114 646719 42174 688685
rect 42495 684902 42561 684903
rect 42495 684838 42496 684902
rect 42560 684838 42561 684902
rect 42495 684837 42561 684838
rect 42303 678390 42369 678391
rect 42303 678326 42304 678390
rect 42368 678326 42369 678390
rect 42303 678325 42369 678326
rect 42306 668327 42366 678325
rect 42498 668919 42558 684837
rect 42879 682978 42945 682979
rect 42879 682914 42880 682978
rect 42944 682914 42945 682978
rect 42879 682913 42945 682914
rect 42687 670990 42753 670991
rect 42687 670926 42688 670990
rect 42752 670926 42753 670990
rect 42687 670925 42753 670926
rect 42495 668918 42561 668919
rect 42495 668854 42496 668918
rect 42560 668854 42561 668918
rect 42495 668853 42561 668854
rect 42303 668326 42369 668327
rect 42303 668262 42304 668326
rect 42368 668262 42369 668326
rect 42303 668261 42369 668262
rect 42690 663443 42750 670925
rect 42882 666551 42942 682913
rect 43071 670990 43137 670991
rect 43071 670926 43072 670990
rect 43136 670926 43137 670990
rect 43071 670925 43137 670926
rect 42879 666550 42945 666551
rect 42879 666486 42880 666550
rect 42944 666486 42945 666550
rect 42879 666485 42945 666486
rect 43074 665367 43134 670925
rect 43071 665366 43137 665367
rect 43071 665302 43072 665366
rect 43136 665302 43137 665366
rect 43071 665301 43137 665302
rect 42687 663442 42753 663443
rect 42687 663378 42688 663442
rect 42752 663378 42753 663442
rect 42687 663377 42753 663378
rect 673986 648495 674046 697269
rect 674178 666995 674238 741373
rect 674370 670103 674430 743297
rect 675519 740402 675585 740403
rect 675519 740338 675520 740402
rect 675584 740338 675585 740402
rect 675519 740337 675585 740338
rect 674751 739366 674817 739367
rect 674751 739302 674752 739366
rect 674816 739302 674817 739366
rect 674751 739301 674817 739302
rect 674559 694670 674625 694671
rect 674559 694606 674560 694670
rect 674624 694606 674625 694670
rect 674559 694605 674625 694606
rect 674367 670102 674433 670103
rect 674367 670038 674368 670102
rect 674432 670038 674433 670102
rect 674367 670037 674433 670038
rect 674175 666994 674241 666995
rect 674175 666930 674176 666994
rect 674240 666930 674241 666994
rect 674175 666929 674241 666930
rect 673983 648494 674049 648495
rect 673983 648430 673984 648494
rect 674048 648430 674049 648494
rect 673983 648429 674049 648430
rect 674175 648346 674241 648347
rect 674175 648282 674176 648346
rect 674240 648282 674241 648346
rect 674175 648281 674241 648282
rect 42111 646718 42177 646719
rect 42111 646654 42112 646718
rect 42176 646654 42177 646718
rect 42111 646653 42177 646654
rect 674178 642387 674238 648281
rect 674367 645534 674433 645535
rect 674367 645470 674368 645534
rect 674432 645470 674433 645534
rect 674367 645469 674433 645470
rect 673794 642327 674238 642387
rect 42879 635914 42945 635915
rect 42879 635850 42880 635914
rect 42944 635850 42945 635914
rect 42879 635849 42945 635850
rect 42495 634434 42561 634435
rect 42495 634370 42496 634434
rect 42560 634370 42561 634434
rect 42495 634369 42561 634370
rect 42303 627626 42369 627627
rect 42303 627562 42304 627626
rect 42368 627562 42369 627626
rect 42303 627561 42369 627562
rect 42111 627478 42177 627479
rect 42111 627414 42112 627478
rect 42176 627414 42177 627478
rect 42111 627413 42177 627414
rect 42114 624519 42174 627413
rect 42111 624518 42177 624519
rect 42111 624454 42112 624518
rect 42176 624454 42177 624518
rect 42111 624453 42177 624454
rect 42111 624370 42177 624371
rect 42111 624306 42112 624370
rect 42176 624306 42177 624370
rect 42111 624305 42177 624306
rect 42114 620967 42174 624305
rect 42111 620966 42177 620967
rect 42111 620902 42112 620966
rect 42176 620902 42177 620966
rect 42111 620901 42177 620902
rect 42306 620819 42366 627561
rect 42498 622151 42558 634369
rect 42495 622150 42561 622151
rect 42495 622086 42496 622150
rect 42560 622086 42561 622150
rect 42495 622085 42561 622086
rect 42303 620818 42369 620819
rect 42303 620754 42304 620818
rect 42368 620754 42369 620818
rect 42303 620753 42369 620754
rect 42882 618303 42942 635849
rect 673794 630399 673854 642327
rect 674370 637839 674430 645469
rect 674367 637838 674433 637839
rect 674367 637774 674368 637838
rect 674432 637774 674433 637838
rect 674367 637773 674433 637774
rect 674175 630438 674241 630439
rect 673794 630339 674046 630399
rect 674175 630374 674176 630438
rect 674240 630374 674241 630438
rect 674175 630373 674241 630374
rect 673986 624963 674046 630339
rect 673983 624962 674049 624963
rect 673983 624898 673984 624962
rect 674048 624898 674049 624962
rect 673983 624897 674049 624898
rect 674178 618895 674238 630373
rect 674562 621707 674622 694605
rect 674754 666699 674814 739301
rect 675327 738626 675393 738627
rect 675327 738562 675328 738626
rect 675392 738562 675393 738626
rect 675327 738561 675393 738562
rect 675135 697926 675201 697927
rect 675135 697862 675136 697926
rect 675200 697862 675201 697926
rect 675135 697861 675201 697862
rect 674943 696890 675009 696891
rect 674943 696826 674944 696890
rect 675008 696826 675009 696890
rect 674943 696825 675009 696826
rect 674751 666698 674817 666699
rect 674751 666634 674752 666698
rect 674816 666634 674817 666698
rect 674751 666633 674817 666634
rect 674751 652194 674817 652195
rect 674751 652130 674752 652194
rect 674816 652130 674817 652194
rect 674751 652129 674817 652130
rect 674754 639911 674814 652129
rect 674751 639910 674817 639911
rect 674751 639846 674752 639910
rect 674816 639846 674817 639910
rect 674751 639845 674817 639846
rect 674946 639723 675006 696825
rect 675138 641983 675198 697861
rect 675330 665959 675390 738561
rect 675522 669807 675582 740337
rect 675711 734482 675777 734483
rect 675711 734418 675712 734482
rect 675776 734418 675777 734482
rect 675711 734417 675777 734418
rect 675519 669806 675585 669807
rect 675519 669742 675520 669806
rect 675584 669742 675585 669806
rect 675519 669741 675585 669742
rect 675327 665958 675393 665959
rect 675327 665894 675328 665958
rect 675392 665894 675393 665958
rect 675327 665893 675393 665894
rect 675714 664331 675774 734417
rect 675906 717130 675966 786661
rect 676095 784210 676161 784211
rect 676095 784146 676096 784210
rect 676160 784146 676161 784210
rect 676095 784145 676161 784146
rect 675903 717129 675969 717130
rect 675903 717065 675904 717129
rect 675968 717065 675969 717129
rect 675903 717064 675969 717065
rect 676098 711987 676158 784145
rect 676290 715835 676350 787845
rect 676479 781990 676545 781991
rect 676479 781926 676480 781990
rect 676544 781926 676545 781990
rect 676479 781925 676545 781926
rect 676482 736703 676542 781925
rect 676674 757423 676734 876349
rect 677055 780510 677121 780511
rect 677055 780446 677056 780510
rect 677120 780446 677121 780510
rect 677055 780445 677121 780446
rect 677058 780249 677118 780445
rect 677058 780189 677310 780249
rect 677055 777550 677121 777551
rect 677055 777486 677056 777550
rect 677120 777486 677121 777550
rect 677055 777485 677121 777486
rect 676863 777402 676929 777403
rect 676863 777338 676864 777402
rect 676928 777338 676929 777402
rect 676863 777337 676929 777338
rect 676866 773111 676926 777337
rect 676863 773110 676929 773111
rect 676863 773046 676864 773110
rect 676928 773046 676929 773110
rect 676863 773045 676929 773046
rect 676863 772962 676929 772963
rect 676863 772898 676864 772962
rect 676928 772898 676929 772962
rect 676863 772897 676929 772898
rect 676671 757422 676737 757423
rect 676671 757358 676672 757422
rect 676736 757358 676737 757422
rect 676671 757357 676737 757358
rect 676866 753871 676926 772897
rect 676863 753870 676929 753871
rect 676863 753806 676864 753870
rect 676928 753806 676929 753870
rect 676863 753805 676929 753806
rect 676671 741734 676737 741735
rect 676671 741670 676672 741734
rect 676736 741670 676737 741734
rect 676671 741669 676737 741670
rect 676479 736702 676545 736703
rect 676479 736638 676480 736702
rect 676544 736638 676545 736702
rect 676479 736637 676545 736638
rect 676287 715834 676353 715835
rect 676287 715770 676288 715834
rect 676352 715770 676353 715834
rect 676287 715769 676353 715770
rect 676095 711986 676161 711987
rect 676095 711922 676096 711986
rect 676160 711922 676161 711986
rect 676095 711921 676161 711922
rect 676095 694818 676161 694819
rect 676095 694754 676096 694818
rect 676160 694754 676161 694818
rect 676095 694753 676161 694754
rect 675903 693486 675969 693487
rect 675903 693422 675904 693486
rect 675968 693422 675969 693486
rect 675903 693421 675969 693422
rect 675711 664330 675777 664331
rect 675711 664266 675712 664330
rect 675776 664266 675777 664330
rect 675711 664265 675777 664266
rect 675711 659446 675777 659447
rect 675711 659382 675712 659446
rect 675776 659382 675777 659446
rect 675711 659381 675777 659382
rect 675519 659298 675585 659299
rect 675519 659234 675520 659298
rect 675584 659234 675585 659298
rect 675519 659233 675585 659234
rect 675522 652787 675582 659233
rect 675519 652786 675585 652787
rect 675519 652722 675520 652786
rect 675584 652722 675585 652786
rect 675519 652721 675585 652722
rect 675519 652638 675585 652639
rect 675519 652574 675520 652638
rect 675584 652574 675585 652638
rect 675519 652573 675585 652574
rect 675327 651010 675393 651011
rect 675327 650946 675328 651010
rect 675392 650946 675393 651010
rect 675327 650945 675393 650946
rect 675135 641982 675201 641983
rect 675135 641918 675136 641982
rect 675200 641918 675201 641982
rect 675135 641917 675201 641918
rect 674754 639663 675006 639723
rect 674754 627331 674814 639663
rect 674943 639466 675009 639467
rect 674943 639402 674944 639466
rect 675008 639402 675009 639466
rect 674943 639401 675009 639402
rect 674751 627330 674817 627331
rect 674751 627266 674752 627330
rect 674816 627266 674817 627330
rect 674751 627265 674817 627266
rect 674559 621706 674625 621707
rect 674559 621642 674560 621706
rect 674624 621642 674625 621706
rect 674559 621641 674625 621642
rect 674946 620409 675006 639401
rect 675135 638578 675201 638579
rect 675135 638514 675136 638578
rect 675200 638514 675201 638578
rect 675135 638513 675201 638514
rect 674754 620349 675006 620409
rect 674175 618894 674241 618895
rect 674175 618830 674176 618894
rect 674240 618830 674241 618894
rect 674175 618829 674241 618830
rect 41919 618302 41985 618303
rect 41919 618238 41920 618302
rect 41984 618238 41985 618302
rect 41919 618237 41985 618238
rect 42879 618302 42945 618303
rect 42879 618238 42880 618302
rect 42944 618238 42945 618302
rect 42879 618237 42945 618238
rect 41922 575087 41982 618237
rect 674367 607794 674433 607795
rect 674367 607730 674368 607794
rect 674432 607730 674433 607794
rect 674367 607729 674433 607730
rect 673983 604982 674049 604983
rect 673983 604918 673984 604982
rect 674048 604918 674049 604982
rect 673983 604917 674049 604918
rect 42111 603206 42177 603207
rect 42111 603142 42112 603206
rect 42176 603142 42177 603206
rect 42111 603141 42177 603142
rect 41919 575086 41985 575087
rect 41919 575022 41920 575086
rect 41984 575022 41985 575086
rect 41919 575021 41985 575022
rect 41727 574938 41793 574939
rect 41727 574874 41728 574938
rect 41792 574874 41793 574938
rect 41727 574873 41793 574874
rect 41343 573902 41409 573903
rect 41343 573838 41344 573902
rect 41408 573838 41409 573902
rect 41343 573837 41409 573838
rect 40575 573310 40641 573311
rect 40575 573246 40576 573310
rect 40640 573246 40641 573310
rect 40575 573245 40641 573246
rect 40575 556734 40641 556735
rect 40575 556670 40576 556734
rect 40640 556670 40641 556734
rect 40575 556669 40641 556670
rect 40578 532315 40638 556669
rect 40959 553626 41025 553627
rect 40959 553562 40960 553626
rect 41024 553562 41025 553626
rect 40959 553561 41025 553562
rect 40962 532611 41022 553561
rect 40959 532610 41025 532611
rect 40959 532546 40960 532610
rect 41024 532546 41025 532610
rect 40959 532545 41025 532546
rect 40575 532314 40641 532315
rect 40575 532250 40576 532314
rect 40640 532250 40641 532314
rect 40575 532249 40641 532250
rect 41730 531723 41790 574873
rect 41727 531722 41793 531723
rect 41727 531658 41728 531722
rect 41792 531658 41793 531722
rect 41727 531657 41793 531658
rect 40575 431970 40641 431971
rect 40575 431906 40576 431970
rect 40640 431906 40641 431970
rect 40575 431905 40641 431906
rect 40383 425162 40449 425163
rect 40383 425098 40384 425162
rect 40448 425098 40449 425162
rect 40383 425097 40449 425098
rect 40386 402519 40446 425097
rect 40383 402518 40449 402519
rect 40383 402454 40384 402518
rect 40448 402454 40449 402518
rect 40383 402453 40449 402454
rect 40578 388607 40638 431905
rect 40959 430786 41025 430787
rect 40959 430722 40960 430786
rect 41024 430722 41025 430786
rect 40959 430721 41025 430722
rect 40767 429454 40833 429455
rect 40767 429390 40768 429454
rect 40832 429390 40833 429454
rect 40767 429389 40833 429390
rect 40770 398819 40830 429389
rect 40962 400151 41022 430721
rect 41343 428418 41409 428419
rect 41343 428354 41344 428418
rect 41408 428354 41409 428418
rect 41343 428353 41409 428354
rect 41151 426346 41217 426347
rect 41151 426282 41152 426346
rect 41216 426282 41217 426346
rect 41151 426281 41217 426282
rect 40959 400150 41025 400151
rect 40959 400086 40960 400150
rect 41024 400086 41025 400150
rect 40959 400085 41025 400086
rect 41154 399559 41214 426281
rect 41346 402075 41406 428353
rect 41535 427678 41601 427679
rect 41535 427614 41536 427678
rect 41600 427614 41601 427678
rect 41535 427613 41601 427614
rect 41538 406071 41598 427613
rect 41730 419095 41790 531657
rect 41922 531279 41982 575021
rect 42114 561027 42174 603141
rect 43071 586630 43137 586631
rect 43071 586566 43072 586630
rect 43136 586566 43137 586630
rect 43071 586565 43137 586566
rect 42495 585002 42561 585003
rect 42495 584938 42496 585002
rect 42560 584938 42561 585002
rect 42495 584937 42561 584938
rect 42303 584262 42369 584263
rect 42303 584198 42304 584262
rect 42368 584198 42369 584262
rect 42303 584197 42369 584198
rect 42306 581303 42366 584197
rect 42303 581302 42369 581303
rect 42303 581238 42304 581302
rect 42368 581238 42369 581302
rect 42303 581237 42369 581238
rect 42498 577011 42558 584937
rect 42879 584410 42945 584411
rect 42879 584346 42880 584410
rect 42944 584346 42945 584410
rect 42879 584345 42945 584346
rect 42882 578343 42942 584345
rect 42879 578342 42945 578343
rect 42879 578278 42880 578342
rect 42944 578278 42945 578342
rect 42879 578277 42945 578278
rect 43074 577603 43134 586565
rect 673986 584559 674046 604917
rect 674175 604834 674241 604835
rect 674175 604770 674176 604834
rect 674240 604770 674241 604834
rect 674175 604769 674241 604770
rect 674178 584559 674238 604769
rect 673983 584558 674049 584559
rect 673983 584494 673984 584558
rect 674048 584494 674049 584558
rect 673983 584493 674049 584494
rect 674175 584558 674241 584559
rect 674175 584494 674176 584558
rect 674240 584494 674241 584558
rect 674175 584493 674241 584494
rect 673983 584114 674049 584115
rect 673983 584050 673984 584114
rect 674048 584050 674049 584114
rect 673983 584049 674049 584050
rect 43071 577602 43137 577603
rect 43071 577538 43072 577602
rect 43136 577538 43137 577602
rect 43071 577537 43137 577538
rect 42495 577010 42561 577011
rect 42495 576946 42496 577010
rect 42560 576946 42561 577010
rect 42495 576945 42561 576946
rect 42111 561026 42177 561027
rect 42111 560962 42112 561026
rect 42176 560962 42177 561026
rect 42111 560961 42177 560962
rect 42687 541342 42753 541343
rect 42687 541278 42688 541342
rect 42752 541278 42753 541342
rect 42687 541277 42753 541278
rect 42111 541194 42177 541195
rect 42111 541130 42112 541194
rect 42176 541130 42177 541194
rect 42111 541129 42177 541130
rect 42114 538975 42174 541129
rect 42111 538974 42177 538975
rect 42111 538910 42112 538974
rect 42176 538910 42177 538974
rect 42111 538909 42177 538910
rect 42690 538679 42750 541277
rect 43071 541046 43137 541047
rect 43071 540982 43072 541046
rect 43136 540982 43137 541046
rect 43071 540981 43137 540982
rect 42687 538678 42753 538679
rect 42687 538614 42688 538678
rect 42752 538614 42753 538678
rect 42687 538613 42753 538614
rect 43074 536903 43134 540981
rect 43071 536902 43137 536903
rect 43071 536838 43072 536902
rect 43136 536838 43137 536902
rect 43071 536837 43137 536838
rect 673986 534091 674046 584049
rect 674175 561766 674241 561767
rect 674175 561702 674176 561766
rect 674240 561702 674241 561766
rect 674175 561701 674241 561702
rect 673983 534090 674049 534091
rect 673983 534026 673984 534090
rect 674048 534026 674049 534090
rect 673983 534025 674049 534026
rect 41919 531278 41985 531279
rect 41919 531214 41920 531278
rect 41984 531214 41985 531278
rect 41919 531213 41985 531214
rect 41727 419094 41793 419095
rect 41727 419030 41728 419094
rect 41792 419030 41793 419094
rect 41727 419029 41793 419030
rect 41535 406070 41601 406071
rect 41535 406006 41536 406070
rect 41600 406006 41601 406070
rect 41535 406005 41601 406006
rect 41922 405291 41982 531213
rect 674178 487767 674238 561701
rect 674370 534905 674430 607729
rect 674559 607498 674625 607499
rect 674559 607434 674560 607498
rect 674624 607434 674625 607498
rect 674559 607433 674625 607434
rect 674367 534904 674433 534905
rect 674367 534840 674368 534904
rect 674432 534840 674433 534904
rect 674367 534839 674433 534840
rect 674562 532315 674622 607433
rect 674754 577307 674814 620349
rect 674943 599210 675009 599211
rect 674943 599146 674944 599210
rect 675008 599146 675009 599210
rect 674943 599145 675009 599146
rect 674946 578195 675006 599145
rect 675138 578195 675198 638513
rect 675330 581747 675390 650945
rect 675327 581746 675393 581747
rect 675327 581682 675328 581746
rect 675392 581682 675393 581746
rect 675327 581681 675393 581682
rect 675522 580415 675582 652573
rect 675714 640799 675774 659381
rect 675906 645091 675966 693421
rect 675903 645090 675969 645091
rect 675903 645026 675904 645090
rect 675968 645026 675969 645090
rect 675903 645025 675969 645026
rect 675711 640798 675777 640799
rect 675711 640734 675712 640798
rect 675776 640734 675777 640798
rect 675711 640733 675777 640734
rect 676098 633251 676158 694753
rect 676482 691711 676542 736637
rect 676479 691710 676545 691711
rect 676479 691646 676480 691710
rect 676544 691646 676545 691710
rect 676479 691645 676545 691646
rect 676287 679722 676353 679723
rect 676287 679658 676288 679722
rect 676352 679658 676353 679722
rect 676287 679657 676353 679658
rect 676290 672323 676350 679657
rect 676287 672322 676353 672323
rect 676287 672258 676288 672322
rect 676352 672258 676353 672322
rect 676287 672257 676353 672258
rect 676482 659299 676542 691645
rect 676674 689343 676734 741669
rect 676863 732558 676929 732559
rect 676863 732494 676864 732558
rect 676928 732494 676929 732558
rect 676863 732493 676929 732494
rect 676671 689342 676737 689343
rect 676671 689278 676672 689342
rect 676736 689278 676737 689342
rect 676671 689277 676737 689278
rect 676671 689194 676737 689195
rect 676671 689130 676672 689194
rect 676736 689130 676737 689194
rect 676671 689129 676737 689130
rect 676674 659447 676734 689129
rect 676866 662407 676926 732493
rect 677058 708435 677118 777485
rect 677250 772963 677310 780189
rect 677823 773110 677889 773111
rect 677823 773046 677824 773110
rect 677888 773046 677889 773110
rect 677823 773045 677889 773046
rect 677247 772962 677313 772963
rect 677247 772898 677248 772962
rect 677312 772898 677313 772962
rect 677247 772897 677313 772898
rect 677247 772666 677313 772667
rect 677247 772602 677248 772666
rect 677312 772602 677313 772666
rect 677247 772601 677313 772602
rect 677250 754463 677310 772601
rect 677247 754462 677313 754463
rect 677247 754398 677248 754462
rect 677312 754398 677313 754462
rect 677247 754397 677313 754398
rect 677826 752983 677886 773045
rect 677823 752982 677889 752983
rect 677823 752918 677824 752982
rect 677888 752918 677889 752982
rect 677823 752917 677889 752918
rect 677055 708434 677121 708435
rect 677055 708370 677056 708434
rect 677120 708370 677121 708434
rect 677055 708369 677121 708370
rect 677055 688306 677121 688307
rect 677055 688242 677056 688306
rect 677120 688242 677121 688306
rect 677055 688241 677121 688242
rect 677058 687675 677118 688241
rect 677058 687615 677310 687675
rect 677055 685642 677121 685643
rect 677055 685578 677056 685642
rect 677120 685578 677121 685642
rect 677055 685577 677121 685578
rect 676863 662406 676929 662407
rect 676863 662342 676864 662406
rect 676928 662342 676929 662406
rect 676863 662341 676929 662342
rect 676671 659446 676737 659447
rect 676671 659382 676672 659446
rect 676736 659382 676737 659446
rect 676671 659381 676737 659382
rect 676479 659298 676545 659299
rect 676479 659234 676480 659298
rect 676544 659234 676545 659298
rect 676479 659233 676545 659234
rect 676287 649678 676353 649679
rect 676287 649614 676288 649678
rect 676352 649614 676353 649678
rect 676287 649613 676353 649614
rect 676095 633250 676161 633251
rect 676095 633186 676096 633250
rect 676160 633186 676161 633250
rect 676095 633185 676161 633186
rect 676095 630142 676161 630143
rect 676095 630078 676096 630142
rect 676160 630078 676161 630142
rect 676095 630077 676161 630078
rect 675711 606462 675777 606463
rect 675711 606398 675712 606462
rect 675776 606398 675777 606462
rect 675711 606397 675777 606398
rect 675519 580414 675585 580415
rect 675519 580350 675520 580414
rect 675584 580350 675585 580414
rect 675519 580349 675585 580350
rect 674943 578194 675009 578195
rect 674943 578130 674944 578194
rect 675008 578130 675009 578194
rect 674943 578129 675009 578130
rect 675135 578194 675201 578195
rect 675135 578130 675136 578194
rect 675200 578130 675201 578194
rect 675135 578129 675201 578130
rect 674751 577306 674817 577307
rect 674751 577242 674752 577306
rect 674816 577242 674817 577306
rect 674751 577241 674817 577242
rect 675519 567390 675585 567391
rect 675519 567326 675520 567390
rect 675584 567326 675585 567390
rect 675519 567325 675585 567326
rect 674943 562950 675009 562951
rect 674943 562886 674944 562950
rect 675008 562886 675009 562950
rect 674943 562885 675009 562886
rect 674751 558954 674817 558955
rect 674751 558890 674752 558954
rect 674816 558890 674817 558954
rect 674751 558889 674817 558890
rect 674559 532314 674625 532315
rect 674559 532250 674560 532314
rect 674624 532250 674625 532314
rect 674559 532249 674625 532250
rect 674175 487766 674241 487767
rect 674175 487702 674176 487766
rect 674240 487702 674241 487766
rect 674175 487701 674241 487702
rect 674754 487471 674814 558889
rect 674946 491467 675006 562885
rect 675135 561618 675201 561619
rect 675135 561554 675136 561618
rect 675200 561554 675201 561618
rect 675135 561553 675201 561554
rect 675138 492799 675198 561553
rect 675522 538383 675582 567325
rect 675519 538382 675585 538383
rect 675519 538318 675520 538382
rect 675584 538318 675585 538382
rect 675519 538317 675585 538318
rect 675714 537051 675774 606397
rect 675903 600246 675969 600247
rect 675903 600182 675904 600246
rect 675968 600182 675969 600246
rect 675903 600181 675969 600182
rect 675711 537050 675777 537051
rect 675711 536986 675712 537050
rect 675776 536986 675777 537050
rect 675711 536985 675777 536986
rect 675906 533795 675966 600181
rect 676098 599211 676158 630077
rect 676095 599210 676161 599211
rect 676095 599146 676096 599210
rect 676160 599146 676161 599210
rect 676095 599145 676161 599146
rect 676095 593438 676161 593439
rect 676095 593374 676096 593438
rect 676160 593374 676161 593438
rect 676095 593373 676161 593374
rect 675903 533794 675969 533795
rect 675903 533730 675904 533794
rect 675968 533730 675969 533794
rect 675903 533729 675969 533730
rect 676098 532759 676158 593373
rect 676290 579675 676350 649613
rect 676479 648494 676545 648495
rect 676479 648430 676480 648494
rect 676544 648430 676545 648494
rect 676479 648429 676545 648430
rect 676482 640503 676542 648429
rect 676863 644942 676929 644943
rect 676863 644878 676864 644942
rect 676928 644878 676929 644942
rect 676863 644877 676929 644878
rect 676671 640798 676737 640799
rect 676671 640734 676672 640798
rect 676736 640734 676737 640798
rect 676671 640733 676737 640734
rect 676479 640502 676545 640503
rect 676479 640438 676480 640502
rect 676544 640438 676545 640502
rect 676479 640437 676545 640438
rect 676479 640354 676545 640355
rect 676479 640290 676480 640354
rect 676544 640290 676545 640354
rect 676479 640289 676545 640290
rect 676482 581303 676542 640289
rect 676674 630399 676734 640733
rect 676866 635027 676926 644877
rect 676863 635026 676929 635027
rect 676863 634962 676864 635026
rect 676928 634962 676929 635026
rect 676863 634961 676929 634962
rect 676863 630438 676929 630439
rect 676863 630399 676864 630438
rect 676674 630374 676864 630399
rect 676928 630374 676929 630438
rect 676674 630373 676929 630374
rect 676674 630339 676926 630373
rect 676671 630142 676737 630143
rect 676671 630078 676672 630142
rect 676736 630078 676737 630142
rect 676671 630077 676737 630078
rect 676674 620967 676734 630077
rect 676671 620966 676737 620967
rect 676671 620902 676672 620966
rect 676736 620902 676737 620966
rect 676671 620901 676737 620902
rect 677058 617859 677118 685577
rect 677250 663591 677310 687615
rect 677247 663590 677313 663591
rect 677247 663526 677248 663590
rect 677312 663526 677313 663590
rect 677247 663525 677313 663526
rect 677055 617858 677121 617859
rect 677055 617794 677056 617858
rect 677120 617794 677121 617858
rect 677055 617793 677121 617794
rect 676671 595362 676737 595363
rect 676671 595298 676672 595362
rect 676736 595298 676737 595362
rect 676671 595297 676737 595298
rect 676479 581302 676545 581303
rect 676479 581238 676480 581302
rect 676544 581238 676545 581302
rect 676479 581237 676545 581238
rect 676287 579674 676353 579675
rect 676287 579610 676288 579674
rect 676352 579610 676353 579674
rect 676287 579609 676353 579610
rect 676287 557770 676353 557771
rect 676287 557706 676288 557770
rect 676352 557706 676353 557770
rect 676287 557705 676353 557706
rect 676095 532758 676161 532759
rect 676095 532694 676096 532758
rect 676160 532694 676161 532758
rect 676095 532693 676161 532694
rect 675135 492798 675201 492799
rect 675135 492734 675136 492798
rect 675200 492734 675201 492798
rect 675135 492733 675201 492734
rect 674943 491466 675009 491467
rect 674943 491402 674944 491466
rect 675008 491402 675009 491466
rect 674943 491401 675009 491402
rect 674751 487470 674817 487471
rect 674751 487406 674752 487470
rect 674816 487406 674817 487470
rect 674751 487405 674817 487406
rect 676290 484067 676350 557705
rect 676674 536311 676734 595297
rect 676863 581894 676929 581895
rect 676863 581830 676864 581894
rect 676928 581830 676929 581894
rect 676863 581829 676929 581830
rect 676866 547115 676926 581829
rect 676863 547114 676929 547115
rect 676863 547050 676864 547114
rect 676928 547050 676929 547114
rect 676863 547049 676929 547050
rect 676671 536310 676737 536311
rect 676671 536246 676672 536310
rect 676736 536246 676737 536310
rect 676671 536245 676737 536246
rect 676287 484066 676353 484067
rect 676287 484002 676288 484066
rect 676352 484002 676353 484066
rect 676287 484001 676353 484002
rect 673983 475334 674049 475335
rect 673983 475270 673984 475334
rect 674048 475270 674049 475334
rect 673983 475269 674049 475270
rect 42111 432710 42177 432711
rect 42111 432646 42112 432710
rect 42176 432646 42177 432710
rect 42111 432645 42177 432646
rect 41538 405231 41982 405291
rect 41538 403851 41598 405231
rect 41727 404294 41793 404295
rect 41727 404230 41728 404294
rect 41792 404230 41793 404294
rect 41727 404229 41793 404230
rect 41535 403850 41601 403851
rect 41535 403786 41536 403850
rect 41600 403786 41601 403850
rect 41535 403785 41601 403786
rect 41343 402074 41409 402075
rect 41343 402010 41344 402074
rect 41408 402010 41409 402074
rect 41343 402009 41409 402010
rect 41151 399558 41217 399559
rect 41151 399494 41152 399558
rect 41216 399494 41217 399558
rect 41151 399493 41217 399494
rect 40767 398818 40833 398819
rect 40767 398754 40768 398818
rect 40832 398754 40833 398818
rect 40767 398753 40833 398754
rect 40575 388606 40641 388607
rect 40575 388542 40576 388606
rect 40640 388542 40641 388606
rect 40575 388541 40641 388542
rect 40578 368775 40638 388541
rect 40959 387570 41025 387571
rect 40959 387506 40960 387570
rect 41024 387506 41025 387570
rect 40959 387505 41025 387506
rect 40767 386090 40833 386091
rect 40767 386026 40768 386090
rect 40832 386026 40833 386090
rect 40767 386025 40833 386026
rect 40575 368774 40641 368775
rect 40575 368710 40576 368774
rect 40640 368710 40641 368774
rect 40575 368709 40641 368710
rect 40383 363002 40449 363003
rect 40383 362938 40384 363002
rect 40448 362938 40449 363002
rect 40383 362937 40449 362938
rect 40386 355341 40446 362937
rect 40770 355603 40830 386025
rect 40962 356935 41022 387505
rect 41343 385202 41409 385203
rect 41343 385138 41344 385202
rect 41408 385138 41409 385202
rect 41343 385137 41409 385138
rect 41151 383130 41217 383131
rect 41151 383066 41152 383130
rect 41216 383066 41217 383130
rect 41151 383065 41217 383066
rect 40959 356934 41025 356935
rect 40959 356870 40960 356934
rect 41024 356870 41025 356934
rect 40959 356869 41025 356870
rect 41154 356491 41214 383065
rect 41346 358711 41406 385137
rect 41535 384462 41601 384463
rect 41535 384398 41536 384462
rect 41600 384398 41601 384462
rect 41535 384397 41601 384398
rect 41538 362855 41598 384397
rect 41730 372657 41790 404229
rect 42114 390235 42174 432645
rect 42303 419094 42369 419095
rect 42303 419030 42304 419094
rect 42368 419030 42369 419094
rect 42303 419029 42369 419030
rect 42306 404295 42366 419029
rect 673986 405923 674046 475269
rect 676671 411990 676737 411991
rect 676671 411926 676672 411990
rect 676736 411926 676737 411990
rect 676671 411925 676737 411926
rect 673983 405922 674049 405923
rect 673983 405858 673984 405922
rect 674048 405858 674049 405922
rect 673983 405857 674049 405858
rect 42303 404294 42369 404295
rect 42303 404230 42304 404294
rect 42368 404230 42369 404294
rect 42303 404229 42369 404230
rect 42687 403850 42753 403851
rect 42687 403786 42688 403850
rect 42752 403786 42753 403850
rect 42687 403785 42753 403786
rect 42111 390234 42177 390235
rect 42111 390170 42112 390234
rect 42176 390170 42177 390234
rect 42111 390169 42177 390170
rect 42495 389494 42561 389495
rect 42495 389430 42496 389494
rect 42560 389430 42561 389494
rect 42495 389429 42561 389430
rect 42111 381946 42177 381947
rect 42111 381882 42112 381946
rect 42176 381882 42177 381946
rect 42111 381881 42177 381882
rect 41730 372597 41982 372657
rect 41727 368626 41793 368627
rect 41727 368562 41728 368626
rect 41792 368562 41793 368626
rect 41727 368561 41793 368562
rect 41730 363151 41790 368561
rect 41922 368331 41982 372597
rect 42114 368775 42174 381881
rect 42111 368774 42177 368775
rect 42111 368710 42112 368774
rect 42176 368710 42177 368774
rect 42111 368709 42177 368710
rect 42111 368478 42177 368479
rect 42111 368414 42112 368478
rect 42176 368414 42177 368478
rect 42111 368413 42177 368414
rect 41919 368330 41985 368331
rect 41919 368266 41920 368330
rect 41984 368266 41985 368330
rect 41919 368265 41985 368266
rect 41727 363150 41793 363151
rect 41727 363086 41728 363150
rect 41792 363086 41793 363150
rect 41727 363085 41793 363086
rect 41535 362854 41601 362855
rect 41535 362790 41536 362854
rect 41600 362790 41601 362854
rect 41535 362789 41601 362790
rect 41727 360634 41793 360635
rect 41727 360570 41728 360634
rect 41792 360570 41793 360634
rect 41727 360569 41793 360570
rect 41343 358710 41409 358711
rect 41343 358646 41344 358710
rect 41408 358646 41409 358710
rect 41343 358645 41409 358646
rect 41151 356490 41217 356491
rect 41151 356426 41152 356490
rect 41216 356426 41217 356490
rect 41151 356425 41217 356426
rect 40767 355602 40833 355603
rect 40767 355538 40768 355602
rect 40832 355538 40833 355602
rect 40767 355537 40833 355538
rect 40386 355281 41406 355341
rect 41346 345983 41406 355281
rect 41343 345982 41409 345983
rect 41343 345918 41344 345982
rect 41408 345918 41409 345982
rect 41343 345917 41409 345918
rect 40767 344354 40833 344355
rect 40767 344290 40768 344354
rect 40832 344290 40833 344354
rect 40767 344289 40833 344290
rect 40383 338730 40449 338731
rect 40383 338666 40384 338730
rect 40448 338666 40449 338730
rect 40383 338665 40449 338666
rect 40386 316087 40446 338665
rect 40383 316086 40449 316087
rect 40383 316022 40384 316086
rect 40448 316022 40449 316086
rect 40383 316021 40449 316022
rect 40770 313719 40830 344289
rect 40959 342874 41025 342875
rect 40959 342810 40960 342874
rect 41024 342810 41025 342874
rect 40959 342809 41025 342810
rect 40767 313718 40833 313719
rect 40767 313654 40768 313718
rect 40832 313654 40833 313718
rect 40767 313653 40833 313654
rect 40962 312387 41022 342809
rect 41343 341986 41409 341987
rect 41343 341922 41344 341986
rect 41408 341922 41409 341986
rect 41343 341921 41409 341922
rect 41151 339914 41217 339915
rect 41151 339850 41152 339914
rect 41216 339850 41217 339914
rect 41151 339849 41217 339850
rect 41154 313275 41214 339849
rect 41346 315643 41406 341921
rect 41535 341246 41601 341247
rect 41535 341182 41536 341246
rect 41600 341182 41601 341246
rect 41535 341181 41601 341182
rect 41538 319787 41598 341181
rect 41535 319786 41601 319787
rect 41535 319722 41536 319786
rect 41600 319722 41601 319786
rect 41535 319721 41601 319722
rect 41535 318750 41601 318751
rect 41535 318686 41536 318750
rect 41600 318686 41601 318750
rect 41535 318685 41601 318686
rect 41343 315642 41409 315643
rect 41343 315578 41344 315642
rect 41408 315578 41409 315642
rect 41343 315577 41409 315578
rect 41151 313274 41217 313275
rect 41151 313210 41152 313274
rect 41216 313210 41217 313274
rect 41151 313209 41217 313210
rect 40959 312386 41025 312387
rect 40959 312322 40960 312386
rect 41024 312322 41025 312386
rect 40959 312321 41025 312322
rect 40575 302766 40641 302767
rect 40575 302702 40576 302766
rect 40640 302702 40641 302766
rect 40575 302701 40641 302702
rect 40383 295514 40449 295515
rect 40383 295450 40384 295514
rect 40448 295450 40449 295514
rect 40383 295449 40449 295450
rect 40386 272871 40446 295449
rect 40383 272870 40449 272871
rect 40383 272806 40384 272870
rect 40448 272806 40449 272870
rect 40383 272805 40449 272806
rect 40578 259551 40638 302701
rect 40959 301138 41025 301139
rect 40959 301074 40960 301138
rect 41024 301074 41025 301138
rect 40959 301073 41025 301074
rect 40767 299658 40833 299659
rect 40767 299594 40768 299658
rect 40832 299594 40833 299658
rect 40767 299593 40833 299594
rect 40770 269171 40830 299593
rect 40962 270651 41022 301073
rect 41538 298771 41598 318685
rect 41730 318011 41790 360569
rect 42114 359451 42174 368413
rect 42303 368330 42369 368331
rect 42303 368266 42304 368330
rect 42368 368266 42369 368330
rect 42303 368265 42369 368266
rect 42306 360931 42366 368265
rect 42303 360930 42369 360931
rect 42303 360866 42304 360930
rect 42368 360866 42369 360930
rect 42303 360865 42369 360866
rect 42111 359450 42177 359451
rect 42111 359386 42112 359450
rect 42176 359386 42177 359450
rect 42111 359385 42177 359386
rect 42306 346683 42366 360865
rect 42498 346871 42558 389429
rect 42690 360635 42750 403785
rect 673986 360783 674046 405857
rect 676674 405331 676734 411925
rect 675327 405330 675393 405331
rect 675327 405266 675328 405330
rect 675392 405266 675393 405330
rect 675327 405265 675393 405266
rect 676671 405330 676737 405331
rect 676671 405266 676672 405330
rect 676736 405266 676737 405330
rect 676671 405265 676737 405266
rect 674175 403554 674241 403555
rect 674175 403490 674176 403554
rect 674240 403490 674241 403554
rect 674175 403489 674241 403490
rect 674178 373955 674238 403489
rect 674559 400594 674625 400595
rect 674559 400530 674560 400594
rect 674624 400530 674625 400594
rect 674559 400529 674625 400530
rect 674367 400446 674433 400447
rect 674367 400382 674368 400446
rect 674432 400382 674433 400446
rect 674367 400381 674433 400382
rect 674175 373954 674241 373955
rect 674175 373890 674176 373954
rect 674240 373890 674241 373954
rect 674175 373889 674241 373890
rect 674370 372031 674430 400381
rect 674562 378839 674622 400529
rect 674559 378838 674625 378839
rect 674559 378774 674560 378838
rect 674624 378774 674625 378838
rect 674559 378773 674625 378774
rect 674367 372030 674433 372031
rect 674367 371966 674368 372030
rect 674432 371966 674433 372030
rect 674367 371965 674433 371966
rect 674175 361448 674241 361449
rect 674175 361384 674176 361448
rect 674240 361384 674241 361448
rect 674175 361383 674241 361384
rect 673983 360782 674049 360783
rect 673983 360718 673984 360782
rect 674048 360718 674049 360782
rect 673983 360717 674049 360718
rect 42687 360634 42753 360635
rect 42687 360570 42688 360634
rect 42752 360570 42753 360634
rect 42687 360569 42753 360570
rect 42495 346870 42561 346871
rect 42495 346806 42496 346870
rect 42560 346806 42561 346870
rect 42495 346805 42561 346806
rect 42306 346623 42558 346683
rect 42111 346130 42177 346131
rect 42111 346066 42112 346130
rect 42176 346066 42177 346130
rect 42111 346065 42177 346066
rect 41919 335622 41985 335623
rect 41919 335558 41920 335622
rect 41984 335558 41985 335622
rect 41919 335557 41985 335558
rect 41727 318010 41793 318011
rect 41727 317946 41728 318010
rect 41792 317946 41793 318010
rect 41727 317945 41793 317946
rect 41730 313867 41790 317945
rect 41922 317419 41982 335557
rect 41919 317418 41985 317419
rect 41919 317354 41920 317418
rect 41984 317354 41985 317418
rect 41919 317353 41985 317354
rect 41727 313866 41793 313867
rect 41727 313802 41728 313866
rect 41792 313802 41793 313866
rect 41727 313801 41793 313802
rect 42114 302767 42174 346065
rect 42303 345982 42369 345983
rect 42303 345918 42304 345982
rect 42368 345918 42369 345982
rect 42303 345917 42369 345918
rect 42306 302767 42366 345917
rect 42498 342727 42558 346623
rect 42495 342726 42561 342727
rect 42495 342662 42496 342726
rect 42560 342662 42561 342726
rect 42495 342661 42561 342662
rect 43071 342726 43137 342727
rect 43071 342662 43072 342726
rect 43136 342662 43137 342726
rect 43071 342661 43137 342662
rect 43074 318751 43134 342661
rect 43071 318750 43137 318751
rect 43071 318686 43072 318750
rect 43136 318686 43137 318750
rect 43071 318685 43137 318686
rect 674178 317271 674238 361383
rect 675330 360191 675390 405265
rect 675519 374546 675585 374547
rect 675519 374482 675520 374546
rect 675584 374482 675585 374546
rect 675519 374481 675585 374482
rect 675327 360190 675393 360191
rect 675327 360126 675328 360190
rect 675392 360126 675393 360190
rect 675327 360125 675393 360126
rect 674367 358266 674433 358267
rect 674367 358202 674368 358266
rect 674432 358202 674433 358266
rect 674367 358201 674433 358202
rect 674370 328371 674430 358201
rect 674751 355454 674817 355455
rect 674751 355390 674752 355454
rect 674816 355390 674817 355454
rect 674751 355389 674817 355390
rect 674559 354566 674625 354567
rect 674559 354502 674560 354566
rect 674624 354502 674625 354566
rect 674559 354501 674625 354502
rect 674367 328370 674433 328371
rect 674367 328306 674368 328370
rect 674432 328306 674433 328370
rect 674367 328305 674433 328306
rect 674562 326891 674622 354501
rect 674754 333551 674814 355389
rect 675135 351458 675201 351459
rect 675135 351394 675136 351458
rect 675200 351394 675201 351458
rect 675135 351393 675201 351394
rect 674943 345538 675009 345539
rect 674943 345474 674944 345538
rect 675008 345474 675009 345538
rect 674943 345473 675009 345474
rect 674751 333550 674817 333551
rect 674751 333486 674752 333550
rect 674816 333486 674817 333550
rect 674751 333485 674817 333486
rect 674559 326890 674625 326891
rect 674559 326826 674560 326890
rect 674624 326826 674625 326890
rect 674559 326825 674625 326826
rect 674175 317270 674241 317271
rect 674175 317206 674176 317270
rect 674240 317206 674241 317270
rect 674175 317205 674241 317206
rect 674175 316456 674241 316457
rect 674175 316392 674176 316456
rect 674240 316392 674241 316456
rect 674175 316391 674241 316392
rect 673983 314902 674049 314903
rect 673983 314838 673984 314902
rect 674048 314838 674049 314902
rect 673983 314837 674049 314838
rect 43071 313866 43137 313867
rect 43071 313802 43072 313866
rect 43136 313802 43137 313866
rect 43071 313801 43137 313802
rect 42111 302766 42177 302767
rect 42111 302702 42112 302766
rect 42176 302702 42177 302766
rect 42111 302701 42177 302702
rect 42303 302766 42369 302767
rect 42303 302702 42304 302766
rect 42368 302702 42369 302766
rect 42303 302701 42369 302702
rect 41343 298770 41409 298771
rect 41343 298706 41344 298770
rect 41408 298706 41409 298770
rect 41343 298705 41409 298706
rect 41535 298770 41601 298771
rect 41535 298706 41536 298770
rect 41600 298706 41601 298770
rect 41535 298705 41601 298706
rect 41151 296698 41217 296699
rect 41151 296634 41152 296698
rect 41216 296634 41217 296698
rect 41151 296633 41217 296634
rect 40959 270650 41025 270651
rect 40959 270586 40960 270650
rect 41024 270586 41025 270650
rect 40959 270585 41025 270586
rect 41154 270059 41214 296633
rect 41346 272427 41406 298705
rect 41535 298030 41601 298031
rect 41535 297966 41536 298030
rect 41600 297966 41601 298030
rect 41535 297965 41601 297966
rect 41538 276571 41598 297965
rect 41919 282342 41985 282343
rect 41919 282278 41920 282342
rect 41984 282278 41985 282342
rect 41919 282277 41985 282278
rect 41535 276570 41601 276571
rect 41535 276506 41536 276570
rect 41600 276506 41601 276570
rect 41535 276505 41601 276506
rect 41922 274795 41982 282277
rect 41919 274794 41985 274795
rect 41919 274730 41920 274794
rect 41984 274730 41985 274794
rect 41919 274729 41985 274730
rect 41727 274054 41793 274055
rect 41727 273990 41728 274054
rect 41792 273990 41793 274054
rect 41727 273989 41793 273990
rect 41343 272426 41409 272427
rect 41343 272362 41344 272426
rect 41408 272362 41409 272426
rect 41343 272361 41409 272362
rect 41151 270058 41217 270059
rect 41151 269994 41152 270058
rect 41216 269994 41217 270058
rect 41151 269993 41217 269994
rect 40767 269170 40833 269171
rect 40767 269106 40768 269170
rect 40832 269106 40833 269170
rect 40767 269105 40833 269106
rect 40575 259550 40641 259551
rect 40575 259486 40576 259550
rect 40640 259486 40641 259550
rect 40575 259485 40641 259486
rect 40383 257922 40449 257923
rect 40383 257858 40384 257922
rect 40448 257858 40449 257922
rect 40383 257857 40449 257858
rect 40386 227287 40446 257857
rect 40575 256442 40641 256443
rect 40575 256378 40576 256442
rect 40640 256378 40641 256442
rect 40575 256377 40641 256378
rect 40578 247859 40638 256377
rect 40959 255702 41025 255703
rect 40959 255638 40960 255702
rect 41024 255638 41025 255702
rect 40959 255637 41025 255638
rect 40767 253482 40833 253483
rect 40767 253418 40768 253482
rect 40832 253418 40833 253482
rect 40767 253417 40833 253418
rect 40575 247858 40641 247859
rect 40575 247794 40576 247858
rect 40640 247794 40641 247858
rect 40575 247793 40641 247794
rect 40575 227582 40641 227583
rect 40575 227518 40576 227582
rect 40640 227518 40641 227582
rect 40575 227517 40641 227518
rect 40383 227286 40449 227287
rect 40383 227222 40384 227286
rect 40448 227222 40449 227286
rect 40383 227221 40449 227222
rect 40578 225955 40638 227517
rect 40770 226843 40830 253417
rect 40962 229063 41022 255637
rect 41343 254814 41409 254815
rect 41343 254750 41344 254814
rect 41408 254750 41409 254814
rect 41343 254749 41409 254750
rect 41151 252446 41217 252447
rect 41151 252382 41152 252446
rect 41216 252382 41217 252446
rect 41151 252381 41217 252382
rect 41154 229803 41214 252381
rect 41346 233355 41406 254749
rect 41535 247710 41601 247711
rect 41535 247646 41536 247710
rect 41600 247646 41601 247710
rect 41535 247645 41601 247646
rect 41343 233354 41409 233355
rect 41343 233290 41344 233354
rect 41408 233290 41409 233354
rect 41343 233289 41409 233290
rect 41151 229802 41217 229803
rect 41151 229738 41152 229802
rect 41216 229738 41217 229802
rect 41151 229737 41217 229738
rect 40959 229062 41025 229063
rect 40959 228998 40960 229062
rect 41024 228998 41025 229062
rect 40959 228997 41025 228998
rect 41538 227583 41598 247645
rect 41730 231727 41790 273989
rect 41727 231726 41793 231727
rect 41727 231662 41728 231726
rect 41792 231662 41793 231726
rect 41727 231661 41793 231662
rect 41535 227582 41601 227583
rect 41535 227518 41536 227582
rect 41600 227518 41601 227582
rect 41535 227517 41601 227518
rect 40767 226842 40833 226843
rect 40767 226778 40768 226842
rect 40832 226778 40833 226842
rect 40767 226777 40833 226778
rect 40575 225954 40641 225955
rect 40575 225890 40576 225954
rect 40640 225890 40641 225954
rect 40575 225889 40641 225890
rect 40575 214706 40641 214707
rect 40575 214642 40576 214706
rect 40640 214642 40641 214706
rect 40575 214641 40641 214642
rect 40383 213226 40449 213227
rect 40383 213162 40384 213226
rect 40448 213162 40449 213226
rect 40383 213161 40449 213162
rect 40386 182887 40446 213161
rect 40578 184219 40638 214641
rect 40959 212486 41025 212487
rect 40959 212422 40960 212486
rect 41024 212422 41025 212486
rect 40959 212421 41025 212422
rect 40767 210414 40833 210415
rect 40767 210350 40768 210414
rect 40832 210350 40833 210414
rect 40767 210349 40833 210350
rect 40575 184218 40641 184219
rect 40575 184154 40576 184218
rect 40640 184154 40641 184218
rect 40575 184153 40641 184154
rect 40770 183627 40830 210349
rect 40962 185995 41022 212421
rect 41151 211598 41217 211599
rect 41151 211534 41152 211598
rect 41216 211534 41217 211598
rect 41151 211533 41217 211534
rect 41154 190139 41214 211533
rect 41151 190138 41217 190139
rect 41151 190074 41152 190138
rect 41216 190074 41217 190138
rect 41151 190073 41217 190074
rect 41730 188363 41790 231661
rect 41922 231579 41982 274729
rect 42114 264879 42174 302701
rect 42495 298770 42561 298771
rect 42495 298706 42496 298770
rect 42560 298706 42561 298770
rect 42495 298705 42561 298706
rect 42303 283674 42369 283675
rect 42303 283610 42304 283674
rect 42368 283610 42369 283674
rect 42303 283609 42369 283610
rect 42306 281603 42366 283609
rect 42498 282343 42558 298705
rect 42495 282342 42561 282343
rect 42495 282278 42496 282342
rect 42560 282278 42561 282342
rect 42495 282277 42561 282278
rect 42303 281602 42369 281603
rect 42303 281538 42304 281602
rect 42368 281538 42369 281602
rect 42303 281537 42369 281538
rect 43074 274055 43134 313801
rect 43071 274054 43137 274055
rect 43071 273990 43072 274054
rect 43136 273990 43137 274054
rect 43071 273989 43137 273990
rect 287871 273906 287937 273907
rect 287871 273842 287872 273906
rect 287936 273842 287937 273906
rect 287871 273841 287937 273842
rect 284799 267838 284865 267839
rect 284799 267774 284800 267838
rect 284864 267774 284865 267838
rect 284799 267773 284865 267774
rect 284415 267542 284481 267543
rect 284415 267478 284416 267542
rect 284480 267478 284481 267542
rect 284415 267477 284481 267478
rect 284031 266062 284097 266063
rect 284031 265998 284032 266062
rect 284096 265998 284097 266062
rect 284031 265997 284097 265998
rect 42111 264878 42177 264879
rect 42111 264814 42112 264878
rect 42176 264814 42177 264878
rect 42111 264813 42177 264814
rect 204927 254962 204993 254963
rect 204927 254898 204928 254962
rect 204992 254898 204993 254962
rect 204927 254897 204993 254898
rect 204735 254814 204801 254815
rect 204735 254750 204736 254814
rect 204800 254750 204801 254814
rect 204735 254749 204801 254750
rect 145407 250670 145473 250671
rect 145407 250606 145408 250670
rect 145472 250606 145473 250670
rect 145407 250605 145473 250606
rect 42303 240754 42369 240755
rect 42303 240690 42304 240754
rect 42368 240690 42369 240754
rect 42303 240689 42369 240690
rect 42306 234835 42366 240689
rect 42303 234834 42369 234835
rect 42303 234770 42304 234834
rect 42368 234770 42369 234834
rect 42303 234769 42369 234770
rect 41919 231578 41985 231579
rect 41919 231514 41920 231578
rect 41984 231514 41985 231578
rect 41919 231513 41985 231514
rect 41922 189103 41982 231513
rect 42495 197686 42561 197687
rect 42495 197622 42496 197686
rect 42560 197622 42561 197686
rect 42495 197621 42561 197622
rect 42498 195763 42558 197621
rect 42495 195762 42561 195763
rect 42495 195698 42496 195762
rect 42560 195698 42561 195762
rect 42495 195697 42561 195698
rect 41919 189102 41985 189103
rect 41919 189038 41920 189102
rect 41984 189038 41985 189102
rect 41919 189037 41985 189038
rect 41727 188362 41793 188363
rect 41727 188298 41728 188362
rect 41792 188298 41793 188362
rect 41727 188297 41793 188298
rect 40959 185994 41025 185995
rect 40959 185930 40960 185994
rect 41024 185930 41025 185994
rect 40959 185929 41025 185930
rect 40767 183626 40833 183627
rect 40767 183562 40768 183626
rect 40832 183562 40833 183626
rect 40767 183561 40833 183562
rect 40383 182886 40449 182887
rect 40383 182822 40384 182886
rect 40448 182822 40449 182886
rect 40383 182821 40449 182822
rect 31743 177114 31809 177115
rect 31743 177050 31744 177114
rect 31808 177050 31809 177114
rect 31743 177049 31809 177050
rect 31746 125315 31806 177049
rect 31743 125314 31809 125315
rect 31743 125250 31744 125314
rect 31808 125250 31809 125314
rect 31743 125249 31809 125250
rect 145410 50871 145470 250605
rect 145599 244454 145665 244455
rect 145599 244390 145600 244454
rect 145664 244390 145665 244454
rect 145599 244389 145665 244390
rect 145602 51315 145662 244389
rect 145791 240902 145857 240903
rect 145791 240838 145792 240902
rect 145856 240838 145857 240902
rect 145791 240837 145857 240838
rect 145599 51314 145665 51315
rect 145599 51250 145600 51314
rect 145664 51250 145665 51314
rect 145599 51249 145665 51250
rect 145794 51019 145854 240837
rect 145983 236758 146049 236759
rect 145983 236694 145984 236758
rect 146048 236694 146049 236758
rect 145983 236693 146049 236694
rect 145986 51167 146046 236693
rect 204738 230247 204798 254749
rect 204930 230395 204990 254897
rect 283071 253334 283137 253335
rect 283071 253270 283072 253334
rect 283136 253270 283137 253334
rect 283071 253269 283137 253270
rect 208383 252150 208449 252151
rect 208383 252086 208384 252150
rect 208448 252086 208449 252150
rect 208383 252085 208449 252086
rect 207423 252002 207489 252003
rect 207423 251938 207424 252002
rect 207488 251938 207489 252002
rect 207423 251937 207489 251938
rect 207426 230395 207486 251937
rect 208386 230395 208446 252085
rect 283074 248895 283134 253269
rect 283071 248894 283137 248895
rect 283071 248830 283072 248894
rect 283136 248830 283137 248894
rect 283071 248829 283137 248830
rect 284034 248451 284094 265997
rect 284223 254666 284289 254667
rect 284223 254602 284224 254666
rect 284288 254602 284289 254666
rect 284223 254601 284289 254602
rect 284031 248450 284097 248451
rect 284031 248386 284032 248450
rect 284096 248386 284097 248450
rect 284031 248385 284097 248386
rect 284226 245787 284286 254601
rect 284418 246971 284478 267477
rect 284802 248599 284862 267773
rect 284991 266210 285057 266211
rect 284991 266146 284992 266210
rect 285056 266146 285057 266210
rect 284991 266145 285057 266146
rect 284799 248598 284865 248599
rect 284799 248534 284800 248598
rect 284864 248534 284865 248598
rect 284799 248533 284865 248534
rect 284799 248450 284865 248451
rect 284799 248386 284800 248450
rect 284864 248386 284865 248450
rect 284799 248385 284865 248386
rect 284802 247415 284862 248385
rect 284994 248007 285054 266145
rect 287679 264878 287745 264879
rect 287679 264814 287680 264878
rect 287744 264814 287745 264878
rect 287679 264813 287745 264814
rect 287487 262214 287553 262215
rect 287487 262150 287488 262214
rect 287552 262150 287553 262214
rect 287487 262149 287553 262150
rect 287103 256886 287169 256887
rect 287103 256822 287104 256886
rect 287168 256822 287169 256886
rect 287103 256821 287169 256822
rect 286911 256442 286977 256443
rect 286911 256378 286912 256442
rect 286976 256378 286977 256442
rect 286911 256377 286977 256378
rect 286719 256294 286785 256295
rect 286719 256230 286720 256294
rect 286784 256230 286785 256294
rect 286719 256229 286785 256230
rect 286527 253038 286593 253039
rect 286527 252974 286528 253038
rect 286592 252974 286593 253038
rect 286527 252973 286593 252974
rect 285759 248154 285825 248155
rect 285759 248090 285760 248154
rect 285824 248090 285825 248154
rect 285759 248089 285825 248090
rect 284991 248006 285057 248007
rect 284991 247942 284992 248006
rect 285056 247942 285057 248006
rect 284991 247941 285057 247942
rect 284799 247414 284865 247415
rect 284799 247350 284800 247414
rect 284864 247350 284865 247414
rect 284799 247349 284865 247350
rect 285762 247267 285822 248089
rect 285759 247266 285825 247267
rect 285759 247202 285760 247266
rect 285824 247202 285825 247266
rect 285759 247201 285825 247202
rect 284415 246970 284481 246971
rect 284415 246906 284416 246970
rect 284480 246906 284481 246970
rect 284415 246905 284481 246906
rect 284223 245786 284289 245787
rect 284223 245722 284224 245786
rect 284288 245722 284289 245786
rect 284223 245721 284289 245722
rect 286530 242235 286590 252973
rect 286527 242234 286593 242235
rect 286527 242170 286528 242234
rect 286592 242170 286593 242234
rect 286527 242169 286593 242170
rect 204927 230394 204993 230395
rect 204927 230330 204928 230394
rect 204992 230330 204993 230394
rect 204927 230329 204993 230330
rect 207423 230394 207489 230395
rect 207423 230330 207424 230394
rect 207488 230330 207489 230394
rect 207423 230329 207489 230330
rect 208383 230394 208449 230395
rect 208383 230330 208384 230394
rect 208448 230330 208449 230394
rect 208383 230329 208449 230330
rect 204735 230246 204801 230247
rect 204735 230182 204736 230246
rect 204800 230182 204801 230246
rect 204735 230181 204801 230182
rect 286722 229211 286782 256229
rect 286914 237351 286974 256377
rect 286911 237350 286977 237351
rect 286911 237286 286912 237350
rect 286976 237286 286977 237350
rect 286911 237285 286977 237286
rect 287106 232171 287166 256821
rect 287295 254518 287361 254519
rect 287295 254454 287296 254518
rect 287360 254454 287361 254518
rect 287295 254453 287361 254454
rect 287103 232170 287169 232171
rect 287103 232106 287104 232170
rect 287168 232106 287169 232170
rect 287103 232105 287169 232106
rect 286719 229210 286785 229211
rect 286719 229146 286720 229210
rect 286784 229146 286785 229210
rect 286719 229145 286785 229146
rect 287298 229063 287358 254453
rect 287490 239571 287550 262149
rect 287487 239570 287553 239571
rect 287487 239506 287488 239570
rect 287552 239506 287553 239570
rect 287487 239505 287553 239506
rect 287682 235131 287742 264813
rect 287874 238683 287934 273841
rect 442239 270650 442305 270651
rect 442239 270586 442240 270650
rect 442304 270586 442305 270650
rect 442239 270585 442305 270586
rect 450687 270650 450753 270651
rect 450687 270586 450688 270650
rect 450752 270586 450753 270650
rect 450687 270585 450753 270586
rect 442047 270058 442113 270059
rect 442047 269994 442048 270058
rect 442112 269994 442113 270058
rect 442047 269993 442113 269994
rect 290367 269022 290433 269023
rect 290367 268958 290368 269022
rect 290432 268958 290433 269022
rect 290367 268957 290433 268958
rect 290175 268874 290241 268875
rect 290175 268810 290176 268874
rect 290240 268810 290241 268874
rect 290175 268809 290241 268810
rect 289983 267690 290049 267691
rect 289983 267626 289984 267690
rect 290048 267626 290049 267690
rect 289983 267625 290049 267626
rect 289215 267246 289281 267247
rect 289215 267182 289216 267246
rect 289280 267182 289281 267246
rect 289215 267181 289281 267182
rect 289023 263398 289089 263399
rect 289023 263334 289024 263398
rect 289088 263334 289089 263398
rect 289023 263333 289089 263334
rect 288063 254074 288129 254075
rect 288063 254010 288064 254074
rect 288128 254010 288129 254074
rect 288063 254009 288129 254010
rect 287871 238682 287937 238683
rect 287871 238618 287872 238682
rect 287936 238618 287937 238682
rect 287871 238617 287937 238618
rect 287679 235130 287745 235131
rect 287679 235066 287680 235130
rect 287744 235066 287745 235130
rect 287679 235065 287745 235066
rect 287295 229062 287361 229063
rect 287295 228998 287296 229062
rect 287360 228998 287361 229062
rect 287295 228997 287361 228998
rect 288066 228915 288126 254009
rect 288255 253778 288321 253779
rect 288255 253714 288256 253778
rect 288320 253714 288321 253778
rect 288255 253713 288321 253714
rect 288258 230395 288318 253713
rect 288447 253630 288513 253631
rect 288447 253566 288448 253630
rect 288512 253566 288513 253630
rect 288447 253565 288513 253566
rect 288450 232023 288510 253565
rect 288831 253482 288897 253483
rect 288831 253418 288832 253482
rect 288896 253418 288897 253482
rect 288831 253417 288897 253418
rect 288639 253038 288705 253039
rect 288639 252974 288640 253038
rect 288704 252974 288705 253038
rect 288639 252973 288705 252974
rect 288642 248895 288702 252973
rect 288639 248894 288705 248895
rect 288639 248830 288640 248894
rect 288704 248830 288705 248894
rect 288639 248829 288705 248830
rect 288639 248746 288705 248747
rect 288639 248682 288640 248746
rect 288704 248682 288705 248746
rect 288639 248681 288705 248682
rect 288642 246675 288702 248681
rect 288639 246674 288705 246675
rect 288639 246610 288640 246674
rect 288704 246610 288705 246674
rect 288639 246609 288705 246610
rect 288639 242234 288705 242235
rect 288639 242170 288640 242234
rect 288704 242170 288705 242234
rect 288639 242169 288705 242170
rect 288642 239423 288702 242169
rect 288639 239422 288705 239423
rect 288639 239358 288640 239422
rect 288704 239358 288705 239422
rect 288639 239357 288705 239358
rect 288447 232022 288513 232023
rect 288447 231958 288448 232022
rect 288512 231958 288513 232022
rect 288447 231957 288513 231958
rect 288834 231875 288894 253417
rect 289026 235575 289086 263333
rect 289023 235574 289089 235575
rect 289023 235510 289024 235574
rect 289088 235510 289089 235574
rect 289023 235509 289089 235510
rect 289218 235427 289278 267181
rect 289791 262954 289857 262955
rect 289791 262890 289792 262954
rect 289856 262890 289857 262954
rect 289791 262889 289857 262890
rect 289599 257478 289665 257479
rect 289599 257414 289600 257478
rect 289664 257414 289665 257478
rect 289599 257413 289665 257414
rect 289407 253038 289473 253039
rect 289407 252974 289408 253038
rect 289472 252974 289473 253038
rect 289407 252973 289473 252974
rect 289410 239571 289470 252973
rect 289407 239570 289473 239571
rect 289407 239506 289408 239570
rect 289472 239506 289473 239570
rect 289407 239505 289473 239506
rect 289602 236019 289662 257413
rect 289599 236018 289665 236019
rect 289599 235954 289600 236018
rect 289664 235954 289665 236018
rect 289599 235953 289665 235954
rect 289794 235871 289854 262889
rect 289791 235870 289857 235871
rect 289791 235806 289792 235870
rect 289856 235806 289857 235870
rect 289791 235805 289857 235806
rect 289986 235723 290046 267625
rect 290178 239571 290238 268809
rect 290175 239570 290241 239571
rect 290175 239506 290176 239570
rect 290240 239506 290241 239570
rect 290175 239505 290241 239506
rect 290370 236167 290430 268957
rect 290751 268726 290817 268727
rect 290751 268662 290752 268726
rect 290816 268662 290817 268726
rect 290751 268661 290817 268662
rect 290559 268578 290625 268579
rect 290559 268514 290560 268578
rect 290624 268514 290625 268578
rect 290559 268513 290625 268514
rect 290562 239127 290622 268513
rect 290754 257479 290814 268661
rect 292863 267394 292929 267395
rect 292863 267330 292864 267394
rect 292928 267330 292929 267394
rect 292863 267329 292929 267330
rect 291519 263102 291585 263103
rect 291519 263038 291520 263102
rect 291584 263038 291585 263102
rect 291519 263037 291585 263038
rect 290751 257478 290817 257479
rect 290751 257414 290752 257478
rect 290816 257414 290817 257478
rect 290751 257413 290817 257414
rect 290751 256146 290817 256147
rect 290751 256082 290752 256146
rect 290816 256082 290817 256146
rect 290751 256081 290817 256082
rect 290754 239423 290814 256081
rect 290943 255998 291009 255999
rect 290943 255934 290944 255998
rect 291008 255934 291009 255998
rect 290943 255933 291009 255934
rect 290946 239571 291006 255933
rect 291327 255850 291393 255851
rect 291327 255786 291328 255850
rect 291392 255786 291393 255850
rect 291327 255785 291393 255786
rect 291135 253038 291201 253039
rect 291135 252974 291136 253038
rect 291200 252974 291201 253038
rect 291135 252973 291201 252974
rect 291138 239571 291198 252973
rect 291330 239571 291390 255785
rect 290943 239570 291009 239571
rect 290943 239506 290944 239570
rect 291008 239506 291009 239570
rect 290943 239505 291009 239506
rect 291135 239570 291201 239571
rect 291135 239506 291136 239570
rect 291200 239506 291201 239570
rect 291135 239505 291201 239506
rect 291327 239570 291393 239571
rect 291327 239506 291328 239570
rect 291392 239506 291393 239570
rect 291327 239505 291393 239506
rect 290751 239422 290817 239423
rect 290751 239358 290752 239422
rect 290816 239358 290817 239422
rect 290751 239357 290817 239358
rect 290559 239126 290625 239127
rect 290559 239062 290560 239126
rect 290624 239062 290625 239126
rect 290559 239061 290625 239062
rect 291522 238979 291582 263037
rect 292095 256590 292161 256591
rect 292095 256526 292096 256590
rect 292160 256526 292161 256590
rect 292095 256525 292161 256526
rect 291711 255702 291777 255703
rect 291711 255638 291712 255702
rect 291776 255638 291777 255702
rect 291711 255637 291777 255638
rect 291714 239571 291774 255637
rect 291903 255554 291969 255555
rect 291903 255490 291904 255554
rect 291968 255490 291969 255554
rect 291903 255489 291969 255490
rect 291906 239571 291966 255489
rect 291711 239570 291777 239571
rect 291711 239506 291712 239570
rect 291776 239506 291777 239570
rect 291711 239505 291777 239506
rect 291903 239570 291969 239571
rect 291903 239506 291904 239570
rect 291968 239506 291969 239570
rect 291903 239505 291969 239506
rect 291519 238978 291585 238979
rect 291519 238914 291520 238978
rect 291584 238914 291585 238978
rect 291519 238913 291585 238914
rect 292098 238239 292158 256525
rect 292287 255406 292353 255407
rect 292287 255342 292288 255406
rect 292352 255342 292353 255406
rect 292287 255341 292353 255342
rect 292290 239571 292350 255341
rect 292671 255258 292737 255259
rect 292671 255194 292672 255258
rect 292736 255194 292737 255258
rect 292671 255193 292737 255194
rect 292479 253334 292545 253335
rect 292479 253270 292480 253334
rect 292544 253270 292545 253334
rect 292479 253269 292545 253270
rect 292287 239570 292353 239571
rect 292287 239506 292288 239570
rect 292352 239506 292353 239570
rect 292287 239505 292353 239506
rect 292095 238238 292161 238239
rect 292095 238174 292096 238238
rect 292160 238174 292161 238238
rect 292095 238173 292161 238174
rect 292482 236463 292542 253269
rect 292674 239571 292734 255193
rect 292671 239570 292737 239571
rect 292671 239506 292672 239570
rect 292736 239506 292737 239570
rect 292671 239505 292737 239506
rect 292866 239275 292926 267329
rect 441471 257330 441537 257331
rect 441471 257266 441472 257330
rect 441536 257266 441537 257330
rect 441471 257265 441537 257266
rect 351423 257182 351489 257183
rect 351423 257118 351424 257182
rect 351488 257118 351489 257182
rect 351423 257117 351489 257118
rect 337215 255998 337281 255999
rect 337215 255934 337216 255998
rect 337280 255934 337281 255998
rect 337215 255933 337281 255934
rect 337218 255441 337278 255933
rect 351426 255851 351486 257117
rect 351423 255850 351489 255851
rect 351423 255786 351424 255850
rect 351488 255786 351489 255850
rect 351423 255785 351489 255786
rect 337218 255381 337662 255441
rect 293055 255110 293121 255111
rect 293055 255046 293056 255110
rect 293120 255046 293121 255110
rect 293055 255045 293121 255046
rect 293058 239571 293118 255045
rect 293247 254962 293313 254963
rect 293247 254898 293248 254962
rect 293312 254898 293313 254962
rect 293247 254897 293313 254898
rect 293055 239570 293121 239571
rect 293055 239506 293056 239570
rect 293120 239506 293121 239570
rect 293055 239505 293121 239506
rect 293250 239423 293310 254897
rect 337602 254667 337662 255381
rect 337599 254666 337665 254667
rect 337599 254602 337600 254666
rect 337664 254602 337665 254666
rect 337599 254601 337665 254602
rect 293439 254222 293505 254223
rect 293439 254158 293440 254222
rect 293504 254158 293505 254222
rect 293439 254157 293505 254158
rect 293247 239422 293313 239423
rect 293247 239358 293248 239422
rect 293312 239358 293313 239422
rect 293247 239357 293313 239358
rect 292863 239274 292929 239275
rect 292863 239210 292864 239274
rect 292928 239210 292929 239274
rect 292863 239209 292929 239210
rect 293442 237647 293502 254157
rect 441474 239568 441534 257265
rect 441855 254518 441921 254519
rect 441855 254454 441856 254518
rect 441920 254454 441921 254518
rect 441855 254453 441921 254454
rect 441663 253630 441729 253631
rect 441663 253566 441664 253630
rect 441728 253566 441729 253630
rect 441663 253565 441729 253566
rect 441282 239508 441534 239568
rect 441087 239422 441153 239423
rect 441087 239358 441088 239422
rect 441152 239358 441153 239422
rect 441087 239357 441153 239358
rect 400575 238534 400641 238535
rect 400575 238470 400576 238534
rect 400640 238470 400641 238534
rect 400575 238469 400641 238470
rect 293439 237646 293505 237647
rect 293439 237582 293440 237646
rect 293504 237582 293505 237646
rect 293439 237581 293505 237582
rect 399231 237054 399297 237055
rect 399231 236990 399232 237054
rect 399296 236990 399297 237054
rect 399231 236989 399297 236990
rect 399234 236881 399294 236989
rect 400578 236907 400638 238469
rect 400575 236906 400641 236907
rect 400575 236842 400576 236906
rect 400640 236842 400641 236906
rect 411327 236906 411393 236907
rect 411327 236881 411328 236906
rect 411392 236881 411393 236906
rect 400575 236841 400641 236842
rect 292479 236462 292545 236463
rect 292479 236398 292480 236462
rect 292544 236398 292545 236462
rect 292479 236397 292545 236398
rect 290367 236166 290433 236167
rect 290367 236102 290368 236166
rect 290432 236102 290433 236166
rect 290367 236101 290433 236102
rect 289983 235722 290049 235723
rect 289983 235658 289984 235722
rect 290048 235658 290049 235722
rect 289983 235657 290049 235658
rect 289215 235426 289281 235427
rect 289215 235362 289216 235426
rect 289280 235362 289281 235426
rect 289215 235361 289281 235362
rect 441090 234243 441150 239357
rect 441087 234242 441153 234243
rect 441087 234178 441088 234242
rect 441152 234178 441153 234242
rect 441087 234177 441153 234178
rect 288831 231874 288897 231875
rect 288831 231810 288832 231874
rect 288896 231810 288897 231874
rect 288831 231809 288897 231810
rect 288255 230394 288321 230395
rect 288255 230330 288256 230394
rect 288320 230330 288321 230394
rect 288255 230329 288321 230330
rect 288063 228914 288129 228915
rect 288063 228850 288064 228914
rect 288128 228850 288129 228914
rect 288063 228849 288129 228850
rect 413247 228174 413313 228175
rect 413247 228110 413248 228174
rect 413312 228110 413313 228174
rect 413247 228109 413313 228110
rect 207615 227730 207681 227731
rect 207615 227666 207616 227730
rect 207680 227666 207681 227730
rect 207615 227665 207681 227666
rect 207039 224030 207105 224031
rect 207039 223966 207040 224030
rect 207104 223966 207105 224030
rect 207039 223965 207105 223966
rect 206655 223882 206721 223883
rect 206655 223818 206656 223882
rect 206720 223818 206721 223882
rect 206655 223817 206721 223818
rect 206271 223734 206337 223735
rect 206271 223670 206272 223734
rect 206336 223670 206337 223734
rect 206271 223669 206337 223670
rect 206274 206823 206334 223669
rect 206274 206763 206526 206823
rect 206466 201495 206526 206763
rect 205890 201435 206526 201495
rect 205890 181515 205950 201435
rect 205890 181455 206334 181515
rect 200895 181406 200961 181407
rect 200895 181342 200896 181406
rect 200960 181342 200961 181406
rect 200895 181341 200961 181342
rect 200898 166903 200958 181341
rect 206274 168195 206334 181455
rect 206082 168135 206334 168195
rect 200895 166902 200961 166903
rect 200895 166838 200896 166902
rect 200960 166838 200961 166902
rect 200895 166837 200961 166838
rect 206082 146883 206142 168135
rect 206082 146823 206334 146883
rect 206274 126903 206334 146823
rect 206274 126843 206526 126903
rect 206466 120909 206526 126843
rect 206274 120849 206526 120909
rect 206274 90939 206334 120849
rect 206274 90879 206526 90939
rect 204351 86686 204417 86687
rect 204351 86622 204352 86686
rect 204416 86622 204417 86686
rect 204351 86621 204417 86622
rect 204159 62266 204225 62267
rect 204159 62202 204160 62266
rect 204224 62202 204225 62266
rect 204159 62201 204225 62202
rect 204162 52499 204222 62201
rect 204159 52498 204225 52499
rect 204159 52434 204160 52498
rect 204224 52434 204225 52498
rect 204159 52433 204225 52434
rect 204354 51907 204414 86621
rect 206466 86277 206526 90879
rect 205890 86217 206526 86277
rect 205890 75621 205950 86217
rect 205890 75561 206334 75621
rect 206274 65631 206334 75561
rect 206082 65571 206334 65631
rect 204735 58862 204801 58863
rect 204735 58798 204736 58862
rect 204800 58798 204801 58862
rect 204735 58797 204801 58798
rect 204738 53831 204798 58797
rect 204927 56790 204993 56791
rect 204927 56726 204928 56790
rect 204992 56726 204993 56790
rect 204927 56725 204993 56726
rect 204735 53830 204801 53831
rect 204735 53766 204736 53830
rect 204800 53766 204801 53830
rect 204735 53765 204801 53766
rect 204930 53239 204990 56725
rect 206082 54719 206142 65571
rect 206658 57639 206718 223817
rect 206847 222994 206913 222995
rect 206847 222930 206848 222994
rect 206912 222930 206913 222994
rect 206847 222929 206913 222930
rect 206274 57579 206718 57639
rect 206079 54718 206145 54719
rect 206079 54654 206080 54718
rect 206144 54654 206145 54718
rect 206079 54653 206145 54654
rect 206274 54423 206334 57579
rect 206850 56307 206910 222929
rect 206658 56247 206910 56307
rect 206271 54422 206337 54423
rect 206271 54358 206272 54422
rect 206336 54358 206337 54422
rect 206271 54357 206337 54358
rect 206658 53683 206718 56247
rect 207042 55641 207102 223965
rect 207423 223882 207489 223883
rect 207423 223818 207424 223882
rect 207488 223818 207489 223882
rect 207423 223817 207489 223818
rect 207231 222698 207297 222699
rect 207231 222634 207232 222698
rect 207296 222634 207297 222698
rect 207231 222633 207297 222634
rect 206850 55581 207102 55641
rect 206655 53682 206721 53683
rect 206655 53618 206656 53682
rect 206720 53618 206721 53682
rect 206655 53617 206721 53618
rect 204927 53238 204993 53239
rect 204927 53174 204928 53238
rect 204992 53174 204993 53238
rect 206850 53236 206910 55581
rect 207234 54975 207294 222633
rect 207042 54915 207294 54975
rect 207042 53387 207102 54915
rect 207426 54275 207486 223817
rect 207423 54274 207489 54275
rect 207423 54210 207424 54274
rect 207488 54210 207489 54274
rect 207423 54209 207489 54210
rect 207618 53979 207678 227665
rect 207999 226842 208065 226843
rect 207999 226778 208000 226842
rect 208064 226778 208065 226842
rect 207999 226777 208065 226778
rect 207807 226694 207873 226695
rect 207807 226630 207808 226694
rect 207872 226630 207873 226694
rect 207807 226629 207873 226630
rect 207615 53978 207681 53979
rect 207615 53914 207616 53978
rect 207680 53914 207681 53978
rect 207615 53913 207681 53914
rect 207810 53535 207870 226629
rect 208002 54127 208062 226777
rect 208191 226546 208257 226547
rect 208191 226482 208192 226546
rect 208256 226482 208257 226546
rect 208191 226481 208257 226482
rect 207999 54126 208065 54127
rect 207999 54062 208000 54126
rect 208064 54062 208065 54126
rect 207999 54061 208065 54062
rect 207231 53534 207297 53535
rect 207231 53470 207232 53534
rect 207296 53470 207297 53534
rect 207231 53469 207297 53470
rect 207807 53534 207873 53535
rect 207807 53470 207808 53534
rect 207872 53470 207873 53534
rect 207807 53469 207873 53470
rect 207039 53386 207105 53387
rect 207039 53322 207040 53386
rect 207104 53322 207105 53386
rect 207039 53321 207105 53322
rect 207234 53236 207294 53469
rect 206850 53176 207294 53236
rect 204927 53173 204993 53174
rect 208194 52351 208254 226481
rect 388671 224770 388737 224771
rect 388671 224706 388672 224770
rect 388736 224706 388737 224770
rect 388671 224705 388737 224706
rect 391743 224770 391809 224771
rect 391743 224706 391744 224770
rect 391808 224706 391809 224770
rect 391743 224705 391809 224706
rect 388674 223883 388734 224705
rect 391746 223883 391806 224705
rect 400191 224030 400257 224031
rect 400191 223966 400192 224030
rect 400256 223966 400257 224030
rect 400191 223965 400257 223966
rect 349311 223882 349377 223883
rect 349311 223818 349312 223882
rect 349376 223818 349377 223882
rect 349311 223817 349377 223818
rect 359679 223882 359745 223883
rect 359679 223818 359680 223882
rect 359744 223818 359745 223882
rect 359679 223817 359745 223818
rect 362751 223882 362817 223883
rect 362751 223818 362752 223882
rect 362816 223818 362817 223882
rect 362751 223817 362817 223818
rect 388671 223882 388737 223883
rect 388671 223818 388672 223882
rect 388736 223818 388737 223882
rect 388671 223817 388737 223818
rect 391743 223882 391809 223883
rect 391743 223818 391744 223882
rect 391808 223818 391809 223882
rect 391743 223817 391809 223818
rect 302463 223586 302529 223587
rect 302463 223522 302464 223586
rect 302528 223522 302529 223586
rect 302463 223521 302529 223522
rect 302466 223143 302526 223521
rect 302463 223142 302529 223143
rect 302463 223078 302464 223142
rect 302528 223078 302529 223142
rect 302463 223077 302529 223078
rect 349314 222699 349374 223817
rect 359682 222995 359742 223817
rect 359679 222994 359745 222995
rect 359679 222930 359680 222994
rect 359744 222930 359745 222994
rect 359679 222929 359745 222930
rect 362754 222847 362814 223817
rect 380031 223586 380097 223587
rect 380031 223522 380032 223586
rect 380096 223522 380097 223586
rect 380031 223521 380097 223522
rect 380034 223143 380094 223521
rect 400194 223439 400254 223965
rect 405567 223882 405633 223883
rect 405567 223818 405568 223882
rect 405632 223880 405633 223882
rect 405951 223882 406017 223883
rect 405951 223880 405952 223882
rect 405632 223820 405952 223880
rect 405632 223818 405633 223820
rect 405567 223817 405633 223818
rect 405951 223818 405952 223820
rect 406016 223818 406017 223882
rect 405951 223817 406017 223818
rect 413250 223735 413310 228109
rect 441282 228027 441342 239508
rect 441666 237351 441726 253565
rect 441663 237350 441729 237351
rect 441663 237286 441664 237350
rect 441728 237286 441729 237350
rect 441663 237285 441729 237286
rect 441858 230395 441918 254453
rect 442050 238831 442110 269993
rect 442242 238979 442302 270585
rect 446463 270502 446529 270503
rect 446463 270438 446464 270502
rect 446528 270438 446529 270502
rect 446463 270437 446529 270438
rect 449535 270502 449601 270503
rect 449535 270438 449536 270502
rect 449600 270438 449601 270502
rect 449535 270437 449601 270438
rect 443583 270354 443649 270355
rect 443583 270290 443584 270354
rect 443648 270290 443649 270354
rect 443583 270289 443649 270290
rect 443007 270206 443073 270207
rect 443007 270142 443008 270206
rect 443072 270142 443073 270206
rect 443007 270141 443073 270142
rect 442623 258958 442689 258959
rect 442623 258894 442624 258958
rect 442688 258894 442689 258958
rect 442623 258893 442689 258894
rect 442431 254370 442497 254371
rect 442431 254306 442432 254370
rect 442496 254306 442497 254370
rect 442431 254305 442497 254306
rect 442434 239423 442494 254305
rect 442626 253631 442686 258893
rect 442815 258810 442881 258811
rect 442815 258746 442816 258810
rect 442880 258746 442881 258810
rect 442815 258745 442881 258746
rect 442623 253630 442689 253631
rect 442623 253566 442624 253630
rect 442688 253566 442689 253630
rect 442623 253565 442689 253566
rect 442623 253038 442689 253039
rect 442623 252974 442624 253038
rect 442688 252974 442689 253038
rect 442623 252973 442689 252974
rect 442626 239571 442686 252973
rect 442818 246117 442878 258745
rect 443010 256147 443070 270141
rect 443391 268282 443457 268283
rect 443391 268218 443392 268282
rect 443456 268218 443457 268282
rect 443391 268217 443457 268218
rect 443199 259106 443265 259107
rect 443199 259042 443200 259106
rect 443264 259042 443265 259106
rect 443199 259041 443265 259042
rect 443007 256146 443073 256147
rect 443007 256082 443008 256146
rect 443072 256082 443073 256146
rect 443007 256081 443073 256082
rect 442818 246057 443070 246117
rect 442623 239570 442689 239571
rect 442623 239506 442624 239570
rect 442688 239506 442689 239570
rect 442623 239505 442689 239506
rect 442431 239422 442497 239423
rect 442431 239358 442432 239422
rect 442496 239358 442497 239422
rect 442431 239357 442497 239358
rect 442239 238978 442305 238979
rect 442239 238914 442240 238978
rect 442304 238914 442305 238978
rect 442239 238913 442305 238914
rect 442431 238978 442497 238979
rect 442431 238914 442432 238978
rect 442496 238914 442497 238978
rect 442431 238913 442497 238914
rect 442047 238830 442113 238831
rect 442047 238766 442048 238830
rect 442112 238766 442113 238830
rect 442047 238765 442113 238766
rect 442434 236759 442494 238913
rect 442623 238830 442689 238831
rect 442623 238766 442624 238830
rect 442688 238766 442689 238830
rect 442623 238765 442689 238766
rect 442431 236758 442497 236759
rect 442431 236694 442432 236758
rect 442496 236694 442497 236758
rect 442431 236693 442497 236694
rect 442626 230839 442686 238765
rect 442815 237350 442881 237351
rect 442815 237286 442816 237350
rect 442880 237286 442881 237350
rect 442815 237285 442881 237286
rect 442818 233651 442878 237285
rect 442815 233650 442881 233651
rect 442815 233586 442816 233650
rect 442880 233586 442881 233650
rect 442815 233585 442881 233586
rect 443010 233503 443070 246057
rect 443007 233502 443073 233503
rect 443007 233438 443008 233502
rect 443072 233438 443073 233502
rect 443007 233437 443073 233438
rect 442623 230838 442689 230839
rect 442623 230774 442624 230838
rect 442688 230774 442689 230838
rect 442623 230773 442689 230774
rect 441855 230394 441921 230395
rect 441855 230330 441856 230394
rect 441920 230330 441921 230394
rect 441855 230329 441921 230330
rect 441279 228026 441345 228027
rect 441279 227962 441280 228026
rect 441344 227962 441345 228026
rect 441279 227961 441345 227962
rect 443202 227435 443262 259041
rect 443394 232171 443454 268217
rect 443586 258105 443646 270289
rect 445695 269466 445761 269467
rect 445695 269402 445696 269466
rect 445760 269402 445761 269466
rect 445695 269401 445761 269402
rect 443586 258045 445566 258105
rect 445119 257034 445185 257035
rect 445119 256970 445120 257034
rect 445184 256970 445185 257034
rect 445119 256969 445185 256970
rect 443775 256738 443841 256739
rect 443775 256674 443776 256738
rect 443840 256674 443841 256738
rect 443775 256673 443841 256674
rect 443583 253038 443649 253039
rect 443583 252974 443584 253038
rect 443648 252974 443649 253038
rect 443583 252973 443649 252974
rect 443586 239275 443646 252973
rect 443583 239274 443649 239275
rect 443583 239210 443584 239274
rect 443648 239210 443649 239274
rect 443583 239209 443649 239210
rect 443583 236166 443649 236167
rect 443583 236102 443584 236166
rect 443648 236102 443649 236166
rect 443583 236101 443649 236102
rect 443391 232170 443457 232171
rect 443391 232106 443392 232170
rect 443456 232106 443457 232170
rect 443391 232105 443457 232106
rect 443586 230395 443646 236101
rect 443583 230394 443649 230395
rect 443583 230330 443584 230394
rect 443648 230330 443649 230394
rect 443583 230329 443649 230330
rect 443778 227879 443838 256673
rect 444159 254518 444225 254519
rect 444159 254454 444160 254518
rect 444224 254454 444225 254518
rect 444159 254453 444225 254454
rect 443967 254074 444033 254075
rect 443967 254010 443968 254074
rect 444032 254010 444033 254074
rect 443967 254009 444033 254010
rect 443970 239423 444030 254009
rect 443967 239422 444033 239423
rect 443967 239358 443968 239422
rect 444032 239358 444033 239422
rect 443967 239357 444033 239358
rect 444162 239275 444222 254453
rect 444351 254370 444417 254371
rect 444351 254306 444352 254370
rect 444416 254306 444417 254370
rect 444351 254305 444417 254306
rect 444354 239423 444414 254305
rect 444543 254222 444609 254223
rect 444543 254158 444544 254222
rect 444608 254158 444609 254222
rect 444543 254157 444609 254158
rect 444351 239422 444417 239423
rect 444351 239358 444352 239422
rect 444416 239358 444417 239422
rect 444351 239357 444417 239358
rect 444159 239274 444225 239275
rect 444159 239210 444160 239274
rect 444224 239210 444225 239274
rect 444159 239209 444225 239210
rect 444546 237499 444606 254157
rect 444927 253482 444993 253483
rect 444927 253418 444928 253482
rect 444992 253418 444993 253482
rect 444927 253417 444993 253418
rect 444735 253334 444801 253335
rect 444735 253270 444736 253334
rect 444800 253270 444801 253334
rect 444735 253269 444801 253270
rect 444543 237498 444609 237499
rect 444543 237434 444544 237498
rect 444608 237434 444609 237498
rect 444543 237433 444609 237434
rect 444738 236907 444798 253269
rect 444735 236906 444801 236907
rect 444735 236842 444736 236906
rect 444800 236842 444801 236906
rect 444735 236841 444801 236842
rect 444930 236611 444990 253417
rect 445122 239275 445182 256969
rect 445311 256886 445377 256887
rect 445311 256822 445312 256886
rect 445376 256822 445377 256886
rect 445311 256821 445377 256822
rect 445314 239423 445374 256821
rect 445311 239422 445377 239423
rect 445311 239358 445312 239422
rect 445376 239358 445377 239422
rect 445311 239357 445377 239358
rect 445119 239274 445185 239275
rect 445119 239210 445120 239274
rect 445184 239210 445185 239274
rect 445119 239209 445185 239210
rect 445506 237943 445566 258045
rect 445698 238387 445758 269401
rect 446079 258366 446145 258367
rect 446079 258302 446080 258366
rect 446144 258302 446145 258366
rect 446079 258301 446145 258302
rect 445887 253630 445953 253631
rect 445887 253566 445888 253630
rect 445952 253566 445953 253630
rect 445887 253565 445953 253566
rect 445890 238979 445950 253565
rect 445887 238978 445953 238979
rect 445887 238914 445888 238978
rect 445952 238914 445953 238978
rect 445887 238913 445953 238914
rect 445695 238386 445761 238387
rect 445695 238322 445696 238386
rect 445760 238322 445761 238386
rect 445695 238321 445761 238322
rect 445503 237942 445569 237943
rect 445503 237878 445504 237942
rect 445568 237878 445569 237942
rect 445503 237877 445569 237878
rect 446082 237055 446142 258301
rect 446271 253038 446337 253039
rect 446271 252974 446272 253038
rect 446336 252974 446337 253038
rect 446271 252973 446337 252974
rect 446274 239571 446334 252973
rect 446271 239570 446337 239571
rect 446271 239506 446272 239570
rect 446336 239506 446337 239570
rect 446271 239505 446337 239506
rect 446079 237054 446145 237055
rect 446079 236990 446080 237054
rect 446144 236990 446145 237054
rect 446079 236989 446145 236990
rect 444927 236610 444993 236611
rect 444927 236546 444928 236610
rect 444992 236546 444993 236610
rect 444927 236545 444993 236546
rect 446079 232762 446145 232763
rect 446079 232698 446080 232762
rect 446144 232698 446145 232762
rect 446079 232697 446145 232698
rect 443775 227878 443841 227879
rect 443775 227814 443776 227878
rect 443840 227814 443841 227878
rect 443775 227813 443841 227814
rect 443199 227434 443265 227435
rect 443199 227370 443200 227434
rect 443264 227370 443265 227434
rect 443199 227369 443265 227370
rect 419199 226990 419265 226991
rect 419199 226926 419200 226990
rect 419264 226926 419265 226990
rect 419199 226925 419265 226926
rect 419202 226695 419262 226925
rect 419007 226694 419073 226695
rect 419007 226630 419008 226694
rect 419072 226630 419073 226694
rect 419007 226629 419073 226630
rect 419199 226694 419265 226695
rect 419199 226630 419200 226694
rect 419264 226630 419265 226694
rect 419199 226629 419265 226630
rect 419010 226137 419070 226629
rect 419010 226077 419262 226137
rect 419202 225807 419262 226077
rect 419199 225806 419265 225807
rect 419199 225742 419200 225806
rect 419264 225742 419265 225806
rect 419199 225741 419265 225742
rect 428994 224745 429438 224805
rect 428994 223735 429054 224745
rect 429378 224327 429438 224745
rect 429183 224326 429249 224327
rect 429183 224262 429184 224326
rect 429248 224262 429249 224326
rect 429183 224261 429249 224262
rect 429375 224326 429441 224327
rect 429375 224262 429376 224326
rect 429440 224262 429441 224326
rect 429375 224261 429441 224262
rect 413055 223734 413121 223735
rect 413055 223670 413056 223734
rect 413120 223670 413121 223734
rect 413055 223669 413121 223670
rect 413247 223734 413313 223735
rect 413247 223670 413248 223734
rect 413312 223670 413313 223734
rect 413247 223669 413313 223670
rect 428991 223734 429057 223735
rect 428991 223670 428992 223734
rect 429056 223670 429057 223734
rect 428991 223669 429057 223670
rect 400191 223438 400257 223439
rect 400191 223374 400192 223438
rect 400256 223374 400257 223438
rect 400191 223373 400257 223374
rect 413058 223291 413118 223669
rect 429186 223473 429246 224261
rect 439551 224030 439617 224031
rect 439551 223966 439552 224030
rect 439616 223966 439617 224030
rect 439551 223965 439617 223966
rect 440127 224030 440193 224031
rect 440127 223966 440128 224030
rect 440192 223966 440193 224030
rect 440127 223965 440193 223966
rect 440895 224030 440961 224031
rect 440895 223966 440896 224030
rect 440960 223966 440961 224030
rect 440895 223965 440961 223966
rect 429567 223882 429633 223883
rect 429567 223818 429568 223882
rect 429632 223818 429633 223882
rect 429567 223817 429633 223818
rect 429570 223587 429630 223817
rect 429567 223586 429633 223587
rect 429567 223522 429568 223586
rect 429632 223522 429633 223586
rect 429567 223521 429633 223522
rect 429186 223439 429438 223473
rect 429186 223438 429441 223439
rect 429186 223413 429376 223438
rect 429375 223374 429376 223413
rect 429440 223374 429441 223438
rect 429375 223373 429441 223374
rect 413055 223290 413121 223291
rect 413055 223226 413056 223290
rect 413120 223226 413121 223290
rect 413055 223225 413121 223226
rect 417471 223290 417537 223291
rect 417471 223226 417472 223290
rect 417536 223288 417537 223290
rect 417663 223290 417729 223291
rect 417663 223288 417664 223290
rect 417536 223228 417664 223288
rect 417536 223226 417537 223228
rect 417471 223225 417537 223226
rect 417663 223226 417664 223228
rect 417728 223226 417729 223290
rect 417663 223225 417729 223226
rect 380031 223142 380097 223143
rect 380031 223078 380032 223142
rect 380096 223078 380097 223142
rect 380031 223077 380097 223078
rect 380271 223142 380337 223143
rect 380271 223078 380272 223142
rect 380336 223140 380337 223142
rect 400191 223142 400257 223143
rect 380336 223080 380478 223140
rect 380336 223078 380337 223080
rect 380271 223077 380337 223078
rect 380418 222895 380478 223080
rect 400191 223078 400192 223142
rect 400256 223078 400257 223142
rect 400191 223077 400257 223078
rect 400194 222895 400254 223077
rect 439554 222995 439614 223965
rect 439551 222994 439617 222995
rect 439551 222930 439552 222994
rect 439616 222930 439617 222994
rect 439551 222929 439617 222930
rect 362751 222846 362817 222847
rect 362751 222782 362752 222846
rect 362816 222782 362817 222846
rect 362751 222781 362817 222782
rect 349311 222698 349377 222699
rect 349311 222634 349312 222698
rect 349376 222634 349377 222698
rect 440130 222847 440190 223965
rect 440127 222846 440193 222847
rect 440127 222782 440128 222846
rect 440192 222782 440193 222846
rect 440127 222781 440193 222782
rect 440898 222699 440958 223965
rect 446082 223291 446142 232697
rect 446466 223439 446526 270437
rect 447231 269022 447297 269023
rect 447231 268958 447232 269022
rect 447296 268958 447297 269022
rect 447231 268957 447297 268958
rect 446655 268134 446721 268135
rect 446655 268070 446656 268134
rect 446720 268070 446721 268134
rect 446655 268069 446721 268070
rect 446658 259437 446718 268069
rect 446658 259377 447102 259437
rect 446847 258662 446913 258663
rect 446847 258598 446848 258662
rect 446912 258598 446913 258662
rect 446847 258597 446913 258598
rect 446655 255998 446721 255999
rect 446655 255934 446656 255998
rect 446720 255934 446721 255998
rect 446655 255933 446721 255934
rect 446658 237647 446718 255933
rect 446655 237646 446721 237647
rect 446655 237582 446656 237646
rect 446720 237582 446721 237646
rect 446655 237581 446721 237582
rect 446850 226399 446910 258597
rect 447042 238683 447102 259377
rect 447039 238682 447105 238683
rect 447039 238618 447040 238682
rect 447104 238618 447105 238682
rect 447039 238617 447105 238618
rect 447234 238535 447294 268957
rect 449343 268430 449409 268431
rect 449343 268366 449344 268430
rect 449408 268366 449409 268430
rect 449343 268365 449409 268366
rect 448383 257182 448449 257183
rect 448383 257118 448384 257182
rect 448448 257118 448449 257182
rect 448383 257117 448449 257118
rect 447807 256590 447873 256591
rect 447807 256526 447808 256590
rect 447872 256526 447873 256590
rect 447807 256525 447873 256526
rect 447615 254370 447681 254371
rect 447615 254306 447616 254370
rect 447680 254306 447681 254370
rect 447615 254305 447681 254306
rect 447423 253038 447489 253039
rect 447423 252974 447424 253038
rect 447488 252974 447489 253038
rect 447423 252973 447489 252974
rect 447231 238534 447297 238535
rect 447231 238470 447232 238534
rect 447296 238470 447297 238534
rect 447231 238469 447297 238470
rect 447231 237646 447297 237647
rect 447231 237582 447232 237646
rect 447296 237582 447297 237646
rect 447231 237581 447297 237582
rect 446847 226398 446913 226399
rect 446847 226334 446848 226398
rect 446912 226334 446913 226398
rect 446847 226333 446913 226334
rect 447234 224919 447294 237581
rect 447426 225659 447486 252973
rect 447618 239275 447678 254305
rect 447810 239423 447870 256525
rect 448191 255554 448257 255555
rect 448191 255490 448192 255554
rect 448256 255490 448257 255554
rect 448191 255489 448257 255490
rect 447999 254222 448065 254223
rect 447999 254158 448000 254222
rect 448064 254158 448065 254222
rect 447999 254157 448065 254158
rect 447807 239422 447873 239423
rect 447807 239358 447808 239422
rect 447872 239358 447873 239422
rect 447807 239357 447873 239358
rect 447615 239274 447681 239275
rect 447615 239210 447616 239274
rect 447680 239210 447681 239274
rect 447615 239209 447681 239210
rect 448002 233799 448062 254157
rect 448194 237647 448254 255489
rect 448191 237646 448257 237647
rect 448191 237582 448192 237646
rect 448256 237582 448257 237646
rect 448191 237581 448257 237582
rect 447999 233798 448065 233799
rect 447999 233734 448000 233798
rect 448064 233734 448065 233798
rect 447999 233733 448065 233734
rect 448386 226695 448446 257117
rect 448767 256294 448833 256295
rect 448767 256230 448768 256294
rect 448832 256230 448833 256294
rect 448767 256229 448833 256230
rect 448575 255850 448641 255851
rect 448575 255786 448576 255850
rect 448640 255786 448641 255850
rect 448575 255785 448641 255786
rect 448383 226694 448449 226695
rect 448383 226630 448384 226694
rect 448448 226630 448449 226694
rect 448383 226629 448449 226630
rect 447423 225658 447489 225659
rect 447423 225594 447424 225658
rect 447488 225594 447489 225658
rect 447423 225593 447489 225594
rect 447231 224918 447297 224919
rect 447231 224854 447232 224918
rect 447296 224854 447297 224918
rect 447231 224853 447297 224854
rect 448578 224771 448638 255785
rect 448770 239275 448830 256229
rect 448959 256146 449025 256147
rect 448959 256082 448960 256146
rect 449024 256082 449025 256146
rect 448959 256081 449025 256082
rect 448767 239274 448833 239275
rect 448767 239210 448768 239274
rect 448832 239210 448833 239274
rect 448767 239209 448833 239210
rect 448962 238831 449022 256081
rect 449346 252111 449406 268365
rect 449538 252777 449598 270437
rect 449727 269762 449793 269763
rect 449727 269698 449728 269762
rect 449792 269698 449793 269762
rect 449727 269697 449793 269698
rect 449730 254960 449790 269697
rect 449730 254900 450366 254960
rect 449919 254814 449985 254815
rect 449919 254750 449920 254814
rect 449984 254750 449985 254814
rect 449919 254749 449985 254750
rect 449538 252717 449790 252777
rect 449346 252051 449598 252111
rect 448959 238830 449025 238831
rect 448959 238766 448960 238830
rect 449024 238766 449025 238830
rect 448959 238765 449025 238766
rect 448575 224770 448641 224771
rect 448575 224706 448576 224770
rect 448640 224706 448641 224770
rect 448575 224705 448641 224706
rect 449538 223883 449598 252051
rect 449730 225215 449790 252717
rect 449922 237203 449982 254749
rect 450111 253482 450177 253483
rect 450111 253418 450112 253482
rect 450176 253418 450177 253482
rect 450111 253417 450177 253418
rect 450114 239423 450174 253417
rect 450111 239422 450177 239423
rect 450111 239358 450112 239422
rect 450176 239358 450177 239422
rect 450111 239357 450177 239358
rect 450306 239127 450366 254900
rect 450495 253334 450561 253335
rect 450495 253270 450496 253334
rect 450560 253270 450561 253334
rect 450495 253269 450561 253270
rect 450303 239126 450369 239127
rect 450303 239062 450304 239126
rect 450368 239062 450369 239126
rect 450303 239061 450369 239062
rect 449919 237202 449985 237203
rect 449919 237138 449920 237202
rect 449984 237138 449985 237202
rect 449919 237137 449985 237138
rect 449727 225214 449793 225215
rect 449727 225150 449728 225214
rect 449792 225150 449793 225214
rect 449727 225149 449793 225150
rect 449535 223882 449601 223883
rect 449535 223818 449536 223882
rect 449600 223818 449601 223882
rect 449535 223817 449601 223818
rect 450498 223587 450558 253269
rect 450690 237795 450750 270585
rect 673986 269911 674046 314837
rect 674178 272279 674238 316391
rect 674946 315939 675006 345473
rect 675138 330591 675198 351393
rect 675522 335179 675582 374481
rect 675711 371586 675777 371587
rect 675711 371522 675712 371586
rect 675776 371522 675777 371586
rect 675711 371521 675777 371522
rect 675519 335178 675585 335179
rect 675519 335114 675520 335178
rect 675584 335114 675585 335178
rect 675519 335113 675585 335114
rect 675714 334029 675774 371521
rect 675903 360190 675969 360191
rect 675903 360126 675904 360190
rect 675968 360126 675969 360190
rect 675903 360125 675969 360126
rect 675330 333969 675774 334029
rect 675330 333847 675390 333969
rect 675327 333846 675393 333847
rect 675327 333782 675328 333846
rect 675392 333782 675393 333846
rect 675327 333781 675393 333782
rect 675135 330590 675201 330591
rect 675135 330526 675136 330590
rect 675200 330526 675201 330590
rect 675135 330525 675201 330526
rect 674943 315938 675009 315939
rect 674943 315874 674944 315938
rect 675008 315874 675009 315938
rect 674943 315873 675009 315874
rect 674367 315790 674433 315791
rect 674367 315726 674368 315790
rect 674432 315726 674433 315790
rect 674367 315725 674433 315726
rect 674175 272278 674241 272279
rect 674175 272214 674176 272278
rect 674240 272214 674241 272278
rect 674175 272213 674241 272214
rect 674370 270799 674430 315725
rect 674751 312682 674817 312683
rect 674751 312618 674752 312682
rect 674816 312618 674817 312682
rect 674751 312617 674817 312618
rect 674559 309574 674625 309575
rect 674559 309510 674560 309574
rect 674624 309510 674625 309574
rect 674559 309509 674625 309510
rect 674562 281899 674622 309509
rect 674754 283675 674814 312617
rect 674943 306466 675009 306467
rect 674943 306402 674944 306466
rect 675008 306402 675009 306466
rect 674943 306401 675009 306402
rect 674946 285303 675006 306401
rect 675330 289595 675390 333781
rect 675519 329554 675585 329555
rect 675519 329490 675520 329554
rect 675584 329490 675585 329554
rect 675519 329489 675585 329490
rect 675522 290187 675582 329489
rect 675906 315199 675966 360125
rect 675903 315198 675969 315199
rect 675903 315134 675904 315198
rect 675968 315134 675969 315198
rect 675903 315133 675969 315134
rect 675519 290186 675585 290187
rect 675519 290122 675520 290186
rect 675584 290122 675585 290186
rect 675519 290121 675585 290122
rect 675327 289594 675393 289595
rect 675327 289530 675328 289594
rect 675392 289530 675393 289594
rect 675327 289529 675393 289530
rect 674943 285302 675009 285303
rect 674943 285238 674944 285302
rect 675008 285238 675009 285302
rect 674943 285237 675009 285238
rect 674751 283674 674817 283675
rect 674751 283610 674752 283674
rect 674816 283610 674817 283674
rect 674751 283609 674817 283610
rect 674751 282342 674817 282343
rect 674751 282278 674752 282342
rect 674816 282278 674817 282342
rect 674751 282277 674817 282278
rect 674559 281898 674625 281899
rect 674559 281834 674560 281898
rect 674624 281834 674625 281898
rect 674559 281833 674625 281834
rect 674754 273611 674814 282277
rect 674751 273610 674817 273611
rect 674751 273546 674752 273610
rect 674816 273546 674817 273610
rect 674751 273545 674817 273546
rect 674943 273610 675009 273611
rect 674943 273546 674944 273610
rect 675008 273546 675009 273610
rect 674943 273545 675009 273546
rect 674754 272723 674814 273545
rect 674751 272722 674817 272723
rect 674751 272658 674752 272722
rect 674816 272658 674817 272722
rect 674751 272657 674817 272658
rect 674367 270798 674433 270799
rect 674367 270734 674368 270798
rect 674432 270734 674433 270798
rect 674367 270733 674433 270734
rect 673983 269910 674049 269911
rect 673983 269846 673984 269910
rect 674048 269846 674049 269910
rect 673983 269845 674049 269846
rect 452223 269318 452289 269319
rect 452223 269254 452224 269318
rect 452288 269254 452289 269318
rect 452223 269253 452289 269254
rect 451071 258514 451137 258515
rect 451071 258450 451072 258514
rect 451136 258450 451137 258514
rect 451071 258449 451137 258450
rect 450879 253186 450945 253187
rect 450879 253122 450880 253186
rect 450944 253122 450945 253186
rect 450879 253121 450945 253122
rect 450687 237794 450753 237795
rect 450687 237730 450688 237794
rect 450752 237730 450753 237794
rect 450687 237729 450753 237730
rect 450882 232763 450942 253121
rect 450879 232762 450945 232763
rect 450879 232698 450880 232762
rect 450944 232698 450945 232762
rect 450879 232697 450945 232698
rect 451074 225511 451134 258449
rect 451263 254074 451329 254075
rect 451263 254010 451264 254074
rect 451328 254010 451329 254074
rect 451263 254009 451329 254010
rect 451266 233947 451326 254009
rect 451263 233946 451329 233947
rect 451263 233882 451264 233946
rect 451328 233882 451329 233946
rect 451263 233881 451329 233882
rect 452226 227287 452286 269253
rect 452415 269170 452481 269171
rect 452415 269106 452416 269170
rect 452480 269106 452481 269170
rect 452415 269105 452481 269106
rect 452223 227286 452289 227287
rect 452223 227222 452224 227286
rect 452288 227222 452289 227286
rect 452223 227221 452289 227222
rect 452418 226547 452478 269105
rect 673986 255703 674046 269845
rect 674751 268578 674817 268579
rect 674751 268514 674752 268578
rect 674816 268514 674817 268578
rect 674751 268513 674817 268514
rect 674559 265470 674625 265471
rect 674559 265406 674560 265470
rect 674624 265406 674625 265470
rect 674559 265405 674625 265406
rect 674367 265174 674433 265175
rect 674367 265110 674368 265174
rect 674432 265110 674433 265174
rect 674367 265109 674433 265110
rect 452991 255702 453057 255703
rect 452991 255638 452992 255702
rect 453056 255638 453057 255702
rect 452991 255637 453057 255638
rect 673983 255702 674049 255703
rect 673983 255638 673984 255702
rect 674048 255638 674049 255702
rect 673983 255637 674049 255638
rect 452607 253926 452673 253927
rect 452607 253862 452608 253926
rect 452672 253862 452673 253926
rect 452607 253861 452673 253862
rect 452415 226546 452481 226547
rect 452415 226482 452416 226546
rect 452480 226482 452481 226546
rect 452415 226481 452481 226482
rect 451071 225510 451137 225511
rect 451071 225446 451072 225510
rect 451136 225446 451137 225510
rect 451071 225445 451137 225446
rect 452610 225363 452670 253861
rect 452799 253778 452865 253779
rect 452799 253714 452800 253778
rect 452864 253714 452865 253778
rect 452799 253713 452865 253714
rect 452802 226399 452862 253713
rect 452994 226843 453054 255637
rect 453759 255406 453825 255407
rect 453759 255342 453760 255406
rect 453824 255342 453825 255406
rect 453759 255341 453825 255342
rect 453183 255258 453249 255259
rect 453183 255194 453184 255258
rect 453248 255194 453249 255258
rect 453183 255193 453249 255194
rect 453186 227139 453246 255193
rect 453375 255110 453441 255111
rect 453375 255046 453376 255110
rect 453440 255046 453441 255110
rect 453375 255045 453441 255046
rect 453183 227138 453249 227139
rect 453183 227074 453184 227138
rect 453248 227074 453249 227138
rect 453183 227073 453249 227074
rect 452991 226842 453057 226843
rect 452991 226778 452992 226842
rect 453056 226778 453057 226842
rect 452991 226777 453057 226778
rect 452799 226398 452865 226399
rect 452799 226334 452800 226398
rect 452864 226334 452865 226398
rect 452799 226333 452865 226334
rect 453378 226251 453438 255045
rect 453567 253038 453633 253039
rect 453567 252974 453568 253038
rect 453632 252974 453633 253038
rect 453567 252973 453633 252974
rect 453375 226250 453441 226251
rect 453375 226186 453376 226250
rect 453440 226186 453441 226250
rect 453375 226185 453441 226186
rect 453570 226103 453630 252973
rect 453567 226102 453633 226103
rect 453567 226038 453568 226102
rect 453632 226038 453633 226102
rect 453567 226037 453633 226038
rect 452607 225362 452673 225363
rect 452607 225298 452608 225362
rect 452672 225298 452673 225362
rect 452607 225297 452673 225298
rect 453762 225067 453822 255341
rect 454143 254962 454209 254963
rect 454143 254898 454144 254962
rect 454208 254898 454209 254962
rect 454143 254897 454209 254898
rect 453951 254666 454017 254667
rect 453951 254602 453952 254666
rect 454016 254602 454017 254666
rect 453951 254601 454017 254602
rect 453954 226991 454014 254601
rect 453951 226990 454017 226991
rect 453951 226926 453952 226990
rect 454016 226926 454017 226990
rect 453951 226925 454017 226926
rect 454146 225807 454206 254897
rect 454143 225806 454209 225807
rect 454143 225742 454144 225806
rect 454208 225742 454209 225806
rect 454143 225741 454209 225742
rect 453759 225066 453825 225067
rect 453759 225002 453760 225066
rect 453824 225002 453825 225066
rect 453759 225001 453825 225002
rect 673986 224771 674046 255637
rect 674370 236907 674430 265109
rect 674562 243567 674622 265405
rect 674754 249635 674814 268513
rect 674946 257331 675006 273545
rect 675903 270946 675969 270947
rect 675903 270882 675904 270946
rect 675968 270882 675969 270946
rect 675903 270881 675969 270882
rect 675711 268134 675777 268135
rect 675711 268070 675712 268134
rect 675776 268070 675777 268134
rect 675711 268069 675777 268070
rect 675327 262214 675393 262215
rect 675327 262150 675328 262214
rect 675392 262150 675393 262214
rect 675327 262149 675393 262150
rect 674943 257330 675009 257331
rect 674943 257266 674944 257330
rect 675008 257266 675009 257330
rect 674943 257265 675009 257266
rect 674751 249634 674817 249635
rect 674751 249570 674752 249634
rect 674816 249570 674817 249634
rect 674751 249569 674817 249570
rect 675330 245047 675390 262149
rect 675519 257330 675585 257331
rect 675519 257266 675520 257330
rect 675584 257266 675585 257330
rect 675519 257265 675585 257266
rect 674943 245046 675009 245047
rect 674943 244982 674944 245046
rect 675008 244982 675009 245046
rect 674943 244981 675009 244982
rect 675327 245046 675393 245047
rect 675327 244982 675328 245046
rect 675392 244982 675393 245046
rect 675327 244981 675393 244982
rect 674559 243566 674625 243567
rect 674559 243502 674560 243566
rect 674624 243502 674625 243566
rect 674559 243501 674625 243502
rect 674751 238978 674817 238979
rect 674751 238914 674752 238978
rect 674816 238914 674817 238978
rect 674751 238913 674817 238914
rect 674367 236906 674433 236907
rect 674367 236842 674368 236906
rect 674432 236842 674433 236906
rect 674367 236841 674433 236842
rect 674175 226250 674241 226251
rect 674175 226186 674176 226250
rect 674240 226186 674241 226250
rect 674175 226185 674241 226186
rect 673983 224770 674049 224771
rect 673983 224706 673984 224770
rect 674048 224706 674049 224770
rect 673983 224705 674049 224706
rect 633471 224178 633537 224179
rect 633471 224114 633472 224178
rect 633536 224114 633537 224178
rect 633471 224113 633537 224114
rect 632511 224030 632577 224031
rect 632511 223966 632512 224030
rect 632576 223966 632577 224030
rect 632511 223965 632577 223966
rect 632703 224030 632769 224031
rect 632703 223966 632704 224030
rect 632768 223966 632769 224030
rect 632703 223965 632769 223966
rect 632127 223882 632193 223883
rect 632127 223818 632128 223882
rect 632192 223818 632193 223882
rect 632127 223817 632193 223818
rect 632319 223882 632385 223883
rect 632319 223818 632320 223882
rect 632384 223818 632385 223882
rect 632319 223817 632385 223818
rect 450495 223586 450561 223587
rect 446463 223438 446529 223439
rect 446463 223374 446464 223438
rect 446528 223374 446529 223438
rect 446463 223373 446529 223374
rect 450495 223522 450496 223586
rect 450560 223522 450561 223586
rect 450495 223521 450561 223522
rect 446079 223290 446145 223291
rect 446079 223226 446080 223290
rect 446144 223226 446145 223290
rect 446079 223225 446145 223226
rect 447810 222995 447870 223325
rect 447807 222994 447873 222995
rect 447807 222930 447808 222994
rect 447872 222930 447873 222994
rect 447807 222929 447873 222930
rect 440895 222698 440961 222699
rect 349311 222633 349377 222634
rect 440895 222634 440896 222698
rect 440960 222634 440961 222698
rect 440895 222633 440961 222634
rect 471039 53238 471105 53239
rect 471039 53174 471040 53238
rect 471104 53174 471105 53238
rect 471039 53173 471105 53174
rect 208191 52350 208257 52351
rect 208191 52286 208192 52350
rect 208256 52286 208257 52350
rect 208191 52285 208257 52286
rect 204351 51906 204417 51907
rect 204351 51842 204352 51906
rect 204416 51842 204417 51906
rect 204351 51841 204417 51842
rect 145983 51166 146049 51167
rect 145983 51102 145984 51166
rect 146048 51102 146049 51166
rect 145983 51101 146049 51102
rect 145791 51018 145857 51019
rect 145791 50954 145792 51018
rect 145856 50954 145857 51018
rect 145791 50953 145857 50954
rect 145407 50870 145473 50871
rect 145407 50806 145408 50870
rect 145472 50806 145473 50870
rect 145407 50805 145473 50806
rect 302463 45542 302529 45543
rect 302463 45478 302464 45542
rect 302528 45478 302529 45542
rect 302463 45477 302529 45478
rect 302466 43323 302526 45477
rect 305343 45394 305409 45395
rect 305343 45330 305344 45394
rect 305408 45330 305409 45394
rect 305343 45329 305409 45330
rect 305346 43323 305406 45329
rect 356991 45246 357057 45247
rect 356991 45182 356992 45246
rect 357056 45182 357057 45246
rect 356991 45181 357057 45182
rect 302463 43322 302529 43323
rect 302463 43258 302464 43322
rect 302528 43258 302529 43322
rect 302463 43257 302529 43258
rect 305343 43322 305409 43323
rect 305343 43258 305344 43322
rect 305408 43258 305409 43322
rect 305343 43257 305409 43258
rect 356994 43175 357054 45181
rect 360063 45098 360129 45099
rect 360063 45034 360064 45098
rect 360128 45034 360129 45098
rect 360063 45033 360129 45034
rect 360066 43323 360126 45033
rect 362943 44950 363009 44951
rect 362943 44886 362944 44950
rect 363008 44886 363009 44950
rect 362943 44885 363009 44886
rect 362946 43323 363006 44885
rect 360063 43322 360129 43323
rect 360063 43258 360064 43322
rect 360128 43258 360129 43322
rect 360063 43257 360129 43258
rect 362943 43322 363009 43323
rect 362943 43258 362944 43322
rect 363008 43258 363009 43322
rect 362943 43257 363009 43258
rect 356991 43174 357057 43175
rect 356991 43110 356992 43174
rect 357056 43110 357057 43174
rect 356991 43109 357057 43110
rect 471042 42139 471102 53173
rect 632130 48947 632190 223817
rect 632322 50427 632382 223817
rect 632514 51759 632574 223965
rect 632706 52203 632766 223965
rect 632895 223882 632961 223883
rect 632895 223818 632896 223882
rect 632960 223818 632961 223882
rect 632895 223817 632961 223818
rect 633279 223882 633345 223883
rect 633279 223818 633280 223882
rect 633344 223818 633345 223882
rect 633279 223817 633345 223818
rect 632703 52202 632769 52203
rect 632703 52138 632704 52202
rect 632768 52138 632769 52202
rect 632703 52137 632769 52138
rect 632898 52055 632958 223817
rect 632895 52054 632961 52055
rect 632895 51990 632896 52054
rect 632960 51990 632961 52054
rect 632895 51989 632961 51990
rect 633282 51907 633342 223817
rect 633279 51906 633345 51907
rect 633279 51842 633280 51906
rect 633344 51842 633345 51906
rect 633279 51841 633345 51842
rect 632511 51758 632577 51759
rect 632511 51694 632512 51758
rect 632576 51694 632577 51758
rect 632511 51693 632577 51694
rect 632319 50426 632385 50427
rect 632319 50362 632320 50426
rect 632384 50362 632385 50426
rect 632319 50361 632385 50362
rect 632127 48946 632193 48947
rect 632127 48882 632128 48946
rect 632192 48882 632193 48946
rect 632127 48881 632193 48882
rect 633474 48799 633534 224113
rect 673986 179779 674046 224705
rect 674178 182073 674238 226185
rect 674559 222550 674625 222551
rect 674559 222486 674560 222550
rect 674624 222486 674625 222550
rect 674559 222485 674625 222486
rect 674367 220034 674433 220035
rect 674367 219970 674368 220034
rect 674432 219970 674433 220034
rect 674367 219969 674433 219970
rect 674370 191619 674430 219969
rect 674562 193543 674622 222485
rect 674754 220809 674814 238913
rect 674946 236793 675006 244981
rect 675522 244751 675582 257265
rect 675519 244750 675585 244751
rect 675519 244686 675520 244750
rect 675584 244686 675585 244750
rect 675519 244685 675585 244686
rect 675714 238683 675774 268069
rect 675711 238682 675777 238683
rect 675711 238618 675712 238682
rect 675776 238618 675777 238682
rect 675711 238617 675777 238618
rect 674946 236733 675390 236793
rect 675330 221071 675390 236733
rect 675906 227287 675966 270881
rect 676671 256294 676737 256295
rect 676671 256230 676672 256294
rect 676736 256230 676737 256294
rect 676671 256229 676737 256230
rect 675903 227286 675969 227287
rect 675903 227222 675904 227286
rect 675968 227222 675969 227286
rect 675903 227221 675969 227222
rect 676674 225807 676734 256229
rect 676671 225806 676737 225807
rect 676671 225742 676672 225806
rect 676736 225742 676737 225806
rect 676671 225741 676737 225742
rect 675327 221070 675393 221071
rect 675327 221006 675328 221070
rect 675392 221006 675393 221070
rect 675327 221005 675393 221006
rect 674754 220749 675390 220809
rect 675135 220182 675201 220183
rect 675135 220118 675136 220182
rect 675200 220118 675201 220182
rect 675135 220117 675201 220118
rect 674943 216334 675009 216335
rect 674943 216270 674944 216334
rect 675008 216270 675009 216334
rect 674943 216269 675009 216270
rect 674751 210118 674817 210119
rect 674751 210054 674752 210118
rect 674816 210054 674817 210118
rect 674751 210053 674817 210054
rect 674559 193542 674625 193543
rect 674559 193478 674560 193542
rect 674624 193478 674625 193542
rect 674559 193477 674625 193478
rect 674367 191618 674433 191619
rect 674367 191554 674368 191618
rect 674432 191554 674433 191618
rect 674367 191553 674433 191554
rect 674175 182072 674241 182073
rect 674175 182008 674176 182072
rect 674240 182008 674241 182072
rect 674175 182007 674241 182008
rect 674175 181258 674241 181259
rect 674175 181194 674176 181258
rect 674240 181194 674241 181258
rect 674175 181193 674241 181194
rect 673983 179778 674049 179779
rect 673983 179714 673984 179778
rect 674048 179714 674049 179778
rect 673983 179713 674049 179714
rect 673986 135083 674046 179713
rect 674178 136859 674238 181193
rect 674754 180963 674814 210053
rect 674946 195319 675006 216269
rect 675138 198427 675198 220117
rect 675330 199463 675390 220749
rect 676095 206270 676161 206271
rect 676095 206206 676096 206270
rect 676160 206206 676161 206270
rect 676095 206205 676161 206206
rect 676098 204495 676158 206205
rect 676095 204494 676161 204495
rect 676095 204430 676096 204494
rect 676160 204430 676161 204494
rect 676095 204429 676161 204430
rect 675519 201682 675585 201683
rect 675519 201618 675520 201682
rect 675584 201618 675585 201682
rect 675519 201617 675585 201618
rect 675522 200055 675582 201617
rect 675519 200054 675585 200055
rect 675519 199990 675520 200054
rect 675584 199990 675585 200054
rect 675519 199989 675585 199990
rect 675327 199462 675393 199463
rect 675327 199398 675328 199462
rect 675392 199398 675393 199462
rect 675327 199397 675393 199398
rect 675135 198426 675201 198427
rect 675135 198362 675136 198426
rect 675200 198362 675201 198426
rect 675135 198361 675201 198362
rect 674943 195318 675009 195319
rect 674943 195254 674944 195318
rect 675008 195254 675009 195318
rect 674943 195253 675009 195254
rect 675519 193246 675585 193247
rect 675519 193182 675520 193246
rect 675584 193182 675585 193246
rect 675519 193181 675585 193182
rect 675327 193098 675393 193099
rect 675327 193034 675328 193098
rect 675392 193034 675393 193098
rect 675327 193033 675393 193034
rect 674751 180962 674817 180963
rect 674751 180898 674752 180962
rect 674816 180898 674817 180962
rect 674751 180897 674817 180898
rect 674367 180518 674433 180519
rect 674367 180454 674368 180518
rect 674432 180454 674433 180518
rect 674367 180453 674433 180454
rect 674370 142779 674430 180453
rect 674751 177558 674817 177559
rect 674751 177494 674752 177558
rect 674816 177494 674817 177558
rect 674751 177493 674817 177494
rect 674559 174450 674625 174451
rect 674559 174386 674560 174450
rect 674624 174386 674625 174450
rect 674559 174385 674625 174386
rect 674562 146479 674622 174385
rect 674754 148551 674814 177493
rect 674943 171342 675009 171343
rect 674943 171278 674944 171342
rect 675008 171278 675009 171342
rect 674943 171277 675009 171278
rect 674946 150327 675006 171277
rect 675330 155211 675390 193033
rect 675327 155210 675393 155211
rect 675327 155146 675328 155210
rect 675392 155146 675393 155210
rect 675327 155145 675393 155146
rect 675330 154875 675390 155145
rect 675522 155063 675582 193181
rect 675711 161426 675777 161427
rect 675711 161362 675712 161426
rect 675776 161362 675777 161426
rect 675711 161361 675777 161362
rect 675519 155062 675585 155063
rect 675519 154998 675520 155062
rect 675584 154998 675585 155062
rect 675519 154997 675585 154998
rect 675138 154815 675390 154875
rect 674943 150326 675009 150327
rect 674943 150262 674944 150326
rect 675008 150262 675009 150326
rect 674943 150261 675009 150262
rect 674751 148550 674817 148551
rect 674751 148486 674752 148550
rect 674816 148486 674817 148550
rect 674751 148485 674817 148486
rect 674559 146478 674625 146479
rect 674559 146414 674560 146478
rect 674624 146414 674625 146478
rect 674559 146413 674625 146414
rect 674367 142778 674433 142779
rect 674367 142714 674368 142778
rect 674432 142714 674433 142778
rect 674367 142713 674433 142714
rect 674175 136858 674241 136859
rect 674175 136794 674176 136858
rect 674240 136794 674241 136858
rect 674175 136793 674241 136794
rect 673983 135082 674049 135083
rect 673983 135018 673984 135082
rect 674048 135018 674049 135082
rect 673983 135017 674049 135018
rect 674559 132566 674625 132567
rect 674559 132502 674560 132566
rect 674624 132502 674625 132566
rect 674559 132501 674625 132502
rect 674367 130642 674433 130643
rect 674367 130578 674368 130642
rect 674432 130578 674433 130642
rect 674367 130577 674433 130578
rect 674175 129754 674241 129755
rect 674175 129690 674176 129754
rect 674240 129690 674241 129754
rect 674175 129689 674241 129690
rect 674178 101487 674238 129689
rect 674370 108147 674430 130577
rect 674367 108146 674433 108147
rect 674367 108082 674368 108146
rect 674432 108082 674433 108146
rect 674367 108081 674433 108082
rect 674562 103263 674622 132501
rect 675138 126795 675198 154815
rect 675135 126794 675201 126795
rect 675135 126730 675136 126794
rect 675200 126730 675201 126794
rect 675135 126729 675201 126730
rect 675138 110811 675198 126729
rect 675135 110810 675201 110811
rect 675135 110746 675136 110810
rect 675200 110746 675201 110810
rect 675135 110745 675201 110746
rect 675522 110071 675582 154997
rect 675714 153435 675774 161361
rect 675711 153434 675777 153435
rect 675711 153370 675712 153434
rect 675776 153370 675777 153434
rect 675711 153369 675777 153370
rect 675519 110070 675585 110071
rect 675519 110006 675520 110070
rect 675584 110006 675585 110070
rect 675519 110005 675585 110006
rect 674559 103262 674625 103263
rect 674559 103198 674560 103262
rect 674624 103198 674625 103262
rect 674559 103197 674625 103198
rect 674175 101486 674241 101487
rect 674175 101422 674176 101486
rect 674240 101422 674241 101486
rect 674175 101421 674241 101422
rect 633471 48798 633537 48799
rect 633471 48734 633472 48798
rect 633536 48734 633537 48798
rect 633471 48733 633537 48734
rect 471039 42138 471105 42139
rect 471039 42074 471040 42138
rect 471104 42074 471105 42138
rect 471039 42073 471105 42074
rect 189951 41842 190017 41843
rect 189951 41778 189952 41842
rect 190016 41778 190017 41842
rect 189951 41777 190017 41778
rect 194943 41842 195009 41843
rect 194943 41778 194944 41842
rect 195008 41778 195009 41842
rect 194943 41777 195009 41778
rect 518463 41842 518529 41843
rect 518463 41778 518464 41842
rect 518528 41778 518529 41842
rect 518463 41777 518529 41778
rect 189954 40807 190014 41777
rect 189951 40806 190017 40807
rect 189951 40742 189952 40806
rect 190016 40742 190017 40806
rect 189951 40741 190017 40742
rect 194946 40659 195006 41777
rect 518271 40806 518337 40807
rect 518271 40742 518272 40806
rect 518336 40742 518337 40806
rect 518271 40741 518337 40742
rect 194943 40658 195009 40659
rect 194943 40594 194944 40658
rect 195008 40594 195009 40658
rect 194943 40593 195009 40594
rect 518274 40323 518334 40741
rect 518466 40323 518526 41777
rect 518274 40263 518526 40323
<< via4 >>
rect 399146 236645 399382 236881
rect 411242 236842 411328 236881
rect 411328 236842 411392 236881
rect 411392 236842 411478 236881
rect 411242 236645 411478 236842
rect 427562 223438 427798 223561
rect 427562 223374 427648 223438
rect 427648 223374 427712 223438
rect 427712 223374 427798 223438
rect 427562 223325 427798 223374
rect 380330 222659 380566 222895
rect 400106 222659 400342 222895
rect 447722 223325 447958 223561
<< metal5 >>
rect 399104 236881 411520 236923
rect 399104 236645 399146 236881
rect 399382 236645 411242 236881
rect 411478 236645 411520 236881
rect 399104 236603 411520 236645
rect 427520 223561 448000 223603
rect 427520 223325 427562 223561
rect 427798 223325 447722 223561
rect 447958 223325 448000 223561
rect 427520 223283 448000 223325
rect 380288 222895 400384 222937
rect 380288 222659 380330 222895
rect 380566 222659 400106 222895
rect 400342 222659 400384 222895
rect 380288 222617 400384 222659
use user_id_programming  user_id_value ../mag
timestamp 1608006408
transform 1 0 656625 0 1 80926
box 0 0 7109 7077
use storage  storage ../mag
timestamp 1608006408
transform 1 0 52031 0 1 61392
box 0 0 88934 189234
use mgmt_core  soc ../mag
timestamp 1608006408
transform 1 0 204550 0 1 53700
box 0 0 430000 170000
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level ../mag
timestamp 1608006408
transform 1 0 154753 0 1 51403
box 0 1 5124 5084
use simple_por  por ../mag
timestamp 1608006408
transform 1 0 654176 0 1 104197
box 25 11 11344 8338
use mgmt_protect  mgmt_buffers ../mag
timestamp 1608006408
transform 1 0 288100 0 1 239747
box 0 0 169594 13025
use gpio_control_block  gpio_control_bidir\[1\] ../mag
timestamp 1608006408
transform -1 0 708537 0 1 166200
box 0 0 33934 18344
use gpio_control_block  gpio_control_bidir\[0\]
timestamp 1608006408
transform -1 0 708537 0 1 121000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[37\]
timestamp 1608006408
transform 1 0 8567 0 1 202600
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[36\]
timestamp 1608006408
transform 1 0 8567 0 1 245800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[3\]
timestamp 1608006408
transform -1 0 708537 0 1 256400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[2\]
timestamp 1608006408
transform -1 0 708537 0 1 211200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[35\]
timestamp 1608006408
transform 1 0 8567 0 1 289000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[34\]
timestamp 1608006408
transform 1 0 8567 0 1 332200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[33\]
timestamp 1608006408
transform 1 0 8567 0 1 375400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[5\]
timestamp 1608006408
transform -1 0 708537 0 1 346400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[4\]
timestamp 1608006408
transform -1 0 708537 0 1 301400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[7\]
timestamp 1608006408
transform -1 0 708537 0 1 479800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[6\]
timestamp 1608006408
transform -1 0 708537 0 1 391600
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[32\]
timestamp 1608006408
transform 1 0 8567 0 1 418600
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[31\]
timestamp 1608006408
transform 1 0 8567 0 1 546200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[30\]
timestamp 1608006408
transform 1 0 8567 0 1 589400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[29\]
timestamp 1608006408
transform 1 0 8567 0 1 632600
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[9\]
timestamp 1608006408
transform -1 0 708537 0 1 568800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[8\]
timestamp 1608006408
transform -1 0 708537 0 1 523800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[10\]
timestamp 1608006408
transform -1 0 708537 0 1 614000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[28\]
timestamp 1608006408
transform 1 0 8567 0 1 675800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[27\]
timestamp 1608006408
transform 1 0 8567 0 1 719000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[26\]
timestamp 1608006408
transform 1 0 8567 0 1 762200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[13\]
timestamp 1608006408
transform -1 0 708537 0 1 749200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[12\]
timestamp 1608006408
transform -1 0 708537 0 1 704200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[11\]
timestamp 1608006408
transform -1 0 708537 0 1 659000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[25\]
timestamp 1608006408
transform 1 0 8567 0 1 805400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[24\]
timestamp 1608006408
transform 1 0 8567 0 1 889800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[23\]
timestamp 1608006408
transform 0 1 97200 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[22\]
timestamp 1608006408
transform 0 1 148600 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[21\]
timestamp 1608006408
transform 0 1 200000 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[20\]
timestamp 1608006408
transform 0 1 251400 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[19\]
timestamp 1608006408
transform 0 1 303000 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[18\]
timestamp 1608006408
transform 0 1 353400 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[17\]
timestamp 1608006408
transform 0 1 420800 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[16\]
timestamp 1608006408
transform 0 1 497800 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[15\]
timestamp 1608006408
transform 0 1 549200 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[14\]
timestamp 1608006408
transform -1 0 708537 0 1 927600
box 0 0 33934 18344
use chip_io  padframe ../mag
timestamp 1608006408
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use user_project_wrapper  mprj ../mag
timestamp 1608006408
transform 1 0 65277 0 1 276402
box -8576 -7506 592500 711442
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
