* NGSPICE file created from neuron-test.ext - technology: sky130A

* Include SkyWater sky130 device models
.include "/foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice" 
.include "/foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice" 
.include "/foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice"

.param mc_mm_switch=0 
.param mc_pr_switch=1  

* DC source for current measure
Vdd vpwr gnd DC 0.7V
Vgnd vgnd gnd DC 0.0V
Vth vth gnd DC 0.1V
Vk vk gnd DC 0.15V
Vw vw gnd DC 0.01V
Vr vr gnd DC 0.37V
Vau vau gnd DC 0.08V
Vad vad gnd DC 0.25V

Idc vpwr v DC 10p

.subckt sky130_fd_pr__nfet_01v8_dlksd1 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_s3efqo VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lca7f7 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_u061qr VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_h2n75u VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_zt2j7p VSUBS a_n98_n120# a_n40_n146# a_40_n120# w_n134_n182#
X0 a_40_n120# a_n40_n146# a_n98_n120# w_n134_n182# sky130_fd_pr__pfet_01v8 w=1.2e+06u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ckptud VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_2vaynq VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_wpylm8 VSUBS a_n388_n400# a_n330_n426# a_330_n400#
X0 a_330_n400# a_n330_n426# a_n388_n400# VSUBS sky130_fd_pr__nfet_01v8 w=4e+06u l=3.3e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_9i6r5e VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_9hqhhq VSUBS a_n498_n500# a_n440_n526# a_440_n500#
X0 a_440_n500# a_n440_n526# a_n498_n500# VSUBS sky130_fd_pr__nfet_01v8 w=5e+06u l=4.4e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_h43ndc VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_6z4qh8 VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_tb02ql VSUBS a_n618_n800# a_n560_n826# a_560_n800#
X0 a_560_n800# a_n560_n826# a_n618_n800# VSUBS sky130_fd_pr__nfet_01v8 w=8e+06u l=5.6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_zgaw3c VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends


* Top level circuit neuron-test

XM10 vgnd vgnd vad a# sky130_fd_pr__nfet_01v8_dlksd1
XM11 vgnd v a# vgnd sky130_fd_pr__nfet_01v8_s3efqo
XM1 vgnd a_35_1497# v vth sky130_fd_pr__nfet_01v8_lca7f7
XM2 vgnd a_35_1497# vpwr vpwr a_35_1497# sky130_fd_pr__pfet_01v8_u061qr
XM3 vgnd a_35_1497# vpwr vpwr v sky130_fd_pr__pfet_01v8_h2n75u
XM4 vgnd vpwr a_35_1497# axon vpwr sky130_fd_pr__pfet_01v8_zt2j7p
XM5 vgnd vgnd a_35_1497# axon sky130_fd_pr__nfet_01v8_ckptud
XM6 vgnd vw axon vpwr u# sky130_fd_pr__pfet_01v8_2vaynq
XCu vgnd vgnd u# vgnd sky130_fd_pr__nfet_01v8_wpylm8
XM7 vgnd vgnd vr u# sky130_fd_pr__nfet_01v8_9i6r5e
XCv vgnd vgnd v vgnd sky130_fd_pr__nfet_01v8_9hqhhq
XM8 vgnd v u# vgnd sky130_fd_pr__nfet_01v8_h43ndc
XM9 vgnd vau axon vpwr a# sky130_fd_pr__pfet_01v8_6z4qh8
XCa vgnd vgnd a# vgnd sky130_fd_pr__nfet_01v8_tb02ql
XMk vgnd v vk vgnd sky130_fd_pr__nfet_01v8_zgaw3c

.IC V(v)=0 V(u#)=0 V(a#)=0

.control
* Sweep tran
tran 1u 20m uic
plot v(v)
.endc
.end

