magic
tech sky130A
magscale 1 2
timestamp 1605923309
<< nwell >>
rect -109 -180 109 180
<< pmos >>
rect -15 -80 15 80
<< pdiff >>
rect -73 68 -15 80
rect -73 -68 -61 68
rect -27 -68 -15 68
rect -73 -80 -15 -68
rect 15 68 73 80
rect 15 -68 27 68
rect 61 -68 73 68
rect 15 -80 73 -68
<< pdiffc >>
rect -61 -68 -27 68
rect 27 -68 61 68
<< poly >>
rect -33 161 33 177
rect -33 127 -17 161
rect 17 127 33 161
rect -33 111 33 127
rect -15 80 15 111
rect -15 -111 15 -80
rect -33 -127 33 -111
rect -33 -161 -17 -127
rect 17 -161 33 -127
rect -33 -177 33 -161
<< polycont >>
rect -17 127 17 161
rect -17 -161 17 -127
<< locali >>
rect -33 127 -17 161
rect 17 127 33 161
rect -61 68 -27 84
rect -61 -84 -27 -68
rect 27 68 61 84
rect 27 -84 61 -68
rect -33 -161 -17 -127
rect 17 -161 33 -127
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.8 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0
string library sky130
<< end >>
