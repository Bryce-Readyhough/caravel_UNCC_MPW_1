magic
tech sky130A
magscale 1 2
timestamp 1606526574
<< error_s >>
rect 444 356 456 362
rect 406 350 462 356
rect 400 344 468 350
rect 400 338 418 344
rect 412 312 418 338
rect 450 338 468 344
rect 450 312 462 338
rect 412 306 462 312
rect 444 300 462 306
rect 444 294 456 300
rect 3162 -72 3174 -66
rect 3124 -78 3180 -72
rect 3118 -84 3186 -78
rect 3118 -90 3136 -84
rect 3130 -116 3136 -90
rect 3168 -90 3186 -84
rect 3168 -116 3180 -90
rect 3130 -122 3180 -116
rect 3162 -128 3180 -122
rect 3162 -134 3174 -128
rect 428 -922 440 -916
rect 390 -928 446 -922
rect 384 -934 452 -928
rect 384 -940 402 -934
rect 396 -966 402 -940
rect 434 -940 452 -934
rect 434 -966 446 -940
rect 396 -972 446 -966
rect 428 -978 446 -972
rect 428 -984 440 -978
<< pwell >>
rect 3078 -162 3232 -24
<< metal1 >>
rect 1872 669 2901 711
rect 2859 457 2901 669
rect 2803 -568 2845 -377
rect 1856 -610 2845 -568
use Sw-1  Sw-1_2
timestamp 1606521356
transform 1 0 2850 0 1 -512
box -140 90 1782 1018
use Sw-1  Sw-1_1
timestamp 1606521356
transform 1 0 116 0 1 -1362
box -140 90 1782 1018
use Sw-1  Sw-1_0
timestamp 1606521356
transform 1 0 132 0 1 -84
box -140 90 1782 1018
<< end >>
