.subckt untitled-5
XR1 B A __UNCONNECTED_PIN__ sky130_fd_pr__res_generic_po W=1 L=1 mult=1 m=1
**** begin user architecture code

blabla


blabla

**** end user architecture code
.ends
.end
