magic
tech sky130A
magscale 1 2
timestamp 1604444418
<< nwell >>
rect -92 1604 477 1893
rect -43 1560 477 1604
rect 120 1403 205 1560
rect 930 1260 2051 1890
<< psubdiff >>
rect -57 -330 813 -303
rect -57 -390 -30 -330
rect 30 -390 120 -330
rect 180 -390 270 -330
rect 330 -390 420 -330
rect 480 -390 568 -330
rect 628 -331 813 -330
rect 628 -390 718 -331
rect -57 -391 718 -390
rect 778 -391 813 -331
rect -57 -416 813 -391
rect 930 -330 1470 -300
rect 930 -390 960 -330
rect 1020 -390 1110 -330
rect 1170 -390 1260 -330
rect 1320 -390 1380 -330
rect 1440 -390 1470 -330
rect 930 -420 1470 -390
rect 2460 -330 2580 -300
rect 2460 -390 2490 -330
rect 2550 -390 2580 -330
rect 2460 -420 2580 -390
<< nsubdiff >>
rect 1114 1830 1824 1854
rect -23 1801 385 1826
rect -23 1800 302 1801
rect -23 1740 0 1800
rect 60 1740 149 1800
rect 209 1741 302 1800
rect 362 1741 385 1801
rect 1114 1770 1140 1830
rect 1200 1770 1290 1830
rect 1350 1770 1440 1830
rect 1500 1770 1590 1830
rect 1650 1770 1740 1830
rect 1800 1770 1824 1830
rect 1114 1744 1824 1770
rect 209 1740 385 1741
rect -23 1713 385 1740
<< psubdiffcont >>
rect -30 -390 30 -330
rect 120 -390 180 -330
rect 270 -390 330 -330
rect 420 -390 480 -330
rect 568 -390 628 -330
rect 718 -391 778 -331
rect 960 -390 1020 -330
rect 1110 -390 1170 -330
rect 1260 -390 1320 -330
rect 1380 -390 1440 -330
rect 2490 -390 2550 -330
<< nsubdiffcont >>
rect 0 1740 60 1800
rect 149 1740 209 1800
rect 302 1741 362 1801
rect 1140 1770 1200 1830
rect 1290 1770 1350 1830
rect 1440 1770 1500 1830
rect 1590 1770 1650 1830
rect 1740 1770 1800 1830
<< poly >>
rect 2308 1830 3428 1866
rect 2308 1770 2370 1830
rect 2430 1770 2520 1830
rect 2580 1770 2670 1830
rect 2730 1770 2820 1830
rect 2880 1770 2970 1830
rect 3030 1770 3120 1830
rect 3180 1770 3270 1830
rect 3330 1770 3428 1830
rect 2308 1730 3428 1770
rect 35 1553 242 1577
rect 35 1516 149 1553
rect 184 1516 242 1553
rect 1414 1528 1494 1577
rect 1823 1527 1903 1576
rect 35 1497 242 1516
rect 551 1478 680 1488
rect 551 1418 567 1478
rect 627 1418 680 1478
rect 551 1408 680 1418
rect -62 1290 818 1320
rect -62 1230 -30 1290
rect 30 1230 120 1290
rect 180 1230 270 1290
rect 330 1230 420 1290
rect 480 1230 570 1290
rect 630 1230 720 1290
rect 780 1230 818 1290
rect -62 1202 818 1230
rect 1025 1262 1105 1324
rect 1025 1196 1044 1262
rect 1086 1196 1105 1262
rect 1025 1186 1105 1196
rect 1287 1170 1947 1200
rect 1287 1110 1350 1170
rect 1410 1110 1500 1170
rect 1560 1110 1650 1170
rect 1710 1110 1800 1170
rect 1860 1110 1947 1170
rect 1287 1073 1947 1110
rect 1287 210 1947 247
rect -62 120 818 166
rect 1287 150 1350 210
rect 1410 150 1500 210
rect 1560 150 1650 210
rect 1710 150 1800 210
rect 1860 150 1947 210
rect -62 60 -30 120
rect 30 60 120 120
rect 180 60 270 120
rect 330 60 420 120
rect 480 60 570 120
rect 630 60 720 120
rect 780 60 818 120
rect -62 26 818 60
rect 1026 97 1106 121
rect 1287 120 1947 150
rect 1026 31 1045 97
rect 1087 31 1106 97
rect 1026 -9 1106 31
rect 2308 60 3428 108
rect 1669 13 1735 23
rect 1669 -21 1685 13
rect 1719 -21 1735 13
rect 1669 -31 1735 -21
rect 2308 0 2370 60
rect 2430 0 2520 60
rect 2580 0 2670 60
rect 2730 0 2820 60
rect 2880 0 2970 60
rect 3030 0 3120 60
rect 3180 0 3270 60
rect 3330 0 3428 60
rect 2308 -30 3428 0
rect -80 -188 -42 -108
rect 270 -121 352 -108
rect 241 -131 352 -121
rect 569 -122 655 -108
rect 2984 -115 3050 -105
rect 241 -165 257 -131
rect 291 -165 352 -131
rect 241 -175 352 -165
rect 270 -188 352 -175
rect 543 -132 655 -122
rect 543 -166 559 -132
rect 593 -166 655 -132
rect 1374 -156 1454 -118
rect 2984 -149 3000 -115
rect 3034 -149 3050 -115
rect 2984 -159 3050 -149
rect 543 -176 655 -166
rect 569 -188 655 -176
rect 2546 -256 2626 -207
<< polycont >>
rect 2370 1770 2430 1830
rect 2520 1770 2580 1830
rect 2670 1770 2730 1830
rect 2820 1770 2880 1830
rect 2970 1770 3030 1830
rect 3120 1770 3180 1830
rect 3270 1770 3330 1830
rect 149 1516 184 1553
rect 567 1418 627 1478
rect -30 1230 30 1290
rect 120 1230 180 1290
rect 270 1230 330 1290
rect 420 1230 480 1290
rect 570 1230 630 1290
rect 720 1230 780 1290
rect 1044 1196 1086 1262
rect 1350 1110 1410 1170
rect 1500 1110 1560 1170
rect 1650 1110 1710 1170
rect 1800 1110 1860 1170
rect 1350 150 1410 210
rect 1500 150 1560 210
rect 1650 150 1710 210
rect 1800 150 1860 210
rect -30 60 30 120
rect 120 60 180 120
rect 270 60 330 120
rect 420 60 480 120
rect 570 60 630 120
rect 720 60 780 120
rect 1045 31 1087 97
rect 1685 -21 1719 13
rect 2370 0 2430 60
rect 2520 0 2580 60
rect 2670 0 2730 60
rect 2820 0 2880 60
rect 2970 0 3030 60
rect 3120 0 3180 60
rect 3270 0 3330 60
rect 257 -165 291 -131
rect 559 -166 593 -132
rect 3000 -149 3034 -115
<< locali >>
rect 0 2130 360 2160
rect 60 2070 150 2130
rect 210 2070 300 2130
rect 0 1817 360 2070
rect 1110 2130 1830 2160
rect 1110 2070 1140 2130
rect 1200 2070 1290 2130
rect 1350 2070 1440 2130
rect 1500 2070 1590 2130
rect 1650 2070 1740 2130
rect 1800 2070 1830 2130
rect 1110 1920 1830 2070
rect 978 1883 1830 1920
rect -16 1801 377 1817
rect -16 1800 302 1801
rect -16 1740 0 1800
rect 60 1740 149 1800
rect 209 1741 302 1800
rect 362 1741 377 1801
rect 209 1740 377 1741
rect -16 1737 377 1740
rect -34 1733 377 1737
rect -34 1721 420 1733
rect -34 1608 135 1721
rect 251 1604 420 1721
rect 681 1724 777 1728
rect 681 1674 694 1724
rect 746 1674 777 1724
rect 681 1574 777 1674
rect 132 1553 202 1572
rect 132 1516 149 1553
rect 184 1516 202 1553
rect 132 1485 202 1516
rect 458 1540 777 1574
rect 978 1573 1015 1883
rect 1110 1830 1830 1883
rect 1122 1770 1140 1830
rect 1200 1770 1290 1830
rect 1350 1770 1440 1830
rect 1500 1770 1590 1830
rect 1650 1770 1740 1830
rect 1800 1770 1818 1830
rect 2340 1829 2370 1830
rect 1122 1753 1818 1770
rect 1915 1795 2370 1829
rect 979 1549 1013 1573
rect 1247 1569 1811 1603
rect 458 1485 492 1540
rect 681 1517 777 1540
rect 682 1500 775 1517
rect 1247 1516 1281 1569
rect 567 1488 627 1494
rect -93 1290 75 1464
rect 132 1451 256 1485
rect 390 1451 492 1485
rect 557 1478 637 1488
rect 132 1446 202 1451
rect 557 1418 567 1478
rect 627 1418 637 1478
rect 557 1290 637 1418
rect 1117 1453 1402 1516
rect 1777 1480 1811 1569
rect 1915 1471 1949 1795
rect 2340 1770 2370 1795
rect 2430 1770 2520 1830
rect 2580 1770 2670 1830
rect 2730 1770 2820 1830
rect 2880 1770 2970 1830
rect 3030 1770 3120 1830
rect 3180 1770 3270 1830
rect 3330 1770 3360 1830
rect 2220 1631 2281 1710
rect 3468 1679 3540 1710
rect 3468 1638 3469 1679
rect 3517 1638 3540 1679
rect 2220 1590 2234 1631
rect 2220 1511 2281 1590
rect 3468 1555 3540 1638
rect 3468 1514 3469 1555
rect 3517 1514 3540 1555
rect 1117 1401 1222 1453
rect 1276 1401 1402 1453
rect 767 1362 839 1396
rect 1117 1350 1402 1401
rect 2220 1470 2234 1511
rect 2220 1391 2281 1470
rect 3468 1431 3540 1514
rect -60 1230 -30 1290
rect 30 1230 120 1290
rect 180 1230 270 1290
rect 330 1230 420 1290
rect 480 1230 570 1290
rect 630 1230 720 1290
rect 780 1230 810 1290
rect 1037 1262 1096 1284
rect -150 1129 -90 1200
rect -150 1090 -138 1129
rect -93 1090 -90 1129
rect -150 1041 -90 1090
rect -150 1002 -138 1041
rect -93 1002 -90 1041
rect -150 953 -90 1002
rect -150 914 -138 953
rect -93 914 -90 953
rect -150 865 -90 914
rect -150 826 -138 865
rect -93 826 -90 865
rect -150 777 -90 826
rect -150 738 -138 777
rect -93 738 -90 777
rect -150 689 -90 738
rect -150 650 -138 689
rect -93 650 -90 689
rect -150 601 -90 650
rect -150 562 -138 601
rect -93 562 -90 601
rect -150 513 -90 562
rect -150 474 -138 513
rect -93 474 -90 513
rect -150 425 -90 474
rect -150 386 -138 425
rect -93 386 -90 425
rect -150 337 -90 386
rect -150 298 -138 337
rect -93 298 -90 337
rect -150 249 -90 298
rect -150 210 -138 249
rect -93 210 -90 249
rect -150 180 -90 210
rect 840 1139 900 1200
rect 840 1100 845 1139
rect 890 1100 900 1139
rect 1037 1194 1044 1262
rect 1086 1194 1096 1262
rect 1037 1137 1096 1194
rect 1506 1170 1540 1379
rect 2220 1350 2234 1391
rect 3468 1390 3469 1431
rect 3517 1390 3540 1431
rect 2220 1271 2281 1350
rect 3468 1307 3540 1390
rect 2220 1230 2234 1271
rect 3468 1266 3469 1307
rect 3517 1266 3540 1307
rect 1320 1110 1350 1170
rect 1410 1110 1500 1170
rect 1560 1110 1650 1170
rect 1710 1110 1800 1170
rect 1860 1110 1890 1170
rect 2220 1151 2281 1230
rect 3468 1183 3540 1266
rect 2220 1110 2234 1151
rect 3468 1142 3469 1183
rect 3517 1142 3540 1183
rect 840 1050 900 1100
rect 840 1011 845 1050
rect 890 1011 900 1050
rect 840 961 900 1011
rect 840 922 845 961
rect 890 922 900 961
rect 840 872 900 922
rect 840 833 845 872
rect 890 833 900 872
rect 840 783 900 833
rect 840 744 845 783
rect 890 744 900 783
rect 840 694 900 744
rect 840 655 845 694
rect 890 655 900 694
rect 840 605 900 655
rect 840 566 845 605
rect 890 566 900 605
rect 840 516 900 566
rect 840 477 845 516
rect 890 477 900 516
rect 840 427 900 477
rect 840 388 845 427
rect 890 388 900 427
rect 840 338 900 388
rect 840 299 845 338
rect 890 299 900 338
rect 840 249 900 299
rect 1200 1012 1275 1065
rect 1200 972 1214 1012
rect 1260 972 1275 1012
rect 1200 916 1275 972
rect 1200 876 1214 916
rect 1260 876 1275 916
rect 1200 820 1275 876
rect 1200 780 1214 820
rect 1260 780 1275 820
rect 1200 724 1275 780
rect 1200 684 1214 724
rect 1260 684 1275 724
rect 1200 628 1275 684
rect 1200 588 1214 628
rect 1260 588 1275 628
rect 1200 532 1275 588
rect 1200 492 1214 532
rect 1260 492 1275 532
rect 1200 436 1275 492
rect 1200 396 1214 436
rect 1260 396 1275 436
rect 1200 340 1275 396
rect 1200 300 1214 340
rect 1260 300 1275 340
rect 1200 257 1275 300
rect 1959 1013 2040 1065
rect 1959 972 1979 1013
rect 2026 972 2040 1013
rect 1959 917 2040 972
rect 1959 876 1979 917
rect 2026 876 2040 917
rect 1959 821 2040 876
rect 1959 780 1979 821
rect 2026 780 2040 821
rect 1959 725 2040 780
rect 1959 684 1979 725
rect 2026 684 2040 725
rect 1959 629 2040 684
rect 1959 588 1979 629
rect 2026 588 2040 629
rect 1959 533 2040 588
rect 1959 492 1979 533
rect 2026 492 2040 533
rect 1959 437 2040 492
rect 1959 396 1979 437
rect 2026 396 2040 437
rect 1959 341 2040 396
rect 1959 300 1979 341
rect 2026 300 2040 341
rect 1959 257 2040 300
rect 2220 1031 2281 1110
rect 3468 1059 3540 1142
rect 2220 990 2234 1031
rect 3468 1018 3469 1059
rect 3517 1018 3540 1059
rect 2220 911 2281 990
rect 3468 935 3540 1018
rect 2220 870 2234 911
rect 3468 894 3469 935
rect 3517 894 3540 935
rect 2220 791 2281 870
rect 3468 811 3540 894
rect 2220 750 2234 791
rect 3468 770 3469 811
rect 3517 770 3540 811
rect 2220 671 2281 750
rect 3468 687 3540 770
rect 2220 630 2234 671
rect 3468 646 3469 687
rect 3517 646 3540 687
rect 2220 551 2281 630
rect 3468 563 3540 646
rect 2220 510 2234 551
rect 3468 522 3469 563
rect 3517 522 3540 563
rect 2220 431 2281 510
rect 3468 439 3540 522
rect 2220 390 2234 431
rect 3468 398 3469 439
rect 3517 398 3540 439
rect 2220 311 2281 390
rect 3468 315 3540 398
rect 2220 270 2234 311
rect 3468 274 3469 315
rect 3517 274 3540 315
rect 840 210 845 249
rect 890 210 900 249
rect 840 180 900 210
rect 1320 150 1350 210
rect 1410 150 1500 210
rect 1560 150 1650 210
rect 1710 150 1800 210
rect 1860 150 1890 210
rect 2220 191 2281 270
rect 3468 191 3540 274
rect 2220 150 2234 191
rect 3468 150 3469 191
rect 3517 150 3540 191
rect -60 60 -30 120
rect 30 60 120 120
rect 180 60 270 120
rect 330 60 420 120
rect 480 60 570 120
rect 630 60 720 120
rect 780 60 810 120
rect 1037 98 1096 150
rect -33 -75 59 60
rect 355 -78 449 60
rect 657 -76 749 60
rect 1037 30 1045 98
rect 1087 30 1096 98
rect 1037 14 1096 30
rect 1210 78 1266 80
rect 1264 26 1266 78
rect 1210 -18 1266 26
rect 236 -131 313 -111
rect 236 -165 257 -131
rect 291 -165 313 -131
rect 236 -183 313 -165
rect 538 -132 615 -112
rect 538 -166 559 -132
rect 593 -166 615 -132
rect 538 -184 615 -166
rect -33 -300 59 -213
rect 356 -300 448 -214
rect 658 -300 750 -211
rect 980 -300 1015 -87
rect 1132 -109 1266 -18
rect 1466 -42 1500 150
rect 1683 31 1726 150
rect 2220 120 2281 150
rect 3468 120 3540 150
rect 1663 13 1740 31
rect 1663 -21 1685 13
rect 1719 -21 1740 13
rect 2340 0 2370 60
rect 2430 0 2520 60
rect 2580 0 2670 60
rect 2730 0 2820 60
rect 2880 0 2970 60
rect 3030 0 3120 60
rect 3180 0 3270 60
rect 3330 0 3360 60
rect 1663 -41 1740 -21
rect 1210 -110 1266 -109
rect 1327 -300 1362 -107
rect 2637 -124 2671 0
rect 3000 -97 3037 0
rect 2978 -115 3055 -97
rect 2978 -149 3000 -115
rect 3034 -149 3055 -115
rect 2978 -169 3055 -149
rect 2500 -300 2534 -197
rect -60 -330 810 -300
rect -60 -390 -30 -330
rect 30 -390 120 -330
rect 180 -390 270 -330
rect 330 -390 420 -330
rect 480 -390 568 -330
rect 628 -331 810 -330
rect 628 -390 718 -331
rect -60 -391 718 -390
rect 778 -391 810 -331
rect -60 -450 810 -391
rect -60 -510 -30 -450
rect 30 -510 120 -450
rect 180 -510 270 -450
rect 330 -510 420 -450
rect 480 -510 570 -450
rect 630 -510 720 -450
rect 780 -510 810 -450
rect -60 -540 810 -510
rect 930 -330 1470 -300
rect 930 -390 960 -330
rect 1020 -390 1110 -330
rect 1170 -390 1260 -330
rect 1320 -390 1380 -330
rect 1440 -390 1470 -330
rect 930 -450 1470 -390
rect 930 -510 960 -450
rect 1020 -510 1110 -450
rect 1170 -510 1260 -450
rect 1320 -510 1380 -450
rect 1440 -510 1470 -450
rect 930 -540 1470 -510
rect 2460 -330 2580 -300
rect 2460 -390 2490 -330
rect 2550 -390 2580 -330
rect 2460 -450 2580 -390
rect 2460 -510 2490 -450
rect 2550 -510 2580 -450
rect 2460 -540 2580 -510
<< viali >>
rect 0 2070 60 2130
rect 150 2070 210 2130
rect 300 2070 360 2130
rect 1140 2070 1200 2130
rect 1290 2070 1350 2130
rect 1440 2070 1500 2130
rect 1590 2070 1650 2130
rect 1740 2070 1800 2130
rect 694 1674 746 1724
rect 3469 1638 3517 1679
rect 2234 1590 2282 1631
rect 3469 1514 3517 1555
rect 1222 1401 1276 1453
rect 839 1362 873 1396
rect 2234 1470 2282 1511
rect -138 1090 -93 1129
rect -138 1002 -93 1041
rect -138 914 -93 953
rect -138 826 -93 865
rect -138 738 -93 777
rect -138 650 -93 689
rect -138 562 -93 601
rect -138 474 -93 513
rect -138 386 -93 425
rect -138 298 -93 337
rect -138 210 -93 249
rect 845 1100 890 1139
rect 1044 1196 1086 1261
rect 1044 1194 1086 1196
rect 2234 1350 2282 1391
rect 3469 1390 3517 1431
rect 2234 1230 2282 1271
rect 3469 1266 3517 1307
rect 2234 1110 2282 1151
rect 3469 1142 3517 1183
rect 845 1011 890 1050
rect 845 922 890 961
rect 845 833 890 872
rect 845 744 890 783
rect 845 655 890 694
rect 845 566 890 605
rect 845 477 890 516
rect 845 388 890 427
rect 845 299 890 338
rect 1214 972 1260 1012
rect 1214 876 1260 916
rect 1214 780 1260 820
rect 1214 684 1260 724
rect 1214 588 1260 628
rect 1214 492 1260 532
rect 1214 396 1260 436
rect 1214 300 1260 340
rect 1979 972 2026 1013
rect 1979 876 2026 917
rect 1979 780 2026 821
rect 1979 684 2026 725
rect 1979 588 2026 629
rect 1979 492 2026 533
rect 1979 396 2026 437
rect 1979 300 2026 341
rect 2234 990 2282 1031
rect 3469 1018 3517 1059
rect 2234 870 2282 911
rect 3469 894 3517 935
rect 2234 750 2282 791
rect 3469 770 3517 811
rect 2234 630 2282 671
rect 3469 646 3517 687
rect 2234 510 2282 551
rect 3469 522 3517 563
rect 2234 390 2282 431
rect 3469 398 3517 439
rect 2234 270 2282 311
rect 3469 274 3517 315
rect 845 210 890 249
rect 2234 150 2282 191
rect 3469 150 3517 191
rect 1045 97 1087 98
rect 1045 31 1087 97
rect 1045 30 1087 31
rect 1210 26 1264 78
rect 257 -165 291 -131
rect 559 -166 593 -132
rect 1685 -21 1719 13
rect 3000 -149 3034 -115
rect -30 -510 30 -450
rect 120 -510 180 -450
rect 270 -510 330 -450
rect 420 -510 480 -450
rect 570 -510 630 -450
rect 720 -510 780 -450
rect 960 -510 1020 -450
rect 1110 -510 1170 -450
rect 1260 -510 1320 -450
rect 1380 -510 1440 -450
rect 2490 -510 2550 -450
<< metal1 >>
rect -270 2130 3600 2190
rect -270 2070 0 2130
rect 60 2070 150 2130
rect 210 2070 300 2130
rect 360 2070 1140 2130
rect 1200 2070 1290 2130
rect 1350 2070 1440 2130
rect 1500 2070 1590 2130
rect 1650 2070 1740 2130
rect 1800 2070 3600 2130
rect -270 1950 3600 2070
rect 679 1724 1107 1743
rect 679 1674 694 1724
rect 746 1674 1107 1724
rect 679 1661 1107 1674
rect -330 1396 890 1408
rect -330 1362 839 1396
rect 873 1362 890 1396
rect -330 1350 890 1362
rect 1025 1261 1107 1661
rect 2220 1679 3540 1710
rect 2220 1638 3469 1679
rect 3517 1638 3540 1679
rect 2220 1631 3540 1638
rect 2220 1590 2234 1631
rect 2282 1590 3540 1631
rect 2220 1555 3540 1590
rect 2220 1514 3469 1555
rect 3517 1514 3540 1555
rect 2220 1511 3540 1514
rect 1200 1464 1303 1472
rect 1200 1383 1208 1464
rect 1292 1383 1303 1464
rect 1200 1369 1303 1383
rect 2220 1470 2234 1511
rect 2282 1470 3540 1511
rect 2220 1431 3540 1470
rect 2220 1391 3469 1431
rect -150 1140 -60 1200
rect 810 1140 900 1200
rect -150 1139 900 1140
rect -150 1129 845 1139
rect -150 1090 -138 1129
rect -93 1100 845 1129
rect 890 1100 900 1139
rect -93 1090 900 1100
rect -150 1050 900 1090
rect -150 1041 845 1050
rect -150 1002 -138 1041
rect -93 1011 845 1041
rect 890 1011 900 1050
rect -93 1002 900 1011
rect -150 961 900 1002
rect -150 953 845 961
rect -150 914 -138 953
rect -93 922 845 953
rect 890 922 900 961
rect -93 914 900 922
rect -150 872 900 914
rect -150 865 845 872
rect -150 826 -138 865
rect -93 833 845 865
rect 890 833 900 872
rect -93 826 900 833
rect -150 783 900 826
rect -150 777 845 783
rect -150 738 -138 777
rect -93 744 845 777
rect 890 744 900 783
rect -93 738 900 744
rect -150 694 900 738
rect -150 689 845 694
rect -150 650 -138 689
rect -93 655 845 689
rect 890 655 900 694
rect -93 650 900 655
rect -150 605 900 650
rect -150 601 845 605
rect -150 562 -138 601
rect -93 566 845 601
rect 890 566 900 605
rect -93 562 900 566
rect -150 516 900 562
rect -150 513 845 516
rect -150 474 -138 513
rect -93 477 845 513
rect 890 477 900 516
rect -93 474 900 477
rect -150 427 900 474
rect -150 425 845 427
rect -150 386 -138 425
rect -93 388 845 425
rect 890 388 900 427
rect -93 386 900 388
rect -150 338 900 386
rect -150 337 845 338
rect -150 298 -138 337
rect -93 299 845 337
rect 890 299 900 338
rect -93 298 900 299
rect -150 249 900 298
rect -150 210 -138 249
rect -93 240 845 249
rect -93 210 -60 240
rect -150 180 -60 210
rect 810 210 845 240
rect 890 210 900 249
rect 810 180 900 210
rect 236 -122 313 -111
rect 236 -174 248 -122
rect 300 -174 313 -122
rect 236 -183 313 -174
rect 538 -123 615 -112
rect 538 -175 550 -123
rect 602 -175 615 -123
rect 538 -184 615 -175
rect 840 -300 900 180
rect 1025 1194 1044 1261
rect 1086 1194 1107 1261
rect 1025 98 1107 1194
rect 2220 1350 2234 1391
rect 2282 1390 3469 1391
rect 3517 1390 3540 1431
rect 2282 1350 3540 1390
rect 2220 1307 3540 1350
rect 2220 1271 3469 1307
rect 2220 1230 2234 1271
rect 2282 1266 3469 1271
rect 3517 1266 3540 1307
rect 2282 1230 3540 1266
rect 2220 1183 3540 1230
rect 2220 1151 3469 1183
rect 2220 1110 2234 1151
rect 2282 1142 3469 1151
rect 3517 1142 3540 1183
rect 2282 1110 3540 1142
rect 2220 1059 3540 1110
rect 1200 1013 2040 1050
rect 1200 1012 1979 1013
rect 1200 972 1214 1012
rect 1260 972 1979 1012
rect 2026 972 2040 1013
rect 1200 917 2040 972
rect 1200 916 1979 917
rect 1200 876 1214 916
rect 1260 876 1979 916
rect 2026 876 2040 917
rect 1200 821 2040 876
rect 1200 820 1979 821
rect 1200 780 1214 820
rect 1260 780 1979 820
rect 2026 780 2040 821
rect 1200 725 2040 780
rect 1200 724 1979 725
rect 1200 684 1214 724
rect 1260 684 1979 724
rect 2026 684 2040 725
rect 1200 629 2040 684
rect 1200 628 1979 629
rect 1200 588 1214 628
rect 1260 588 1979 628
rect 2026 588 2040 629
rect 1200 533 2040 588
rect 1200 532 1979 533
rect 1200 492 1214 532
rect 1260 492 1979 532
rect 2026 492 2040 533
rect 1200 437 2040 492
rect 1200 436 1979 437
rect 1200 396 1214 436
rect 1260 396 1979 436
rect 2026 396 2040 437
rect 1200 341 2040 396
rect 1200 340 1979 341
rect 1200 300 1214 340
rect 1260 300 1979 340
rect 2026 300 2040 341
rect 1200 270 2040 300
rect 1025 30 1045 98
rect 1087 30 1107 98
rect 1025 14 1107 30
rect 1188 89 1291 97
rect 1188 8 1196 89
rect 1280 8 1291 89
rect 1188 -6 1291 8
rect 1663 22 1740 31
rect 1663 -30 1676 22
rect 1728 -30 1740 22
rect 1663 -41 1740 -30
rect 1980 -300 2040 270
rect 2220 1031 3469 1059
rect 2220 990 2234 1031
rect 2282 1018 3469 1031
rect 3517 1018 3540 1059
rect 2282 990 3540 1018
rect 2220 935 3540 990
rect 2220 911 3469 935
rect 2220 870 2234 911
rect 2282 894 3469 911
rect 3517 894 3540 935
rect 2282 870 3540 894
rect 2220 811 3540 870
rect 2220 791 3469 811
rect 2220 750 2234 791
rect 2282 770 3469 791
rect 3517 770 3540 811
rect 2282 750 3540 770
rect 2220 687 3540 750
rect 2220 671 3469 687
rect 2220 630 2234 671
rect 2282 646 3469 671
rect 3517 646 3540 687
rect 2282 630 3540 646
rect 2220 563 3540 630
rect 2220 551 3469 563
rect 2220 510 2234 551
rect 2282 522 3469 551
rect 3517 522 3540 563
rect 2282 510 3540 522
rect 2220 439 3540 510
rect 2220 431 3469 439
rect 2220 390 2234 431
rect 2282 398 3469 431
rect 3517 398 3540 439
rect 2282 390 3540 398
rect 2220 315 3540 390
rect 2220 311 3469 315
rect 2220 270 2234 311
rect 2282 274 3469 311
rect 3517 274 3540 315
rect 2282 270 3540 274
rect 2220 191 3540 270
rect 2220 150 2234 191
rect 2282 150 3469 191
rect 3517 150 3540 191
rect 2220 120 3540 150
rect 2978 -106 3055 -97
rect 2978 -158 2991 -106
rect 3043 -158 3055 -106
rect 2978 -169 3055 -158
rect 3450 -300 3540 120
rect -240 -450 3630 -300
rect -240 -510 -30 -450
rect 30 -510 120 -450
rect 180 -510 270 -450
rect 330 -510 420 -450
rect 480 -510 570 -450
rect 630 -510 720 -450
rect 780 -510 960 -450
rect 1020 -510 1110 -450
rect 1170 -510 1260 -450
rect 1320 -510 1380 -450
rect 1440 -510 2490 -450
rect 2550 -510 3630 -450
rect -240 -540 3630 -510
<< via1 >>
rect 1208 1453 1292 1464
rect 1208 1401 1222 1453
rect 1222 1401 1276 1453
rect 1276 1401 1292 1453
rect 1208 1383 1292 1401
rect 248 -131 300 -122
rect 248 -165 257 -131
rect 257 -165 291 -131
rect 291 -165 300 -131
rect 248 -174 300 -165
rect 550 -132 602 -123
rect 550 -166 559 -132
rect 559 -166 593 -132
rect 593 -166 602 -132
rect 550 -175 602 -166
rect 1196 78 1280 89
rect 1196 26 1210 78
rect 1210 26 1264 78
rect 1264 26 1280 78
rect 1196 8 1280 26
rect 1676 13 1728 22
rect 1676 -21 1685 13
rect 1685 -21 1719 13
rect 1719 -21 1728 13
rect 1676 -30 1728 -21
rect 2991 -115 3043 -106
rect 2991 -149 3000 -115
rect 3000 -149 3034 -115
rect 3034 -149 3043 -115
rect 2991 -158 3043 -149
<< metal2 >>
rect 1157 1464 1303 1472
rect 1157 1383 1208 1464
rect 1292 1383 1303 1464
rect 1157 1369 1303 1383
rect 1157 97 1221 1369
rect 1157 89 1291 97
rect 1157 8 1196 89
rect 1280 8 1291 89
rect 1157 -6 1291 8
rect 1663 22 1740 31
rect 1663 -30 1676 22
rect 1728 -30 1740 22
rect 1663 -41 1740 -30
rect 236 -122 313 -111
rect 236 -174 248 -122
rect 300 -174 313 -122
rect 236 -183 313 -174
rect 538 -123 615 -112
rect 538 -175 550 -123
rect 602 -175 615 -123
rect 257 -392 291 -183
rect 538 -184 615 -175
rect 559 -285 593 -184
rect 1686 -285 1720 -41
rect 2978 -106 3055 -97
rect 2978 -158 2991 -106
rect 3043 -158 3055 -106
rect 2978 -169 3055 -158
rect 559 -319 1720 -285
rect 3001 -392 3035 -169
rect 257 -426 3035 -392
use sky130_fd_pr__pfet_01v8_zt2j7p  M4
timestamp 1604306825
transform 1 0 1065 0 1 1460
box -134 -182 134 182
use sky130_fd_pr__nfet_01v8_ckptud  M5
timestamp 1604306825
transform 1 0 1066 0 1 -64
box -98 -68 98 68
use sky130_fd_pr__nfet_01v8_h43ndc  M8
timestamp 1604306825
transform 0 1 703 -1 0 -148
box -98 -68 98 68
use sky130_fd_pr__nfet_01v8_s3efqo  M11
timestamp 1604306825
transform 0 1 402 -1 0 -148
box -98 -68 98 68
use sky130_fd_pr__nfet_01v8_zgaw3c  Mk
timestamp 1604306825
transform 0 1 13 -1 0 -148
box -98 -68 98 68
use sky130_fd_pr__pfet_01v8_u061qr  M2
timestamp 1604371879
transform 0 1 335 -1 0 1537
box -134 -142 134 142
use sky130_fd_pr__nfet_01v8_lca7f7  M1
timestamp 1604306825
transform 0 1 728 -1 0 1448
box -98 -68 98 68
use sky130_fd_pr__nfet_01v8_9hqhhq  Cv
timestamp 1604306825
transform 1 0 378 0 1 688
box -498 -526 498 526
use sky130_fd_pr__pfet_01v8_h2n75u  M3
timestamp 1604306825
transform 0 1 -8 -1 0 1537
box -134 -142 134 142
use sky130_fd_pr__pfet_01v8_6z4qh8  M9
timestamp 1604306825
transform 1 0 1863 0 1 1432
box -134 -142 134 142
use sky130_fd_pr__nfet_01v8_9i6r5e  M7
timestamp 1604306825
transform 1 0 1414 0 1 -65
box -98 -68 98 68
use sky130_fd_pr__pfet_01v8_2vaynq  M6
timestamp 1604306825
transform 1 0 1454 0 1 1432
box -134 -142 134 142
use sky130_fd_pr__nfet_01v8_tb02ql  Ca
timestamp 1604306825
transform 1 0 2868 0 1 916
box -618 -826 618 826
use sky130_fd_pr__nfet_01v8_wpylm8  Cu
timestamp 1604306825
transform 1 0 1617 0 1 661
box -388 -426 388 426
use sky130_fd_pr__nfet_01v8_dlksd1  M10
timestamp 1604306825
transform 1 0 2586 0 1 -154
box -98 -68 98 68
<< labels >>
rlabel metal1 -223 2059 -223 2059 1 vpwr
rlabel metal1 -143 -471 -143 -471 1 vgnd
rlabel metal1 -294 1383 -294 1383 1 vth
rlabel poly -66 -148 -66 -148 1 vk
rlabel poly 1456 1547 1456 1547 1 vw
rlabel poly 1406 -136 1406 -136 1 vr
rlabel poly 1867 1553 1867 1553 1 vau
rlabel poly 2587 -232 2587 -232 1 vad
rlabel locali -45 1274 -45 1274 1 v
rlabel locali 1441 1138 1441 1138 1 u#
rlabel locali 2619 1805 2619 1805 1 a#
rlabel metal2 1185 1178 1185 1178 1 axon
<< end >>
