magic
tech sky130A
timestamp 1608047394
<< metal1 >>
rect 1992 1550 2030 2024
rect 1766 1532 2030 1550
rect 1766 1510 2024 1532
rect 1876 1065 2013 1072
rect 1876 1055 2014 1065
rect 1986 946 2014 1055
rect 1986 920 2016 946
rect 1988 752 2016 920
<< metal2 >>
rect 213 1492 252 1739
rect 213 1465 1346 1492
rect 213 1159 252 1465
<< metal3 >>
rect 886 2015 930 2429
rect 886 1963 1089 2015
rect 886 1783 930 1963
rect 81 1154 122 1561
rect 886 1100 929 1783
rect 1100 1540 1268 1544
rect 1100 1535 1438 1540
rect 1098 1505 1438 1535
rect 1098 1433 1137 1505
rect 1246 1504 1438 1505
rect 1097 1400 1137 1433
rect 1097 1298 1136 1400
rect 886 1062 1095 1100
rect 1057 899 1095 1062
<< metal4 >>
rect 443 1164 488 1310
rect 472 1083 1491 1121
use 2good  2good_0
timestamp 1608047394
transform 1 0 98 0 1 604
box -97 -601 1925 738
use 2good  2good_1
timestamp 1608047394
transform 1 0 103 0 1 1850
box -97 -601 1925 738
use Sw-1  Sw-1_0
timestamp 1608047394
transform 1 0 1185 0 1 1008
box -70 45 891 509
<< end >>
