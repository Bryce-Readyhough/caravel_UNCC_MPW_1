magic
tech sky130A
magscale 1 2
timestamp 1608004133
<< locali >>
rect -180 1366 -114 1382
rect -184 1324 -174 1366
rect -120 1324 -110 1366
rect -180 1316 -114 1324
rect -180 1032 -114 1052
rect -184 988 -174 1032
rect -120 988 -110 1032
rect -180 970 -114 988
rect -184 744 -118 772
rect -188 700 -178 744
rect -122 700 -112 744
rect -184 694 -118 700
rect -184 412 -118 422
rect -188 368 -178 412
rect -124 368 -114 412
rect -184 346 -118 368
rect -100 42 -34 58
rect -104 -2 -94 42
rect -40 -2 -30 42
rect -100 -8 -34 -2
rect -102 -292 -34 -284
rect -106 -340 -96 -292
rect -38 -340 -28 -292
rect -102 -358 -34 -340
rect -180 -552 -114 -524
rect -184 -588 -174 -552
rect -120 -588 -110 -552
rect -180 -594 -114 -588
rect -180 -890 -114 -882
rect -184 -930 -174 -890
rect -120 -930 -110 -890
rect -180 -970 -114 -930
<< viali >>
rect -174 1324 -120 1366
rect -174 988 -120 1032
rect -178 700 -122 744
rect -178 368 -124 412
rect -94 -2 -40 42
rect -96 -340 -38 -292
rect -174 -588 -120 -552
rect -174 -930 -120 -890
<< metal1 >>
rect -194 1366 -100 1476
rect -190 1324 -174 1366
rect -120 1324 -106 1366
rect -190 1316 -106 1324
rect -174 1314 -120 1316
rect -188 1032 -102 1046
rect -188 988 -174 1032
rect -120 988 -102 1032
rect -188 974 -102 988
rect -160 930 -102 974
rect -160 886 148 930
rect -160 760 -102 886
rect -192 744 -102 760
rect -192 700 -178 744
rect -122 706 -102 744
rect -122 700 -108 706
rect -192 692 -108 700
rect -178 690 -122 692
rect 1892 690 2070 706
rect 1892 666 2078 690
rect 2044 534 2078 666
rect -178 420 -124 422
rect -192 416 -106 420
rect -192 412 -58 416
rect -192 368 -178 412
rect -124 368 -58 412
rect -192 354 -58 368
rect -112 56 -58 354
rect -112 52 -20 56
rect -112 42 138 52
rect -112 -2 -94 42
rect -40 4 138 42
rect -40 -2 -20 4
rect -112 -12 -20 -2
rect -96 -284 144 -282
rect -112 -292 144 -284
rect -112 -298 -96 -292
rect -126 -340 -96 -298
rect -38 -330 144 -292
rect -38 -340 -24 -330
rect -126 -348 -24 -340
rect -126 -350 -38 -348
rect -126 -536 -68 -350
rect 2060 -502 2098 -352
rect 1880 -536 2098 -502
rect -190 -552 -68 -536
rect -190 -588 -174 -552
rect -120 -580 -68 -552
rect -120 -588 -104 -580
rect -190 -594 -104 -588
rect -174 -598 -120 -594
rect -190 -890 -104 -878
rect -190 -930 -174 -890
rect -120 -930 -104 -890
rect -190 -944 -104 -930
rect -174 -1164 -116 -944
rect -174 -1190 168 -1164
rect -156 -1200 168 -1190
<< metal2 >>
rect 240 896 292 1146
rect 240 844 434 896
rect 240 522 292 844
rect 240 470 2388 522
rect 240 -310 292 470
rect 240 -362 434 -310
<< metal3 >>
rect -30 -637 31 1148
rect 1916 186 1995 631
<< metal4 >>
rect 693 145 763 1141
rect 638 75 763 145
rect 638 -224 708 75
rect 633 -294 2671 -224
rect 638 -1126 708 -294
use sky130_fd_pr__res_generic_po_0v6cx5  sky130_fd_pr__res_generic_po_0v6cx5_0
timestamp 1606707439
transform 1 0 -67 0 1 -150
box -33 -244 33 244
use sky130_fd_pr__res_generic_po_kabjgr  sky130_fd_pr__res_generic_po_kabjgr_0
timestamp 1606707439
transform 1 0 -151 0 1 556
box -33 -244 33 244
use sky130_fd_pr__res_generic_po_i65fu2  sky130_fd_pr__res_generic_po_i65fu2_0
timestamp 1606707439
transform 1 0 -147 0 1 -742
box -33 -244 33 244
use sky130_fd_pr__res_generic_po_abfehu  sky130_fd_pr__res_generic_po_abfehu_0
timestamp 1606707439
transform 1 0 -147 0 1 1176
box -33 -244 33 244
use Sw-1  Sw-1_2
timestamp 1608004133
transform 1 0 2068 0 1 -460
box -140 90 1782 1018
use Sw-1  Sw-1_1
timestamp 1608004133
transform 1 0 110 0 1 -1292
box -140 90 1782 1018
use Sw-1  Sw-1_0
timestamp 1608004133
transform 1 0 124 0 1 -86
box -140 90 1782 1018
<< end >>
