magic
tech sky130A
magscale 1 2
timestamp 1606262523
<< metal1 >>
rect 5316 27479 6214 27591
rect 6326 27479 6332 27591
rect 5376 27229 6660 27341
rect 6772 27229 6778 27341
rect 5463 26979 7083 27089
rect 7193 26979 7199 27089
rect -3277 26538 -3271 26780
rect -3029 26538 1072 26780
rect -2363 24048 -2357 24290
rect -2115 24048 1052 24290
rect 5401 23763 7527 23873
rect 7637 23763 7643 23873
rect 5480 23535 7934 23647
rect 8046 23535 8052 23647
rect 5464 23273 8356 23385
rect 8468 23273 8474 23385
rect 5410 21657 6214 21769
rect 6326 21657 6332 21769
rect 5322 21407 6664 21519
rect 6776 21407 6782 21519
rect 5475 21157 7087 21267
rect 7197 21157 7203 21267
rect -3277 20712 -3271 20954
rect -3029 20712 1066 20954
rect -2379 18226 -2373 18468
rect -2131 18226 1072 18468
rect 5429 17941 7531 18051
rect 7641 17941 7647 18051
rect 5470 17713 7940 17825
rect 8052 17713 8058 17825
rect 5486 17451 8356 17563
rect 8468 17451 8474 17563
rect 5322 15835 6214 15947
rect 6326 15835 6332 15947
rect 5432 15585 6660 15697
rect 6772 15585 6778 15697
rect 5489 15335 7093 15445
rect 7203 15335 7209 15445
rect -3293 14894 -3287 15136
rect -3045 15015 806 15136
rect -3045 14981 839 15015
rect -3045 14894 806 14981
rect -2363 12404 -2357 12646
rect -2115 12404 1002 12646
rect 5453 12119 7531 12229
rect 7641 12119 7647 12229
rect 5496 11891 7940 12003
rect 8052 11891 8058 12003
rect 5464 11629 8356 11741
rect 8468 11629 8474 11741
rect 5326 10013 6214 10125
rect 6326 10013 6332 10125
rect 5456 9763 6660 9875
rect 6772 9763 6778 9875
rect 5469 9513 7083 9623
rect 7193 9513 7199 9623
rect -3277 9074 -3271 9316
rect -3029 9074 930 9316
rect -2363 6584 -2357 6826
rect -2115 6584 968 6826
rect 5371 6297 7531 6407
rect 7641 6297 7647 6407
rect 5492 6069 7934 6181
rect 8046 6069 8052 6181
rect 5474 5807 8356 5919
rect 8468 5807 8474 5919
rect 5250 4191 6218 4303
rect 6330 4191 6336 4303
rect 5446 3941 6664 4053
rect 6776 3941 6782 4053
rect 5483 3691 7083 3801
rect 7193 3691 7199 3801
rect -3277 3250 -3271 3492
rect -3029 3375 840 3492
rect -3029 3341 895 3375
rect -3029 3250 840 3341
rect -2379 760 -2373 1002
rect -2131 760 842 1002
rect 5411 475 7531 585
rect 7641 475 7647 585
rect 5470 247 7940 359
rect 8052 247 8058 359
rect 5470 -15 8360 97
rect 8472 -15 8478 97
<< via1 >>
rect 6214 27479 6326 27591
rect 6660 27229 6772 27341
rect 7083 26979 7193 27089
rect -3271 26538 -3029 26780
rect -2357 24048 -2115 24290
rect 7527 23763 7637 23873
rect 7934 23535 8046 23647
rect 8356 23273 8468 23385
rect 6214 21657 6326 21769
rect 6664 21407 6776 21519
rect 7087 21157 7197 21267
rect -3271 20712 -3029 20954
rect -2373 18226 -2131 18468
rect 7531 17941 7641 18051
rect 7940 17713 8052 17825
rect 8356 17451 8468 17563
rect 6214 15835 6326 15947
rect 6660 15585 6772 15697
rect 7093 15335 7203 15445
rect -3287 14894 -3045 15136
rect -2357 12404 -2115 12646
rect 7531 12119 7641 12229
rect 7940 11891 8052 12003
rect 8356 11629 8468 11741
rect 6214 10013 6326 10125
rect 6660 9763 6772 9875
rect 7083 9513 7193 9623
rect -3271 9074 -3029 9316
rect -2357 6584 -2115 6826
rect 7531 6297 7641 6407
rect 7934 6069 8046 6181
rect 8356 5807 8468 5919
rect 6218 4191 6330 4303
rect 6664 3941 6776 4053
rect 7083 3691 7193 3801
rect -3271 3250 -3029 3492
rect -2373 760 -2131 1002
rect 7531 475 7641 585
rect 7940 247 8052 359
rect 8360 -15 8472 97
<< metal2 >>
rect -3271 26780 -3029 28725
rect -3271 20954 -3029 26538
rect -3271 15142 -3029 20712
rect -2357 24290 -2115 28709
rect -2357 18474 -2115 24048
rect -2373 18468 -2115 18474
rect -2131 18226 -2115 18468
rect -2373 18220 -2115 18226
rect -3287 15136 -3029 15142
rect -3045 14894 -3029 15136
rect -3287 14888 -3029 14894
rect -3271 9316 -3029 14888
rect -3271 3492 -3029 9074
rect -3271 -1787 -3029 3250
rect -2357 12646 -2115 18220
rect -2357 6826 -2115 12404
rect -2357 1008 -2115 6584
rect -2373 1002 -2115 1008
rect -2131 760 -2115 1002
rect -2373 754 -2115 760
rect -2357 -1787 -2115 754
rect 6214 27591 6326 28460
rect 6214 21769 6326 27479
rect 6214 15947 6326 21657
rect 6214 10125 6326 15835
rect 6214 4309 6326 10013
rect 6660 27341 6772 28480
rect 6660 21525 6772 27229
rect 7083 27089 7193 28487
rect 6660 21519 6776 21525
rect 6660 21407 6664 21519
rect 6660 21401 6776 21407
rect 6660 15697 6772 21401
rect 6660 9875 6772 15585
rect 6214 4303 6330 4309
rect 6214 4191 6218 4303
rect 6214 4185 6330 4191
rect 6214 -1736 6326 4185
rect 6660 4059 6772 9763
rect 7083 21273 7193 26979
rect 7527 23873 7637 28495
rect 7083 21267 7197 21273
rect 7083 21157 7087 21267
rect 7083 21151 7197 21157
rect 7083 15451 7193 21151
rect 7527 18057 7637 23763
rect 7934 23647 8046 28480
rect 7527 18051 7641 18057
rect 7527 17941 7531 18051
rect 7527 17935 7641 17941
rect 7083 15445 7203 15451
rect 7083 15335 7093 15445
rect 7083 15329 7203 15335
rect 7083 9623 7193 15329
rect 6660 4053 6776 4059
rect 6660 3941 6664 4053
rect 6660 3935 6776 3941
rect 6660 -1740 6772 3935
rect 7083 3801 7193 9513
rect 7083 -1745 7193 3691
rect 7527 12235 7637 17935
rect 7934 17831 8046 23535
rect 8356 23385 8468 28490
rect 7934 17825 8052 17831
rect 7934 17713 7940 17825
rect 7934 17707 8052 17713
rect 7527 12229 7641 12235
rect 7527 12119 7531 12229
rect 7527 12113 7641 12119
rect 7527 6413 7637 12113
rect 7934 12009 8046 17707
rect 8356 17563 8468 23273
rect 7934 12003 8052 12009
rect 7934 11891 7940 12003
rect 7934 11885 8052 11891
rect 7527 6407 7641 6413
rect 7527 6297 7531 6407
rect 7527 6291 7641 6297
rect 7527 591 7637 6291
rect 7934 6181 8046 11885
rect 7527 585 7641 591
rect 7527 475 7531 585
rect 7527 469 7641 475
rect 7527 -1759 7637 469
rect 7934 365 8046 6069
rect 8356 11741 8468 17451
rect 8356 5919 8468 11629
rect 7934 359 8052 365
rect 7934 247 7940 359
rect 7934 241 8052 247
rect 7934 -1774 8046 241
rect 8356 103 8468 5807
rect 8356 97 8472 103
rect 8356 -15 8360 97
rect 8356 -21 8472 -15
rect 8356 -1792 8468 -21
use neuron-labeled-extended  neuron-labeled-extended_0
array 0 0 5836 0 4 5822
timestamp 1606259729
transform 1 0 630 0 1 623
box -683 -638 4978 4166
<< end >>
