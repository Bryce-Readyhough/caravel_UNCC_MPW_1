magic
tech sky130A
timestamp 1608004133
<< metal1 >>
rect 16202 22417 16247 23211
rect 16171 22409 16265 22417
rect 16171 22340 16177 22409
rect 16260 22340 16265 22409
rect 16385 22400 16417 23130
rect 16619 23053 16685 23060
rect 16619 23012 16627 23053
rect 16679 23012 16685 23053
rect 16619 23006 16685 23012
rect 16627 22417 16668 23006
rect 16808 22948 16874 22954
rect 16808 22907 16813 22948
rect 16865 22907 16874 22948
rect 16808 22900 16874 22907
rect 16817 22420 16861 22900
rect 16990 22843 17056 22850
rect 16990 22802 16995 22843
rect 17047 22802 17056 22843
rect 16990 22796 17056 22802
rect 16600 22416 16689 22417
rect 16591 22409 16689 22416
rect 16171 22336 16265 22340
rect 16360 22392 16450 22400
rect 16360 22338 16368 22392
rect 16444 22338 16450 22392
rect 16360 22332 16450 22338
rect 16591 22343 16599 22409
rect 16683 22347 16689 22409
rect 16796 22416 16885 22420
rect 17000 22416 17040 22796
rect 17231 22740 17297 22747
rect 17231 22699 17237 22740
rect 17289 22699 17297 22740
rect 17231 22693 17297 22699
rect 16796 22355 16800 22416
rect 16881 22355 16885 22416
rect 16796 22351 16885 22355
rect 16980 22408 17062 22416
rect 17240 22411 17277 22693
rect 17435 22632 17516 22638
rect 17435 22589 17440 22632
rect 17510 22589 17516 22632
rect 17435 22584 17516 22589
rect 17449 22413 17491 22584
rect 18314 22542 18735 22547
rect 18302 22516 18735 22542
rect 16980 22353 16985 22408
rect 17058 22353 17062 22408
rect 16980 22347 17062 22353
rect 17217 22406 17300 22411
rect 16683 22343 16688 22347
rect 16591 22336 16688 22343
rect 17217 22346 17223 22406
rect 17297 22346 17300 22406
rect 17217 22342 17300 22346
rect 17436 22405 17520 22413
rect 17436 22348 17444 22405
rect 17513 22348 17520 22405
rect 17436 22344 17520 22348
rect 9536 22096 9579 22106
rect 18302 22096 18336 22516
rect 9536 22040 18348 22096
rect 19358 22095 19595 22097
rect 19358 22070 19602 22095
rect 9536 21652 9579 22040
rect 9534 21594 9579 21652
rect 9534 21488 9568 21594
rect 19579 21521 19602 22070
rect 19526 21504 19615 21521
<< via1 >>
rect 16177 22340 16260 22409
rect 16627 23012 16679 23053
rect 16813 22907 16865 22948
rect 16995 22802 17047 22843
rect 16368 22338 16444 22392
rect 16599 22343 16683 22409
rect 17237 22699 17289 22740
rect 16800 22355 16881 22416
rect 17440 22589 17510 22632
rect 16985 22353 17058 22408
rect 17223 22346 17297 22406
rect 17444 22348 17513 22405
<< metal2 >>
rect 16197 23228 16265 23234
rect 16197 23191 16203 23228
rect 16259 23191 16265 23228
rect 16197 23185 16265 23191
rect 16371 23140 16430 23149
rect 16371 23110 16380 23140
rect 16423 23110 16430 23140
rect 16371 23102 16430 23110
rect 16617 23055 16686 23062
rect 16617 23011 16625 23055
rect 16680 23011 16686 23055
rect 16617 23005 16686 23011
rect 16807 22948 16873 22954
rect 16807 22906 16813 22948
rect 16867 22906 16873 22948
rect 16807 22900 16873 22906
rect 16989 22844 17055 22850
rect 16989 22802 16995 22844
rect 17049 22802 17055 22844
rect 16989 22796 17055 22802
rect 17230 22741 17296 22747
rect 17230 22699 17236 22741
rect 17290 22699 17296 22741
rect 17230 22693 17296 22699
rect 17434 22632 17516 22638
rect 17434 22589 17440 22632
rect 17510 22589 17516 22632
rect 17434 22583 17516 22589
rect 18436 22483 18824 22523
rect 16169 22409 16268 22415
rect 16169 22340 16177 22409
rect 16260 22340 16268 22409
rect 16590 22409 16689 22417
rect 16169 22337 16179 22340
rect 16259 22337 16268 22340
rect 16169 22331 16268 22337
rect 16359 22397 16453 22401
rect 16359 22395 16463 22397
rect 16359 22332 16367 22395
rect 16449 22332 16463 22395
rect 16590 22338 16599 22409
rect 16683 22343 16689 22409
rect 16794 22416 16889 22422
rect 16794 22414 16800 22416
rect 16881 22414 16889 22416
rect 16794 22353 16799 22414
rect 16883 22353 16889 22414
rect 16794 22347 16889 22353
rect 16978 22408 17066 22414
rect 16978 22348 16985 22408
rect 17058 22407 17066 22408
rect 17061 22348 17066 22407
rect 16978 22344 17066 22348
rect 17216 22406 17306 22413
rect 17216 22346 17223 22406
rect 17216 22345 17225 22346
rect 17297 22345 17306 22406
rect 16680 22338 16689 22343
rect 17216 22339 17306 22345
rect 17437 22405 17521 22413
rect 17437 22346 17444 22405
rect 17515 22346 17521 22405
rect 17437 22341 17521 22346
rect 16590 22332 16689 22338
rect 16359 22328 16463 22332
rect 16360 22323 16463 22328
rect 18447 21594 18492 22483
<< via2 >>
rect 16203 23191 16259 23228
rect 16380 23110 16423 23140
rect 16625 23053 16680 23055
rect 16625 23012 16627 23053
rect 16627 23012 16679 23053
rect 16679 23012 16680 23053
rect 16625 23011 16680 23012
rect 16813 22907 16865 22948
rect 16865 22907 16867 22948
rect 16813 22906 16867 22907
rect 16995 22843 17049 22844
rect 16995 22802 17047 22843
rect 17047 22802 17049 22843
rect 17236 22740 17290 22741
rect 17236 22699 17237 22740
rect 17237 22699 17289 22740
rect 17289 22699 17290 22740
rect 17440 22589 17510 22632
rect 16179 22340 16259 22404
rect 16179 22337 16259 22340
rect 16367 22392 16449 22395
rect 16367 22338 16368 22392
rect 16368 22338 16444 22392
rect 16444 22338 16449 22392
rect 16367 22332 16449 22338
rect 16599 22343 16680 22408
rect 16799 22355 16800 22414
rect 16800 22355 16881 22414
rect 16881 22355 16883 22414
rect 16799 22353 16883 22355
rect 16985 22353 17058 22407
rect 17058 22353 17061 22407
rect 16985 22348 17061 22353
rect 17225 22346 17297 22406
rect 17225 22345 17297 22346
rect 16599 22338 16680 22343
rect 17444 22348 17513 22405
rect 17513 22348 17515 22405
rect 17444 22346 17515 22348
<< metal3 >>
rect 6208 23228 6254 23259
rect 16199 23228 16263 23233
rect 6208 23192 16203 23228
rect 6208 21873 6254 23192
rect 16199 23191 16203 23192
rect 16259 23191 16263 23228
rect 16199 23187 16263 23191
rect 6440 23140 16433 23145
rect 6440 23138 16380 23140
rect 6414 23110 16380 23138
rect 16423 23110 16433 23140
rect 6414 23107 16433 23110
rect 6414 21795 6477 23107
rect 6593 23057 6652 23061
rect 16620 23057 16685 23058
rect 6593 23055 16685 23057
rect 6593 23011 16625 23055
rect 16680 23011 16685 23055
rect 6593 23009 16685 23011
rect 6593 21698 6652 23009
rect 16620 23008 16685 23009
rect 6794 22948 16877 22954
rect 6794 22913 16813 22948
rect 6775 22906 16813 22913
rect 16867 22906 16877 22948
rect 6775 22901 16877 22906
rect 6775 21611 6837 22901
rect 6976 22844 17053 22847
rect 6976 22808 16995 22844
rect 6958 22802 16995 22808
rect 17049 22802 17053 22844
rect 6958 22797 17053 22802
rect 6958 21515 7029 22797
rect 7276 22743 17295 22744
rect 7253 22741 17295 22743
rect 7253 22699 17236 22741
rect 17290 22699 17295 22741
rect 7253 22696 17295 22699
rect 7253 21385 7317 22696
rect 7485 22635 7548 22639
rect 17433 22635 17515 22637
rect 7485 22632 17515 22635
rect 7485 22589 17440 22632
rect 17510 22589 17515 22632
rect 7485 22587 17515 22589
rect 7485 21269 7548 22587
rect 17433 22584 17515 22587
rect 7628 22461 18079 22517
rect 7638 22147 7683 22461
rect 16167 22404 16272 22415
rect 16590 22408 16693 22419
rect 16167 22337 16179 22404
rect 16259 22337 16272 22404
rect 16167 22299 16272 22337
rect 16356 22395 16462 22404
rect 16356 22332 16367 22395
rect 16449 22332 16462 22395
rect 16590 22346 16599 22408
rect 7638 22073 7695 22147
rect 7644 21474 7695 22073
rect 16187 21877 16255 22299
rect 16356 22293 16462 22332
rect 16580 22338 16599 22346
rect 16680 22338 16693 22408
rect 16793 22414 16892 22425
rect 16793 22353 16799 22414
rect 16883 22353 16892 22414
rect 16793 22350 16892 22353
rect 16388 21799 16451 22293
rect 16580 22292 16693 22338
rect 16774 22299 16892 22350
rect 16979 22407 17069 22415
rect 16979 22348 16985 22407
rect 17061 22348 17069 22407
rect 16979 22346 17069 22348
rect 16976 22301 17069 22346
rect 17217 22406 17307 22417
rect 17217 22345 17225 22406
rect 17297 22345 17307 22406
rect 16580 21708 16658 22292
rect 16774 21620 16856 22299
rect 16976 21519 17042 22301
rect 17217 22300 17307 22345
rect 17436 22405 17524 22413
rect 17436 22346 17444 22405
rect 17515 22346 17524 22405
rect 17436 22306 17524 22346
rect 7638 21430 8633 21474
rect 17221 21371 17285 22300
rect 17453 21253 17506 22306
rect 18001 21485 18067 22461
rect 18001 21464 18605 21485
rect 18018 21419 18605 21464
<< metal4 >>
rect 18916 21220 18958 22150
use 8good  8good_0
timestamp 1608004133
transform 1 0 -2 0 1 7
box -1 -8 9928 21979
use 8good  8good_1
timestamp 1608004133
transform 1 0 9983 0 1 10
box -1 -8 9928 21979
use Sw-1  Sw-1_0
timestamp 1608004133
transform 1 0 18665 0 1 22033
box -70 45 891 509
<< end >>
