magic
tech sky130A
magscale 1 2
timestamp 1606105257
<< nwell >>
rect -109 -123 109 123
<< pmos >>
rect -15 -61 15 23
<< pdiff >>
rect -73 11 -15 23
rect -73 -49 -61 11
rect -27 -49 -15 11
rect -73 -61 -15 -49
rect 15 11 73 23
rect 15 -49 27 11
rect 61 -49 73 11
rect 15 -61 73 -49
<< pdiffc >>
rect -61 -49 -27 11
rect 27 -49 61 11
<< poly >>
rect -33 104 33 120
rect -33 70 -17 104
rect 17 70 33 104
rect -33 54 33 70
rect -15 23 15 54
rect -15 -87 15 -61
<< polycont >>
rect -17 70 17 104
<< locali >>
rect -33 70 -17 104
rect 17 70 33 104
rect -61 11 -27 27
rect -61 -65 -27 -49
rect 27 11 61 27
rect 27 -65 61 -49
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.42 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0
string library sky130
<< end >>
