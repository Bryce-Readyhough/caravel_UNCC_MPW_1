* NGSPICE file created from testing.ext - technology: sky130A

* Include SkyWater sky130 device models
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical__lin.spice"
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical.spice"
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"

* DC source for current measure
Vdd vdd gnd DC 0.7V
Vgnd vss gnd DC 0.0V
Vth vth gnd DC 0.1V
Vk vk gnd DC 0.15V
Vw vw gnd DC 0.18V
Vr vr gnd DC 0.2V
Vau vau gnd DC 0.23V
Vad vad gnd DC 0.1V

* DC source for current measure
* Vdd vdd gnd DC 0.7V
* Vgnd vss gnd DC 0.0V
* Vth vth gnd DC 0.1V
* Vk vk gnd DC 0.15V
* Vw vw gnd DC 0.01V
* Vr vr gnd DC 0.37V
* Vau vau gnd DC 0.1V
* Vad vad gnd DC 0.2V

Idc vdd v DC 5p
vsyn0 syn0 gnd DC 0.42
vsyn1 syn1 gnd DC 0.42
Vsel sel gnd DC 0.0

* NGSPICE file created from testing.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_owy61o VSUBS a_n73_n61# w_n109_n123# a_15_n61# a_n33_54#
X0 a_15_n61# a_n33_54# a_n73_n61# w_n109_n123# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_63vi9a VSUBS a_15_n11# a_n33_n99# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt one-way VSUBS li_12_16# w_n37_405# li_100_394#
Xsky130_fd_pr__pfet_01v8_owy61o_0 VSUBS li_12_16# w_n37_405# li_100_394# li_100_394#
+ sky130_fd_pr__pfet_01v8_owy61o
Xsky130_fd_pr__nfet_01v8_63vi9a_0 VSUBS li_100_394# li_12_16# li_12_16# sky130_fd_pr__nfet_01v8_63vi9a
.ends

.subckt sky130_fd_pr__nfet_01v8_8mr83b VSUBS a_n73_n42# a_n15_n68# a_15_n42#
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_ykwexw VSUBS a_n73_n42# w_n109_n104# a_n15_n68# a_15_n42#
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt inverter GND in VPWR out
Xsky130_fd_pr__nfet_01v8_8mr83b_0 GND GND in out sky130_fd_pr__nfet_01v8_8mr83b
Xsky130_fd_pr__pfet_01v8_ykwexw_0 GND VPWR VPWR in out sky130_fd_pr__pfet_01v8_ykwexw
.ends

.subckt sky130_fd_pr__nfet_01v8_dlksd1 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_s3efqo VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lca7f7 VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_u061qr VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_h2n75u VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_zt2j7p VSUBS a_n98_n120# a_n40_n146# a_40_n120# w_n134_n182#
X0 a_40_n120# a_n40_n146# a_n98_n120# w_n134_n182# sky130_fd_pr__pfet_01v8 w=1.2e+06u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ckptud VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_2vaynq VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_wpylm8 VSUBS a_n388_n400# a_n330_n426# a_330_n400#
X0 a_330_n400# a_n330_n426# a_n388_n400# VSUBS sky130_fd_pr__nfet_01v8 w=4e+06u l=3.3e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_9i6r5e VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_9hqhhq VSUBS a_n498_n500# a_n440_n526# a_440_n500#
X0 a_440_n500# a_n440_n526# a_n498_n500# VSUBS sky130_fd_pr__nfet_01v8 w=5e+06u l=4.4e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_h43ndc VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_6z4qh8 VSUBS a_n40_n106# a_n98_n80# w_n134_n142# a_40_n80#
X0 a_40_n80# a_n40_n106# a_n98_n80# w_n134_n142# sky130_fd_pr__pfet_01v8 w=800000u l=400000u
.ends

.subckt sky130_fd_pr__nfet_01v8_tb02ql VSUBS a_n618_n800# a_n560_n826# a_560_n800#
X0 a_560_n800# a_n560_n826# a_n618_n800# VSUBS sky130_fd_pr__nfet_01v8 w=8e+06u l=5.6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_zgaw3c VSUBS a_n98_n42# a_n40_n68# a_40_n42#
X0 a_40_n42# a_n40_n68# a_n98_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=400000u
.ends

.subckt neuron-labeled VPWR VGND vth vk vw vr vau vad v u# a# axon
XM10 VGND VGND vad a# sky130_fd_pr__nfet_01v8_dlksd1
XM11 VGND v a# VGND sky130_fd_pr__nfet_01v8_s3efqo
XM1 VGND a_35_1497# v vth sky130_fd_pr__nfet_01v8_lca7f7
XM2 VGND a_35_1497# VPWR VPWR a_35_1497# sky130_fd_pr__pfet_01v8_u061qr
XM3 VGND a_35_1497# VPWR VPWR v sky130_fd_pr__pfet_01v8_h2n75u
XM4 VGND VPWR a_35_1497# axon VPWR sky130_fd_pr__pfet_01v8_zt2j7p
XM5 VGND VGND a_35_1497# axon sky130_fd_pr__nfet_01v8_ckptud
XM6 VGND vw axon VPWR u# sky130_fd_pr__pfet_01v8_2vaynq
XCu VGND VGND u# VGND sky130_fd_pr__nfet_01v8_wpylm8
XM7 VGND VGND vr u# sky130_fd_pr__nfet_01v8_9i6r5e
XCv VGND VGND v VGND sky130_fd_pr__nfet_01v8_9hqhhq
XM8 VGND v u# VGND sky130_fd_pr__nfet_01v8_h43ndc
XM9 VGND vau axon VPWR a# sky130_fd_pr__pfet_01v8_6z4qh8
XCa VGND VGND a# VGND sky130_fd_pr__nfet_01v8_tb02ql
XMk VGND v vk VGND sky130_fd_pr__nfet_01v8_zgaw3c
.ends

.subckt neuron-labeled-extended vk vdd vss vr vad u v vau vw vth a axon vss vdd v
+ neuron-labeled_0/vth li_3628_2434# neuron-labeled_0/vau neuron-labeled_0/vw neuron-labeled_0/axon
+ vss
Xneuron-labeled_0 vdd vss neuron-labeled_0/vth vk neuron-labeled_0/vw vr neuron-labeled_0/vau
+ vad v u li_3628_2434# neuron-labeled_0/axon neuron-labeled
.ends

.subckt sky130_fd_pr__nfet_01v8_5mkfxl VSUBS a_n73_n42# a_15_n42# a_n33_n130#
X0 a_15_n42# a_n33_n130# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_pa2hmj VSUBS a_n33_n177# a_15_n80# w_n109_n180# a_n73_n80#
X0 a_15_n80# a_n33_n177# a_n73_n80# w_n109_n180# sky130_fd_pr__pfet_01v8 w=800000u l=150000u
.ends

.subckt pass-gate clk clk_bar v_in v_out v_newll v_sub
Xsky130_fd_pr__nfet_01v8_5mkfxl_0 v_sub v_out v_in clk sky130_fd_pr__nfet_01v8_5mkfxl
Xsky130_fd_pr__pfet_01v8_pa2hmj_0 v_sub clk_bar v_out v_newll v_in sky130_fd_pr__pfet_01v8_pa2hmj
.ends

.subckt pass-gate-inv-2 v_in v_out clk clk_bar VPWR VGND v_in2 VGND VPWR v_out clk
+ VGND VPWR
Xinverter_0 VGND clk VPWR clk_bar inverter
Xpass-gate_0 clk clk_bar v_in v_out VPWR VGND pass-gate
Xpass-gate_1 clk_bar clk v_in2 v_out VPWR VGND pass-gate
.ends

.subckt testing vw vth vk vr vad v u a axon sel v# u# a# axon# syn0 syn1 vdd vss vau
Xone-way_0 vss inverter_0/out vdd pass-gate-inv-2_0/v_in one-way
Xone-way_1 vss inverter_1/out vdd pass-gate-inv-2_0/v_in2 one-way
Xinverter_0 vss syn1 vdd inverter_0/out inverter
Xinverter_1 vss syn0 vdd inverter_1/out inverter
Xneuron-labeled-extended_0 vk vdd vss vr vad pass-gate-inv-2_1/v_in pass-gate-inv-2_0/v_in
+ neuron-labeled-extended_0/vau neuron-labeled-extended_0/vw neuron-labeled-extended_0/vth
+ neuron-labeled-extended_0/a neuron-labeled-extended_0/axon vss vdd pass-gate-inv-2_0/v_in
+ vth pass-gate-inv-2_2/v_in vau vw pass-gate-inv-2_3/v_in vss neuron-labeled-extended
Xpass-gate-inv-2_0 pass-gate-inv-2_0/v_in v# sel pass-gate-inv-2_0/clk_bar vdd vss
+ pass-gate-inv-2_0/v_in2 vss vdd v# sel vss pass-gate-inv-2_0/inverter_0/VPWR pass-gate-inv-2
Xneuron-labeled-extended_1 vk vdd vss vr vad pass-gate-inv-2_1/v_in2 pass-gate-inv-2_0/v_in2
+ neuron-labeled-extended_1/vau neuron-labeled-extended_1/vw neuron-labeled-extended_1/vth
+ neuron-labeled-extended_1/a neuron-labeled-extended_1/axon vss vdd pass-gate-inv-2_0/v_in2
+ vth pass-gate-inv-2_2/v_in2 vau vw pass-gate-inv-2_3/v_in2 vss neuron-labeled-extended
Xpass-gate-inv-2_1 pass-gate-inv-2_1/v_in u# sel pass-gate-inv-2_1/clk_bar vdd vss
+ pass-gate-inv-2_1/v_in2 vss vdd u# sel vss vdd pass-gate-inv-2
Xneuron-labeled-extended_2 vk vdd vss vr vad u v neuron-labeled-extended_2/vau neuron-labeled-extended_2/vw
+ neuron-labeled-extended_2/vth neuron-labeled-extended_2/a neuron-labeled-extended_2/axon
+ vss vdd v vth a vau vw axon vss neuron-labeled-extended
Xpass-gate-inv-2_2 pass-gate-inv-2_2/v_in a# sel pass-gate-inv-2_2/clk_bar vdd vss
+ pass-gate-inv-2_2/v_in2 vss vdd a# sel vss pass-gate-inv-2_2/inverter_0/VPWR pass-gate-inv-2
Xpass-gate-inv-2_3 pass-gate-inv-2_3/v_in axon# sel pass-gate-inv-2_3/clk_bar vdd
+ vss pass-gate-inv-2_3/v_in2 vss vdd axon# sel vss pass-gate-inv-2_3/inverter_0/VPWR
+ pass-gate-inv-2
.ends





* instantiate
Xtest vw vth vk vr vad v u a axon sel v# u# a# axon# syn0 syn1 vdd vss vau testing

*.IC V(v)=0 V(u#)=0 V(a#)=0

.control
* Sweep tran
tran 1u 50m uic
plot v(v) v(u)
plot v("xtest.neuron-labeled-extended_0/v") v("xtest.neuron-labeled-extended_0/u")

* dc vsyn0 0 0.7 0.01
* plot v("xtest.inverter_0[0]/out")
.endc
.end


